module fake_netlist_1_8575_n_1319 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1319);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1319;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_659;
wire n_432;
wire n_386;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
BUFx3_ASAP7_75t_L g360 ( .A(n_152), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_334), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_283), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
INVxp33_ASAP7_75t_SL g364 ( .A(n_243), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_48), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_359), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_121), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_114), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_51), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_291), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_183), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_232), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_119), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_270), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_248), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_176), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_133), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_90), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_256), .B(n_119), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_189), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_4), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_100), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_246), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_122), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_118), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_205), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_102), .Y(n_389) );
HB1xp67_ASAP7_75t_SL g390 ( .A(n_227), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_294), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_72), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_82), .Y(n_394) );
INVxp33_ASAP7_75t_SL g395 ( .A(n_274), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_123), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_326), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_279), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_349), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_111), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_79), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_32), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_21), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_39), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_300), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_74), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_130), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_38), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_141), .Y(n_409) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_76), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_153), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_18), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_213), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_106), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_240), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_348), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_320), .B(n_312), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_319), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_341), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_216), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_321), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_199), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_72), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_71), .B(n_147), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_217), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_223), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_12), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_48), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_90), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_89), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_271), .B(n_352), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_112), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_49), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_134), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_22), .B(n_164), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_0), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_78), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_278), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_259), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_54), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_30), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_325), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_203), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_273), .Y(n_444) );
INVxp33_ASAP7_75t_SL g445 ( .A(n_269), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_206), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_191), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_310), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_23), .Y(n_449) );
INVxp33_ASAP7_75t_L g450 ( .A(n_340), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_323), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_182), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_293), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_61), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_113), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_83), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_32), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_126), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_150), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_89), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_184), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_115), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_143), .Y(n_463) );
BUFx2_ASAP7_75t_SL g464 ( .A(n_99), .Y(n_464) );
BUFx2_ASAP7_75t_SL g465 ( .A(n_109), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_170), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_165), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_180), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_0), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_13), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_156), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_212), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_63), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_73), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_45), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_42), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_14), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_238), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_148), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_237), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_219), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_357), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_221), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_263), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_236), .Y(n_485) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_84), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_275), .Y(n_487) );
INVxp33_ASAP7_75t_SL g488 ( .A(n_116), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_124), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_169), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_337), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_47), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_254), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_162), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_267), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_132), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_302), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_140), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_231), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_76), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_353), .Y(n_501) );
INVxp33_ASAP7_75t_SL g502 ( .A(n_25), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_296), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_15), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_84), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_99), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_261), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_142), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_255), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_137), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_260), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_102), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_358), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_324), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_8), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_115), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_42), .B(n_112), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_197), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_6), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_19), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_214), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_34), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_299), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_95), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_168), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_98), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_332), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_88), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_322), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_233), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_245), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_69), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_34), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_215), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_304), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_167), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_16), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_249), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_78), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g540 ( .A(n_52), .B(n_250), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_155), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_262), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_117), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_450), .B(n_1), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_369), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_472), .B(n_1), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_369), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_450), .B(n_2), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_414), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_388), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_507), .B(n_414), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_441), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_457), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_374), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_507), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_449), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_380), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_507), .B(n_3), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_380), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_371), .B(n_375), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_518), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_413), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_449), .B(n_5), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_443), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_362), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_486), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_362), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_527), .B(n_7), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_363), .B(n_9), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_368), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_400), .B(n_10), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_368), .Y(n_573) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_360), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_400), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_372), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_374), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_390), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_372), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_401), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_402), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_578), .B(n_478), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_555), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_555), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_561), .B(n_495), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_552), .B(n_448), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_555), .Y(n_587) );
INVx4_ASAP7_75t_L g588 ( .A(n_558), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_555), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_555), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_555), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_561), .B(n_484), .Y(n_592) );
INVx4_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
INVx4_ASAP7_75t_L g594 ( .A(n_558), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_558), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_560), .B(n_408), .C(n_404), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_554), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_567), .A2(n_404), .B1(n_432), .B2(n_408), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_581), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_544), .B(n_487), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_574), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_566), .Y(n_605) );
BUFx4_ASAP7_75t_L g606 ( .A(n_546), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_568), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_551), .B(n_361), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_574), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_544), .B(n_456), .C(n_432), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_574), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_581), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_563), .B(n_427), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_550), .B(n_523), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_548), .B(n_565), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_549), .Y(n_618) );
OR2x6_ASAP7_75t_L g619 ( .A(n_553), .B(n_464), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_611), .Y(n_620) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_611), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_599), .A2(n_569), .B(n_546), .C(n_553), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_604), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_588), .B(n_563), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
NOR2x1p5_ASAP7_75t_L g627 ( .A(n_592), .B(n_562), .Y(n_627) );
NOR2x1p5_ASAP7_75t_L g628 ( .A(n_592), .B(n_564), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_600), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_585), .B(n_548), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_604), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_614), .B(n_569), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_583), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_604), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_618), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_588), .B(n_563), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_586), .B(n_549), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_597), .B(n_549), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_595), .A2(n_556), .B(n_549), .Y(n_639) );
INVx3_ASAP7_75t_SL g640 ( .A(n_619), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_601), .B(n_556), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_617), .A2(n_572), .B(n_488), .C(n_502), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_618), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_588), .B(n_572), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_609), .B(n_570), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_617), .B(n_556), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_616), .B(n_460), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_583), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_618), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_593), .B(n_572), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_612), .B(n_364), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_593), .B(n_365), .Y(n_653) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_619), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_595), .A2(n_571), .B1(n_573), .B2(n_568), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_598), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_582), .B(n_567), .Y(n_658) );
INVx11_ASAP7_75t_L g659 ( .A(n_606), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_593), .B(n_361), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_619), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_615), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_593), .B(n_391), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_589), .Y(n_664) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_594), .B(n_431), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_589), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_594), .B(n_373), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_615), .A2(n_573), .B1(n_576), .B2(n_571), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_594), .B(n_376), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_615), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_594), .B(n_377), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_596), .B(n_379), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_602), .B(n_460), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_605), .B(n_382), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_605), .Y(n_676) );
OR2x6_ASAP7_75t_L g677 ( .A(n_607), .B(n_465), .Y(n_677) );
AO22x1_ASAP7_75t_L g678 ( .A1(n_607), .A2(n_445), .B1(n_395), .B2(n_462), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_608), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_608), .A2(n_573), .B1(n_576), .B2(n_571), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_584), .A2(n_444), .B1(n_493), .B2(n_378), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_589), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_589), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_584), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_629), .B(n_577), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_676), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_659), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_632), .B(n_383), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_684), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_620), .Y(n_690) );
INVx3_ASAP7_75t_L g691 ( .A(n_620), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_654), .B(n_391), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_620), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_657), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_624), .B(n_576), .Y(n_695) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_681), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_627), .B(n_378), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_642), .A2(n_470), .B(n_473), .C(n_410), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_673), .B(n_462), .Y(n_699) );
OAI22xp5_ASAP7_75t_SL g700 ( .A1(n_658), .A2(n_430), .B1(n_526), .B2(n_383), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_652), .A2(n_424), .B(n_381), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_630), .A2(n_579), .B(n_366), .C(n_384), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_620), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_648), .B(n_430), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_677), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_662), .Y(n_706) );
NAND2xp33_ASAP7_75t_L g707 ( .A(n_640), .B(n_444), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_677), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_621), .Y(n_709) );
CKINVDCx6p67_ASAP7_75t_R g710 ( .A(n_658), .Y(n_710) );
OAI21x1_ASAP7_75t_L g711 ( .A1(n_683), .A2(n_587), .B(n_590), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_621), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_670), .Y(n_713) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_621), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_665), .B(n_505), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_645), .A2(n_579), .B(n_370), .C(n_389), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_645), .A2(n_579), .B(n_393), .C(n_394), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_636), .A2(n_587), .B(n_603), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_665), .A2(n_531), .B1(n_536), .B2(n_535), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_621), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_635), .Y(n_721) );
BUFx12f_ASAP7_75t_L g722 ( .A(n_628), .Y(n_722) );
INVx5_ASAP7_75t_L g723 ( .A(n_679), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_635), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_651), .A2(n_403), .B(n_406), .C(n_387), .Y(n_725) );
INVx4_ASAP7_75t_L g726 ( .A(n_650), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_622), .A2(n_423), .B(n_428), .C(n_412), .Y(n_727) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_650), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_678), .B(n_532), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_647), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_652), .B(n_535), .Y(n_731) );
INVx5_ASAP7_75t_L g732 ( .A(n_661), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_641), .A2(n_433), .B(n_436), .C(n_429), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_636), .A2(n_454), .B1(n_455), .B2(n_437), .Y(n_734) );
INVx4_ASAP7_75t_L g735 ( .A(n_682), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_653), .A2(n_669), .B(n_667), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_660), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_637), .A2(n_533), .B1(n_539), .B2(n_477), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_643), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_663), .B(n_533), .Y(n_740) );
BUFx2_ASAP7_75t_L g741 ( .A(n_639), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_644), .A2(n_469), .B(n_475), .C(n_474), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_668), .B(n_539), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_644), .Y(n_744) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_623), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_683), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_638), .B(n_517), .Y(n_747) );
INVx4_ASAP7_75t_L g748 ( .A(n_623), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_653), .B(n_476), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_623), .Y(n_750) );
AND2x2_ASAP7_75t_SL g751 ( .A(n_668), .B(n_440), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_656), .B(n_396), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_623), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_672), .Y(n_754) );
BUFx12f_ASAP7_75t_L g755 ( .A(n_631), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_656), .A2(n_504), .B1(n_506), .B2(n_500), .Y(n_756) );
NOR2xp67_ASAP7_75t_L g757 ( .A(n_671), .B(n_120), .Y(n_757) );
BUFx2_ASAP7_75t_L g758 ( .A(n_631), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_680), .B(n_575), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_675), .A2(n_512), .B1(n_516), .B2(n_515), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_675), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_680), .Y(n_762) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_631), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_625), .A2(n_386), .B(n_385), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_625), .B(n_519), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_631), .Y(n_766) );
AOI21xp33_ASAP7_75t_L g767 ( .A1(n_626), .A2(n_503), .B(n_405), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_634), .Y(n_768) );
NOR2xp67_ASAP7_75t_SL g769 ( .A(n_634), .B(n_397), .Y(n_769) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_634), .Y(n_770) );
OAI21x1_ASAP7_75t_L g771 ( .A1(n_626), .A2(n_610), .B(n_603), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_634), .B(n_520), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_633), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g774 ( .A(n_646), .B(n_397), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_649), .A2(n_522), .B(n_543), .C(n_524), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_649), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_655), .A2(n_398), .B1(n_415), .B2(n_407), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_674), .Y(n_778) );
BUFx2_ASAP7_75t_L g779 ( .A(n_674), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_664), .B(n_440), .Y(n_780) );
BUFx4f_ASAP7_75t_L g781 ( .A(n_664), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_666), .B(n_528), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_666), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_620), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_620), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_665), .A2(n_537), .B1(n_528), .B2(n_574), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_632), .B(n_399), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_665), .B(n_537), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_673), .B(n_399), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_624), .A2(n_610), .B(n_591), .Y(n_790) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_652), .A2(n_419), .B(n_418), .Y(n_791) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_620), .Y(n_792) );
O2A1O1Ixp33_ASAP7_75t_L g793 ( .A1(n_642), .A2(n_547), .B(n_557), .C(n_545), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_630), .A2(n_540), .B(n_435), .C(n_545), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_710), .A2(n_420), .B1(n_422), .B2(n_421), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_794), .B(n_574), .C(n_589), .Y(n_796) );
AOI21xp33_ASAP7_75t_L g797 ( .A1(n_751), .A2(n_426), .B(n_425), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_744), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_719), .A2(n_557), .B1(n_559), .B2(n_547), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_771), .A2(n_411), .B(n_392), .Y(n_800) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_755), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_790), .A2(n_591), .B(n_411), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_689), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_786), .A2(n_580), .B1(n_559), .B2(n_575), .Y(n_804) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_745), .Y(n_805) );
INVx5_ASAP7_75t_L g806 ( .A(n_690), .Y(n_806) );
OA21x2_ASAP7_75t_L g807 ( .A1(n_711), .A2(n_452), .B(n_392), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_718), .A2(n_591), .B(n_482), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_749), .Y(n_809) );
AOI21xp33_ASAP7_75t_L g810 ( .A1(n_775), .A2(n_439), .B(n_434), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_727), .B(n_591), .C(n_604), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_762), .A2(n_417), .B(n_442), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_705), .B(n_580), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_736), .A2(n_447), .B(n_446), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_688), .B(n_416), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_753), .A2(n_501), .B(n_491), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_719), .A2(n_451), .B1(n_459), .B2(n_458), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_696), .A2(n_461), .B1(n_467), .B2(n_463), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_772), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_753), .A2(n_501), .B(n_491), .Y(n_820) );
NAND2x1p5_ASAP7_75t_L g821 ( .A(n_723), .B(n_360), .Y(n_821) );
AO21x2_ASAP7_75t_L g822 ( .A1(n_764), .A2(n_479), .B(n_471), .Y(n_822) );
AO21x2_ASAP7_75t_L g823 ( .A1(n_764), .A2(n_481), .B(n_480), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_704), .A2(n_489), .B1(n_490), .B2(n_485), .Y(n_824) );
NOR2xp67_ASAP7_75t_L g825 ( .A(n_687), .B(n_10), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_730), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_700), .A2(n_494), .B1(n_497), .B2(n_496), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_694), .Y(n_828) );
OAI21x1_ASAP7_75t_L g829 ( .A1(n_766), .A2(n_534), .B(n_499), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_780), .A2(n_509), .B(n_498), .Y(n_830) );
BUFx3_ASAP7_75t_L g831 ( .A(n_722), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_768), .A2(n_514), .B(n_513), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_759), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_706), .B(n_521), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_723), .Y(n_835) );
OR2x6_ASAP7_75t_L g836 ( .A(n_708), .B(n_525), .Y(n_836) );
INVx3_ASAP7_75t_L g837 ( .A(n_726), .Y(n_837) );
AOI22x1_ASAP7_75t_L g838 ( .A1(n_750), .A2(n_604), .B1(n_613), .B2(n_591), .Y(n_838) );
NAND2x1p5_ASAP7_75t_L g839 ( .A(n_732), .B(n_409), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_713), .Y(n_840) );
AOI21x1_ASAP7_75t_L g841 ( .A1(n_757), .A2(n_530), .B(n_529), .Y(n_841) );
AND2x2_ASAP7_75t_SL g842 ( .A(n_707), .B(n_538), .Y(n_842) );
AO21x2_ASAP7_75t_L g843 ( .A1(n_757), .A2(n_542), .B(n_541), .Y(n_843) );
INVx3_ASAP7_75t_L g844 ( .A(n_726), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_699), .Y(n_845) );
AO21x2_ASAP7_75t_L g846 ( .A1(n_767), .A2(n_613), .B(n_604), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_782), .A2(n_591), .B(n_613), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_745), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_721), .Y(n_849) );
AND2x4_ASAP7_75t_SL g850 ( .A(n_685), .B(n_613), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_686), .B(n_409), .Y(n_851) );
OAI21x1_ASAP7_75t_L g852 ( .A1(n_782), .A2(n_613), .B(n_453), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_695), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_773), .A2(n_613), .B(n_453), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_690), .Y(n_855) );
OA21x2_ASAP7_75t_L g856 ( .A1(n_741), .A2(n_438), .B(n_367), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_716), .A2(n_483), .B(n_468), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_717), .A2(n_508), .B(n_466), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_787), .B(n_510), .Y(n_859) );
INVx1_ASAP7_75t_SL g860 ( .A(n_721), .Y(n_860) );
AO21x2_ASAP7_75t_L g861 ( .A1(n_767), .A2(n_127), .B(n_125), .Y(n_861) );
AOI221x1_ASAP7_75t_L g862 ( .A1(n_791), .A2(n_511), .B1(n_510), .B2(n_13), .C(n_11), .Y(n_862) );
AOI21x1_ASAP7_75t_L g863 ( .A1(n_758), .A2(n_129), .B(n_128), .Y(n_863) );
INVx1_ASAP7_75t_SL g864 ( .A(n_690), .Y(n_864) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_732), .Y(n_865) );
OAI21x1_ASAP7_75t_L g866 ( .A1(n_691), .A2(n_135), .B(n_131), .Y(n_866) );
O2A1O1Ixp33_ASAP7_75t_L g867 ( .A1(n_702), .A2(n_14), .B(n_11), .C(n_12), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_695), .Y(n_868) );
INVx3_ASAP7_75t_L g869 ( .A(n_724), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_SL g870 ( .A1(n_791), .A2(n_138), .B(n_139), .C(n_136), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_777), .A2(n_19), .B1(n_17), .B2(n_18), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_788), .A2(n_21), .B1(n_17), .B2(n_20), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_714), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_732), .B(n_22), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_724), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_788), .B(n_23), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_691), .A2(n_145), .B(n_144), .Y(n_877) );
AO21x1_ASAP7_75t_L g878 ( .A1(n_747), .A2(n_149), .B(n_146), .Y(n_878) );
BUFx10_ASAP7_75t_L g879 ( .A(n_747), .Y(n_879) );
AO22x2_ASAP7_75t_L g880 ( .A1(n_729), .A2(n_756), .B1(n_743), .B2(n_715), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_777), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_714), .Y(n_882) );
NAND2xp33_ASAP7_75t_R g883 ( .A(n_731), .B(n_24), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_742), .Y(n_884) );
INVx8_ASAP7_75t_L g885 ( .A(n_724), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_703), .A2(n_154), .B(n_151), .Y(n_886) );
A2O1A1Ixp33_ASAP7_75t_L g887 ( .A1(n_733), .A2(n_29), .B(n_27), .C(n_28), .Y(n_887) );
OAI21x1_ASAP7_75t_L g888 ( .A1(n_703), .A2(n_158), .B(n_157), .Y(n_888) );
OA21x2_ASAP7_75t_L g889 ( .A1(n_765), .A2(n_160), .B(n_159), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_737), .B(n_27), .Y(n_890) );
OAI21xp5_ASAP7_75t_L g891 ( .A1(n_793), .A2(n_28), .B(n_29), .Y(n_891) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_728), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_697), .B(n_30), .Y(n_893) );
AOI22x1_ASAP7_75t_L g894 ( .A1(n_748), .A2(n_163), .B1(n_166), .B2(n_161), .Y(n_894) );
INVx4_ASAP7_75t_SL g895 ( .A(n_714), .Y(n_895) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_725), .A2(n_31), .B(n_33), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_728), .Y(n_897) );
OAI21x1_ASAP7_75t_L g898 ( .A1(n_712), .A2(n_172), .B(n_171), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_728), .Y(n_899) );
CKINVDCx11_ASAP7_75t_R g900 ( .A(n_735), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_761), .Y(n_901) );
NOR2x1_ASAP7_75t_SL g902 ( .A(n_735), .B(n_35), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_740), .Y(n_903) );
AO31x2_ASAP7_75t_L g904 ( .A1(n_748), .A2(n_38), .A3(n_36), .B(n_37), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_734), .B(n_36), .Y(n_905) );
AO31x2_ASAP7_75t_L g906 ( .A1(n_693), .A2(n_40), .A3(n_37), .B(n_39), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_789), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_698), .B(n_40), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_701), .B(n_41), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_712), .A2(n_174), .B(n_173), .Y(n_910) );
BUFx12f_ASAP7_75t_L g911 ( .A(n_754), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_792), .Y(n_912) );
OAI21x1_ASAP7_75t_L g913 ( .A1(n_720), .A2(n_177), .B(n_175), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_709), .A2(n_179), .B(n_178), .Y(n_914) );
AO21x1_ASAP7_75t_L g915 ( .A1(n_752), .A2(n_185), .B(n_181), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_760), .B(n_41), .Y(n_916) );
AOI222xp33_ASAP7_75t_L g917 ( .A1(n_738), .A2(n_43), .B1(n_44), .B2(n_45), .C1(n_46), .C2(n_47), .Y(n_917) );
OAI21x1_ASAP7_75t_L g918 ( .A1(n_720), .A2(n_187), .B(n_186), .Y(n_918) );
BUFx2_ASAP7_75t_L g919 ( .A(n_792), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_692), .B(n_43), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_739), .A2(n_44), .B1(n_46), .B2(n_49), .Y(n_921) );
OA21x2_ASAP7_75t_L g922 ( .A1(n_779), .A2(n_190), .B(n_188), .Y(n_922) );
OAI21x1_ASAP7_75t_L g923 ( .A1(n_784), .A2(n_193), .B(n_192), .Y(n_923) );
AND2x4_ASAP7_75t_L g924 ( .A(n_784), .B(n_50), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_792), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_739), .A2(n_50), .B1(n_51), .B2(n_52), .C(n_53), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_785), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_842), .A2(n_774), .B1(n_785), .B2(n_781), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_845), .B(n_746), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_802), .A2(n_808), .B(n_847), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_799), .B(n_783), .Y(n_931) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_883), .A2(n_776), .B1(n_770), .B2(n_763), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_827), .A2(n_769), .B1(n_778), .B2(n_770), .C(n_763), .Y(n_933) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_805), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_802), .A2(n_763), .B(n_745), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_880), .A2(n_778), .B1(n_56), .B2(n_57), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_811), .A2(n_195), .B(n_194), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g938 ( .A1(n_808), .A2(n_198), .B(n_196), .Y(n_938) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_903), .A2(n_55), .B(n_56), .C(n_58), .Y(n_939) );
BUFx3_ASAP7_75t_L g940 ( .A(n_801), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_817), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_852), .A2(n_201), .B(n_200), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_907), .B(n_62), .Y(n_943) );
AO31x2_ASAP7_75t_L g944 ( .A1(n_915), .A2(n_62), .A3(n_63), .B(n_64), .Y(n_944) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_811), .A2(n_64), .B(n_65), .Y(n_945) );
OAI22x1_ASAP7_75t_L g946 ( .A1(n_856), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_946) );
BUFx2_ASAP7_75t_L g947 ( .A(n_803), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_909), .Y(n_948) );
INVx11_ASAP7_75t_L g949 ( .A(n_911), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_800), .A2(n_204), .B(n_202), .Y(n_950) );
OAI21x1_ASAP7_75t_L g951 ( .A1(n_854), .A2(n_208), .B(n_207), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_880), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_817), .A2(n_68), .B1(n_70), .B2(n_71), .Y(n_953) );
OAI21xp5_ASAP7_75t_L g954 ( .A1(n_857), .A2(n_74), .B(n_75), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_824), .A2(n_77), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_836), .A2(n_80), .B1(n_81), .B2(n_83), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_909), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_836), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_818), .A2(n_86), .B1(n_87), .B2(n_91), .C(n_92), .Y(n_959) );
INVx11_ASAP7_75t_L g960 ( .A(n_900), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_893), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_908), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_917), .A2(n_94), .B(n_96), .C(n_97), .Y(n_963) );
BUFx2_ASAP7_75t_L g964 ( .A(n_828), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_815), .A2(n_101), .B1(n_103), .B2(n_104), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_795), .A2(n_105), .B(n_106), .C(n_107), .Y(n_966) );
INVx3_ASAP7_75t_L g967 ( .A(n_885), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_809), .B(n_108), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_871), .A2(n_110), .B1(n_113), .B2(n_114), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_840), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_833), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_971) );
AOI222xp33_ASAP7_75t_L g972 ( .A1(n_881), .A2(n_218), .B1(n_220), .B2(n_222), .C1(n_224), .C2(n_225), .Y(n_972) );
AOI211xp5_ASAP7_75t_L g973 ( .A1(n_881), .A2(n_226), .B(n_228), .C(n_229), .Y(n_973) );
BUFx6f_ASAP7_75t_L g974 ( .A(n_805), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_859), .B(n_230), .Y(n_975) );
OAI221xp5_ASAP7_75t_SL g976 ( .A1(n_926), .A2(n_234), .B1(n_235), .B2(n_239), .C(n_241), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_797), .A2(n_242), .B1(n_244), .B2(n_247), .Y(n_977) );
INVx1_ASAP7_75t_SL g978 ( .A(n_835), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g979 ( .A1(n_902), .A2(n_251), .B1(n_252), .B2(n_253), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_901), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_890), .A2(n_257), .B1(n_258), .B2(n_264), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g982 ( .A1(n_846), .A2(n_265), .B(n_266), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_872), .A2(n_268), .B1(n_272), .B2(n_276), .C(n_277), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_872), .A2(n_280), .B1(n_281), .B2(n_282), .Y(n_984) );
OAI21xp33_ASAP7_75t_SL g985 ( .A1(n_891), .A2(n_284), .B(n_285), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_920), .A2(n_286), .B1(n_287), .B2(n_288), .Y(n_986) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_796), .A2(n_289), .B(n_290), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_826), .B(n_292), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_916), .A2(n_295), .B1(n_297), .B2(n_298), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g990 ( .A1(n_857), .A2(n_301), .B1(n_303), .B2(n_305), .C(n_306), .Y(n_990) );
BUFx12f_ASAP7_75t_L g991 ( .A(n_831), .Y(n_991) );
INVx8_ASAP7_75t_L g992 ( .A(n_885), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_804), .A2(n_307), .B1(n_308), .B2(n_309), .C(n_313), .Y(n_993) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_804), .A2(n_314), .B1(n_315), .B2(n_316), .C(n_317), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_798), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_891), .A2(n_318), .B1(n_327), .B2(n_329), .C(n_330), .Y(n_996) );
OA21x2_ASAP7_75t_L g997 ( .A1(n_796), .A2(n_331), .B(n_333), .Y(n_997) );
BUFx6f_ASAP7_75t_L g998 ( .A(n_805), .Y(n_998) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_856), .A2(n_335), .B(n_336), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_905), .A2(n_884), .B1(n_896), .B2(n_876), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_865), .Y(n_1001) );
OAI211xp5_ASAP7_75t_SL g1002 ( .A1(n_867), .A2(n_339), .B(n_342), .C(n_343), .Y(n_1002) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_846), .A2(n_344), .B(n_345), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_810), .A2(n_346), .B1(n_347), .B2(n_350), .C(n_351), .Y(n_1004) );
AOI21xp5_ASAP7_75t_L g1005 ( .A1(n_807), .A2(n_355), .B(n_356), .Y(n_1005) );
OAI21x1_ASAP7_75t_L g1006 ( .A1(n_838), .A2(n_820), .B(n_816), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_813), .B(n_876), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_849), .A2(n_860), .B1(n_812), .B2(n_858), .Y(n_1008) );
OAI22xp5_ASAP7_75t_SL g1009 ( .A1(n_896), .A2(n_874), .B1(n_839), .B2(n_821), .Y(n_1009) );
NAND2xp5_ASAP7_75t_SL g1010 ( .A(n_849), .B(n_860), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_834), .B(n_858), .Y(n_1011) );
OAI211xp5_ASAP7_75t_L g1012 ( .A1(n_862), .A2(n_867), .B(n_921), .C(n_887), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_806), .B(n_895), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_834), .B(n_905), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_807), .A2(n_814), .B(n_812), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_819), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_839), .A2(n_821), .B1(n_850), .B2(n_924), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_830), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g1019 ( .A(n_848), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_806), .B(n_895), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_830), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_885), .Y(n_1022) );
AO21x1_ASAP7_75t_L g1023 ( .A1(n_924), .A2(n_863), .B(n_841), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_904), .Y(n_1024) );
AOI21x1_ASAP7_75t_L g1025 ( .A1(n_922), .A2(n_889), .B(n_829), .Y(n_1025) );
A2O1A1Ixp33_ASAP7_75t_L g1026 ( .A1(n_853), .A2(n_868), .B(n_832), .C(n_844), .Y(n_1026) );
OA21x2_ASAP7_75t_L g1027 ( .A1(n_866), .A2(n_888), .B(n_877), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_851), .A2(n_879), .B1(n_837), .B2(n_844), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_879), .A2(n_837), .B1(n_825), .B2(n_843), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_806), .A2(n_899), .B1(n_892), .B2(n_864), .Y(n_1030) );
AO31x2_ASAP7_75t_L g1031 ( .A1(n_878), .A2(n_912), .A3(n_925), .B(n_882), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_892), .B(n_899), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_822), .Y(n_1033) );
BUFx6f_ASAP7_75t_L g1034 ( .A(n_848), .Y(n_1034) );
INVx4_ASAP7_75t_L g1035 ( .A(n_806), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_822), .Y(n_1036) );
OAI222xp33_ASAP7_75t_L g1037 ( .A1(n_894), .A2(n_864), .B1(n_919), .B2(n_897), .C1(n_869), .C2(n_875), .Y(n_1037) );
NAND2xp33_ASAP7_75t_R g1038 ( .A(n_922), .B(n_889), .Y(n_1038) );
OAI21xp5_ASAP7_75t_L g1039 ( .A1(n_855), .A2(n_873), .B(n_927), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_870), .A2(n_823), .B1(n_843), .B2(n_897), .C(n_869), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_823), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_895), .B(n_875), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_848), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_886), .A2(n_910), .B(n_918), .Y(n_1044) );
OR2x6_ASAP7_75t_L g1045 ( .A(n_898), .B(n_913), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_914), .A2(n_904), .B1(n_906), .B2(n_861), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_906), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_970), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_948), .B(n_906), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_957), .B(n_923), .Y(n_1050) );
INVx3_ASAP7_75t_L g1051 ( .A(n_1013), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_1014), .A2(n_954), .B1(n_969), .B2(n_1009), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1018), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1021), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_942), .Y(n_1055) );
AO21x2_ASAP7_75t_L g1056 ( .A1(n_930), .A2(n_1015), .B(n_1025), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_980), .Y(n_1057) );
NOR2x1_ASAP7_75t_SL g1058 ( .A(n_1017), .B(n_1035), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_1045), .A2(n_1044), .B(n_1009), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_995), .B(n_929), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_978), .B(n_943), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_942), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_931), .Y(n_1063) );
NOR2x1_ASAP7_75t_L g1064 ( .A(n_1001), .B(n_1035), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_1013), .B(n_1020), .Y(n_1065) );
AO21x2_ASAP7_75t_L g1066 ( .A1(n_1047), .A2(n_1024), .B(n_945), .Y(n_1066) );
AOI322xp5_ASAP7_75t_L g1067 ( .A1(n_962), .A2(n_961), .A3(n_953), .B1(n_941), .B2(n_952), .C1(n_947), .C2(n_965), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1033), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_940), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_1043), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_992), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1016), .B(n_1011), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1036), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1000), .B(n_1007), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1041), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1000), .B(n_1032), .Y(n_1076) );
AND2x4_ASAP7_75t_L g1077 ( .A(n_1020), .B(n_1042), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1008), .B(n_1010), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_968), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_992), .Y(n_1080) );
INVx3_ASAP7_75t_L g1081 ( .A(n_934), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_946), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_934), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_934), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_984), .A2(n_956), .B1(n_958), .B2(n_959), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_988), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_974), .Y(n_1087) );
NOR4xp25_ASAP7_75t_SL g1088 ( .A(n_976), .B(n_1038), .C(n_955), .D(n_996), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_973), .B(n_975), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1022), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1028), .B(n_1030), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_974), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_960), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_973), .B(n_944), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_944), .B(n_939), .Y(n_1095) );
NAND2xp5_ASAP7_75t_SL g1096 ( .A(n_985), .B(n_932), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_974), .Y(n_1097) );
BUFx3_ASAP7_75t_L g1098 ( .A(n_967), .Y(n_1098) );
AO21x2_ASAP7_75t_L g1099 ( .A1(n_999), .A2(n_1023), .B(n_1005), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_944), .B(n_1042), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_984), .B(n_963), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_964), .B(n_967), .Y(n_1102) );
INVx3_ASAP7_75t_L g1103 ( .A(n_998), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_966), .Y(n_1104) );
INVx5_ASAP7_75t_L g1105 ( .A(n_1019), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1019), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_936), .B(n_972), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1019), .B(n_1034), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g1109 ( .A(n_1034), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1034), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_1039), .B(n_1026), .Y(n_1111) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_933), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_985), .B(n_1029), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1027), .Y(n_1114) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_949), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_991), .Y(n_1116) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_1045), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_951), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1045), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1012), .B(n_928), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1006), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_987), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_979), .B(n_983), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g1124 ( .A(n_987), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_982), .B(n_1003), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1031), .B(n_937), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g1127 ( .A(n_997), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1040), .B(n_989), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_937), .B(n_1031), .Y(n_1129) );
INVx3_ASAP7_75t_L g1130 ( .A(n_997), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1031), .B(n_971), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_938), .B(n_950), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_990), .A2(n_977), .B1(n_993), .B2(n_994), .Y(n_1133) );
INVx2_ASAP7_75t_L g1134 ( .A(n_981), .Y(n_1134) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_1037), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_935), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1004), .B(n_986), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1002), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1018), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_948), .B(n_957), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_948), .B(n_957), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_948), .B(n_957), .Y(n_1142) );
AO31x2_ASAP7_75t_L g1143 ( .A1(n_1046), .A2(n_1036), .A3(n_1041), .B(n_1033), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1048), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1049), .B(n_1074), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1053), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1053), .Y(n_1147) );
INVx3_ASAP7_75t_L g1148 ( .A(n_1109), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1049), .B(n_1074), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1076), .B(n_1100), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1054), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1057), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1140), .B(n_1141), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_1107), .A2(n_1101), .B1(n_1089), .B2(n_1085), .Y(n_1154) );
NAND2xp5_ASAP7_75t_SL g1155 ( .A(n_1089), .B(n_1052), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1076), .B(n_1100), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1142), .B(n_1060), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1078), .B(n_1139), .Y(n_1158) );
BUFx6f_ASAP7_75t_L g1159 ( .A(n_1109), .Y(n_1159) );
INVx3_ASAP7_75t_L g1160 ( .A(n_1109), .Y(n_1160) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_1080), .Y(n_1161) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_1105), .Y(n_1162) );
AO22x1_ASAP7_75t_L g1163 ( .A1(n_1064), .A2(n_1093), .B1(n_1065), .B2(n_1077), .Y(n_1163) );
AND2x4_ASAP7_75t_L g1164 ( .A(n_1119), .B(n_1117), .Y(n_1164) );
INVxp67_ASAP7_75t_L g1165 ( .A(n_1090), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1068), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1119), .B(n_1059), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1065), .B(n_1069), .Y(n_1168) );
OAI33xp33_ASAP7_75t_L g1169 ( .A1(n_1082), .A2(n_1104), .A3(n_1061), .B1(n_1120), .B2(n_1086), .B3(n_1079), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1072), .B(n_1063), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1070), .B(n_1102), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1073), .Y(n_1172) );
OAI31xp33_ASAP7_75t_SL g1173 ( .A1(n_1096), .A2(n_1113), .A3(n_1094), .B(n_1123), .Y(n_1173) );
OR2x6_ASAP7_75t_SL g1174 ( .A(n_1093), .B(n_1091), .Y(n_1174) );
INVx4_ASAP7_75t_L g1175 ( .A(n_1105), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1073), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1058), .B(n_1108), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1075), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1075), .B(n_1095), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1071), .B(n_1080), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1067), .B(n_1051), .Y(n_1181) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_1143), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_1143), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1051), .B(n_1098), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1114), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1098), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1050), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1050), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1112), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1095), .Y(n_1190) );
OAI211xp5_ASAP7_75t_SL g1191 ( .A1(n_1116), .A2(n_1115), .B(n_1128), .C(n_1138), .Y(n_1191) );
INVx2_ASAP7_75t_SL g1192 ( .A(n_1105), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1066), .B(n_1111), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1105), .B(n_1103), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1083), .B(n_1084), .Y(n_1195) );
AOI21xp5_ASAP7_75t_L g1196 ( .A1(n_1133), .A2(n_1134), .B(n_1088), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g1197 ( .A(n_1143), .Y(n_1197) );
NOR2x1_ASAP7_75t_SL g1198 ( .A(n_1135), .B(n_1092), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1143), .Y(n_1199) );
NAND2xp33_ASAP7_75t_SL g1200 ( .A(n_1134), .B(n_1137), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1185), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1145), .B(n_1149), .Y(n_1202) );
BUFx3_ASAP7_75t_L g1203 ( .A(n_1161), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_1155), .A2(n_1131), .B1(n_1132), .B2(n_1125), .Y(n_1204) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1185), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1145), .B(n_1056), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1166), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1166), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1172), .Y(n_1209) );
INVx3_ASAP7_75t_L g1210 ( .A(n_1177), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1150), .B(n_1156), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1150), .B(n_1129), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1156), .B(n_1129), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1158), .B(n_1129), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1176), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_1167), .B(n_1136), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1167), .B(n_1190), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1179), .B(n_1136), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1179), .B(n_1126), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1176), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1187), .B(n_1110), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1178), .Y(n_1222) );
INVx3_ASAP7_75t_L g1223 ( .A(n_1177), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1188), .B(n_1110), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1170), .B(n_1106), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1226 ( .A(n_1191), .B(n_1081), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1227 ( .A(n_1171), .B(n_1097), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1153), .B(n_1087), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1193), .B(n_1122), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1151), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1173), .B(n_1130), .Y(n_1231) );
INVx4_ASAP7_75t_L g1232 ( .A(n_1175), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1146), .Y(n_1233) );
INVx4_ASAP7_75t_L g1234 ( .A(n_1177), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1235 ( .A(n_1167), .B(n_1130), .Y(n_1235) );
OAI211xp5_ASAP7_75t_SL g1236 ( .A1(n_1165), .A2(n_1130), .B(n_1118), .C(n_1062), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_1147), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1157), .B(n_1099), .Y(n_1238) );
INVx3_ASAP7_75t_L g1239 ( .A(n_1159), .Y(n_1239) );
AOI211xp5_ASAP7_75t_SL g1240 ( .A1(n_1196), .A2(n_1055), .B(n_1062), .C(n_1121), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1217), .B(n_1164), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1202), .B(n_1168), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1206), .B(n_1183), .Y(n_1243) );
INVx3_ASAP7_75t_L g1244 ( .A(n_1234), .Y(n_1244) );
NOR2x1_ASAP7_75t_L g1245 ( .A(n_1232), .B(n_1180), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1206), .B(n_1197), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1211), .B(n_1154), .Y(n_1247) );
NAND2x1p5_ASAP7_75t_L g1248 ( .A(n_1232), .B(n_1162), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1228), .B(n_1152), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1225), .Y(n_1250) );
OAI21xp33_ASAP7_75t_L g1251 ( .A1(n_1231), .A2(n_1181), .B(n_1189), .Y(n_1251) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1217), .B(n_1164), .Y(n_1252) );
OR2x6_ASAP7_75t_L g1253 ( .A(n_1234), .B(n_1163), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1201), .Y(n_1254) );
INVx5_ASAP7_75t_L g1255 ( .A(n_1232), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1205), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1230), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1212), .B(n_1174), .Y(n_1258) );
NAND2x1p5_ASAP7_75t_L g1259 ( .A(n_1203), .B(n_1162), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1219), .B(n_1183), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1213), .B(n_1182), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1227), .B(n_1144), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_1237), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1214), .B(n_1199), .Y(n_1264) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_1251), .A2(n_1169), .B1(n_1200), .B2(n_1238), .C(n_1204), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1249), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1267 ( .A1(n_1245), .A2(n_1200), .B1(n_1217), .B2(n_1226), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_1244), .B(n_1210), .Y(n_1268) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_1255), .A2(n_1223), .B1(n_1210), .B2(n_1203), .Y(n_1269) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1263), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1250), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1257), .Y(n_1272) );
AND4x1_ASAP7_75t_L g1273 ( .A(n_1258), .B(n_1240), .C(n_1184), .D(n_1194), .Y(n_1273) );
INVx3_ASAP7_75t_L g1274 ( .A(n_1255), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1243), .B(n_1218), .Y(n_1275) );
O2A1O1Ixp33_ASAP7_75t_SL g1276 ( .A1(n_1244), .A2(n_1223), .B(n_1192), .C(n_1186), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1243), .B(n_1218), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1246), .B(n_1224), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1242), .B(n_1229), .Y(n_1279) );
OAI22xp33_ASAP7_75t_L g1280 ( .A1(n_1267), .A2(n_1253), .B1(n_1244), .B2(n_1248), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1272), .Y(n_1281) );
INVx1_ASAP7_75t_SL g1282 ( .A(n_1279), .Y(n_1282) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1270), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1266), .B(n_1247), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1271), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1278), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1274), .Y(n_1287) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1274), .Y(n_1288) );
XNOR2xp5_ASAP7_75t_L g1289 ( .A(n_1273), .B(n_1262), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1275), .B(n_1277), .Y(n_1290) );
AOI211xp5_ASAP7_75t_L g1291 ( .A1(n_1280), .A2(n_1276), .B(n_1269), .C(n_1265), .Y(n_1291) );
BUFx4f_ASAP7_75t_SL g1292 ( .A(n_1282), .Y(n_1292) );
INVx5_ASAP7_75t_L g1293 ( .A(n_1287), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1284), .B(n_1260), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1284), .B(n_1261), .Y(n_1295) );
AOI21xp5_ASAP7_75t_L g1296 ( .A1(n_1289), .A2(n_1268), .B(n_1259), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1281), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_1290), .A2(n_1252), .B1(n_1241), .B2(n_1264), .Y(n_1298) );
NAND4xp25_ASAP7_75t_SL g1299 ( .A(n_1291), .B(n_1286), .C(n_1290), .D(n_1288), .Y(n_1299) );
NOR3xp33_ASAP7_75t_SL g1300 ( .A(n_1296), .B(n_1236), .C(n_1285), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1297), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_1292), .A2(n_1283), .B1(n_1235), .B2(n_1229), .Y(n_1302) );
AOI221xp5_ASAP7_75t_L g1303 ( .A1(n_1298), .A2(n_1221), .B1(n_1216), .B2(n_1235), .C(n_1256), .Y(n_1303) );
NAND4xp25_ASAP7_75t_L g1304 ( .A(n_1294), .B(n_1235), .C(n_1216), .D(n_1239), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1305 ( .A(n_1301), .Y(n_1305) );
OAI21xp5_ASAP7_75t_L g1306 ( .A1(n_1299), .A2(n_1293), .B(n_1295), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1302), .Y(n_1307) );
NOR3xp33_ASAP7_75t_SL g1308 ( .A(n_1304), .B(n_1209), .C(n_1233), .Y(n_1308) );
INVxp67_ASAP7_75t_SL g1309 ( .A(n_1305), .Y(n_1309) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_1307), .B(n_1300), .C(n_1303), .Y(n_1310) );
NAND3x1_ASAP7_75t_L g1311 ( .A(n_1306), .B(n_1239), .C(n_1148), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1309), .Y(n_1312) );
AO21x2_ASAP7_75t_L g1313 ( .A1(n_1310), .A2(n_1308), .B(n_1198), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1311), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1312), .Y(n_1315) );
OAI21x1_ASAP7_75t_L g1316 ( .A1(n_1315), .A2(n_1314), .B(n_1313), .Y(n_1316) );
AOI22x1_ASAP7_75t_L g1317 ( .A1(n_1316), .A2(n_1160), .B1(n_1159), .B2(n_1254), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_1317), .A2(n_1195), .B1(n_1127), .B2(n_1124), .Y(n_1318) );
AOI222xp33_ASAP7_75t_L g1319 ( .A1(n_1318), .A2(n_1207), .B1(n_1222), .B2(n_1220), .C1(n_1215), .C2(n_1208), .Y(n_1319) );
endmodule