module real_aes_8433_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_0), .A2(n_26), .B1(n_164), .B2(n_167), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_SL g322 ( .A1(n_1), .A2(n_323), .B(n_324), .C(n_328), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_2), .B(n_265), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_3), .B(n_237), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_4), .A2(n_219), .B(n_256), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_5), .Y(n_106) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_6), .A2(n_253), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g209 ( .A(n_7), .Y(n_209) );
AND2x6_ASAP7_75t_L g224 ( .A(n_7), .B(n_207), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_7), .B(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_8), .A2(n_13), .B1(n_154), .B2(n_159), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_9), .A2(n_189), .B1(n_192), .B2(n_193), .Y(n_188) );
INVx1_ASAP7_75t_L g192 ( .A(n_9), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_9), .A2(n_224), .B(n_228), .C(n_338), .Y(n_337) );
AO22x2_ASAP7_75t_L g87 ( .A1(n_10), .A2(n_22), .B1(n_88), .B2(n_89), .Y(n_87) );
INVx1_ASAP7_75t_L g247 ( .A(n_11), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_12), .B(n_237), .Y(n_275) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_14), .A2(n_25), .B1(n_88), .B2(n_92), .Y(n_91) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_15), .A2(n_228), .B(n_279), .C(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_16), .A2(n_81), .B1(n_179), .B2(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_16), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_17), .A2(n_228), .B(n_272), .C(n_279), .Y(n_271) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_18), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_19), .A2(n_81), .B1(n_178), .B2(n_179), .Y(n_80) );
INVx1_ASAP7_75t_L g178 ( .A(n_19), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_20), .A2(n_219), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g222 ( .A(n_21), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_23), .A2(n_226), .B(n_241), .C(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_SL g544 ( .A1(n_23), .A2(n_81), .B1(n_179), .B2(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_23), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_24), .A2(n_37), .B1(n_142), .B2(n_146), .Y(n_141) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_25), .A2(n_42), .B1(n_55), .B2(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_25), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_27), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_28), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_29), .B(n_296), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_30), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_31), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_32), .B(n_219), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_33), .A2(n_66), .B1(n_171), .B2(n_175), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_34), .A2(n_226), .B(n_231), .C(n_241), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_35), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g325 ( .A(n_36), .Y(n_325) );
INVx1_ASAP7_75t_L g232 ( .A(n_38), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_39), .B(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_40), .Y(n_305) );
OAI22xp5_ASAP7_75t_SL g189 ( .A1(n_41), .A2(n_61), .B1(n_190), .B2(n_191), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_41), .Y(n_191) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_42), .A2(n_64), .B1(n_88), .B2(n_92), .Y(n_95) );
INVxp67_ASAP7_75t_L g204 ( .A(n_42), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
INVx1_ASAP7_75t_L g207 ( .A(n_44), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_45), .B(n_219), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_46), .B(n_265), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_47), .A2(n_259), .B(n_261), .C(n_263), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_L g246 ( .A(n_49), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_50), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_51), .B(n_237), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_52), .B(n_238), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_53), .Y(n_113) );
INVx1_ASAP7_75t_L g195 ( .A(n_54), .Y(n_195) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_55), .A2(n_70), .B1(n_88), .B2(n_89), .Y(n_97) );
OAI22xp5_ASAP7_75t_SL g184 ( .A1(n_56), .A2(n_62), .B1(n_185), .B2(n_186), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_56), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_57), .B(n_234), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_58), .A2(n_228), .B(n_241), .C(n_311), .Y(n_310) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_59), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_60), .B(n_233), .Y(n_300) );
INVx1_ASAP7_75t_L g190 ( .A(n_61), .Y(n_190) );
INVx1_ASAP7_75t_L g186 ( .A(n_62), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_63), .Y(n_291) );
INVx2_ASAP7_75t_L g244 ( .A(n_65), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_67), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_68), .B(n_327), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_69), .B(n_219), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_71), .Y(n_288) );
INVxp67_ASAP7_75t_L g262 ( .A(n_72), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_73), .Y(n_98) );
INVx1_ASAP7_75t_L g88 ( .A(n_74), .Y(n_88) );
INVx1_ASAP7_75t_L g90 ( .A(n_74), .Y(n_90) );
INVx1_ASAP7_75t_L g312 ( .A(n_75), .Y(n_312) );
INVx1_ASAP7_75t_L g335 ( .A(n_76), .Y(n_335) );
AND2x2_ASAP7_75t_L g248 ( .A(n_77), .B(n_243), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_197), .B1(n_210), .B2(n_540), .C(n_543), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_180), .Y(n_79) );
INVx2_ASAP7_75t_SL g179 ( .A(n_81), .Y(n_179) );
AND2x4_ASAP7_75t_L g81 ( .A(n_82), .B(n_139), .Y(n_81) );
NOR3xp33_ASAP7_75t_SL g82 ( .A(n_83), .B(n_112), .C(n_125), .Y(n_82) );
OAI221xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_98), .B1(n_99), .B2(n_106), .C(n_107), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AND2x6_ASAP7_75t_L g85 ( .A(n_86), .B(n_93), .Y(n_85) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_91), .Y(n_86) );
AND2x2_ASAP7_75t_L g105 ( .A(n_87), .B(n_95), .Y(n_105) );
INVx2_ASAP7_75t_L g117 ( .A(n_87), .Y(n_117) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g92 ( .A(n_90), .Y(n_92) );
INVx2_ASAP7_75t_L g104 ( .A(n_91), .Y(n_104) );
OR2x2_ASAP7_75t_L g116 ( .A(n_91), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g124 ( .A(n_91), .B(n_117), .Y(n_124) );
INVx1_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
AND2x6_ASAP7_75t_L g144 ( .A(n_93), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g166 ( .A(n_93), .B(n_152), .Y(n_166) );
AND2x4_ASAP7_75t_L g174 ( .A(n_93), .B(n_124), .Y(n_174) );
AND2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_96), .Y(n_93) );
AND2x2_ASAP7_75t_L g119 ( .A(n_94), .B(n_97), .Y(n_119) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_95), .B(n_97), .Y(n_151) );
AND2x2_ASAP7_75t_L g158 ( .A(n_95), .B(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g103 ( .A(n_97), .Y(n_103) );
INVx1_ASAP7_75t_L g138 ( .A(n_97), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_100), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
INVx1_ASAP7_75t_L g111 ( .A(n_103), .Y(n_111) );
INVx1_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
AND2x2_ASAP7_75t_L g152 ( .A(n_104), .B(n_117), .Y(n_152) );
AND2x4_ASAP7_75t_L g110 ( .A(n_105), .B(n_111), .Y(n_110) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_105), .B(n_130), .Y(n_129) );
BUFx4f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_114), .B1(n_120), .B2(n_121), .Y(n_112) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx2_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g123 ( .A(n_119), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g169 ( .A(n_119), .B(n_152), .Y(n_169) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g157 ( .A(n_124), .B(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_131), .B2(n_132), .Y(n_125) );
INVx3_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
CKINVDCx16_ASAP7_75t_R g133 ( .A(n_134), .Y(n_133) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_162), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_153), .Y(n_140) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
INVx11_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x6_ASAP7_75t_L g160 ( .A(n_151), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g177 ( .A(n_152), .B(n_158), .Y(n_177) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx8_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_170), .Y(n_162) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_182), .B1(n_194), .B2(n_196), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_187), .B2(n_188), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_185), .A2(n_227), .B(n_242), .C(n_322), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g193 ( .A(n_189), .Y(n_193) );
INVx1_ASAP7_75t_L g196 ( .A(n_194), .Y(n_196) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
AND3x1_ASAP7_75t_SL g199 ( .A(n_200), .B(n_205), .C(n_208), .Y(n_199) );
INVxp67_ASAP7_75t_L g549 ( .A(n_200), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_205), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_205), .A2(n_228), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g559 ( .A(n_205), .Y(n_559) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_206), .B(n_209), .Y(n_553) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_SL g558 ( .A(n_208), .B(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR5x1_ASAP7_75t_L g213 ( .A(n_214), .B(n_413), .C(n_491), .D(n_515), .E(n_532), .Y(n_213) );
OAI211xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_280), .B(n_330), .C(n_390), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_249), .Y(n_215) );
AND2x2_ASAP7_75t_L g344 ( .A(n_216), .B(n_251), .Y(n_344) );
INVx5_ASAP7_75t_SL g372 ( .A(n_216), .Y(n_372) );
AND2x2_ASAP7_75t_L g408 ( .A(n_216), .B(n_393), .Y(n_408) );
OR2x2_ASAP7_75t_L g447 ( .A(n_216), .B(n_250), .Y(n_447) );
OR2x2_ASAP7_75t_L g478 ( .A(n_216), .B(n_369), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_216), .B(n_382), .Y(n_514) );
AND2x2_ASAP7_75t_L g526 ( .A(n_216), .B(n_369), .Y(n_526) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_248), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_225), .B(n_243), .Y(n_217) );
BUFx2_ASAP7_75t_L g296 ( .A(n_219), .Y(n_296) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_220), .B(n_224), .Y(n_336) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g263 ( .A(n_221), .Y(n_263) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g229 ( .A(n_222), .Y(n_229) );
INVx1_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g230 ( .A(n_223), .Y(n_230) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
INVx3_ASAP7_75t_L g238 ( .A(n_223), .Y(n_238) );
INVx1_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_223), .Y(n_327) );
INVx4_ASAP7_75t_SL g242 ( .A(n_224), .Y(n_242) );
BUFx3_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_242), .B(n_257), .C(n_258), .Y(n_256) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g542 ( .A(n_228), .B(n_279), .Y(n_542) );
AND2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
BUFx3_ASAP7_75t_L g240 ( .A(n_229), .Y(n_240) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_229), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_236), .C(n_239), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_233), .A2(n_239), .B(n_288), .C(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g260 ( .A(n_235), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_237), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g323 ( .A(n_237), .Y(n_323) );
INVx5_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g328 ( .A(n_240), .Y(n_328) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_243), .A2(n_285), .B(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_243), .Y(n_306) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g254 ( .A(n_244), .B(n_245), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g525 ( .A(n_249), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g388 ( .A(n_250), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_267), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_251), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_251), .Y(n_381) );
INVx3_ASAP7_75t_L g396 ( .A(n_251), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_251), .B(n_267), .Y(n_420) );
OR2x2_ASAP7_75t_L g429 ( .A(n_251), .B(n_372), .Y(n_429) );
AND2x2_ASAP7_75t_L g433 ( .A(n_251), .B(n_393), .Y(n_433) );
AND2x2_ASAP7_75t_L g439 ( .A(n_251), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g476 ( .A(n_251), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_251), .B(n_333), .Y(n_490) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_255), .B(n_264), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx4_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_253), .A2(n_270), .B(n_271), .Y(n_269) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g343 ( .A(n_254), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_259), .A2(n_312), .B(n_313), .C(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
OA21x2_ASAP7_75t_L g319 ( .A1(n_265), .A2(n_320), .B(n_329), .Y(n_319) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_266), .B(n_291), .Y(n_290) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_266), .A2(n_309), .B(n_317), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_266), .B(n_318), .Y(n_317) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_266), .A2(n_334), .B(n_341), .Y(n_333) );
OR2x2_ASAP7_75t_L g382 ( .A(n_267), .B(n_333), .Y(n_382) );
AND2x2_ASAP7_75t_L g393 ( .A(n_267), .B(n_369), .Y(n_393) );
AND2x2_ASAP7_75t_L g405 ( .A(n_267), .B(n_396), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_267), .B(n_333), .Y(n_428) );
INVx1_ASAP7_75t_SL g440 ( .A(n_267), .Y(n_440) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g332 ( .A(n_268), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_268), .B(n_372), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_276), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_276), .A2(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_292), .Y(n_281) );
AND2x2_ASAP7_75t_L g353 ( .A(n_282), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_282), .B(n_307), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_282), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_282), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g385 ( .A(n_282), .B(n_376), .Y(n_385) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_282), .Y(n_404) );
AND2x2_ASAP7_75t_L g425 ( .A(n_282), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g435 ( .A(n_282), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g481 ( .A(n_282), .B(n_364), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_282), .B(n_387), .Y(n_508) );
INVx5_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g378 ( .A(n_283), .Y(n_378) );
AND2x2_ASAP7_75t_L g444 ( .A(n_283), .B(n_376), .Y(n_444) );
AND2x2_ASAP7_75t_L g528 ( .A(n_283), .B(n_396), .Y(n_528) );
OR2x6_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_292), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g517 ( .A(n_292), .Y(n_517) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_307), .Y(n_292) );
AND2x2_ASAP7_75t_L g347 ( .A(n_293), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g356 ( .A(n_293), .B(n_354), .Y(n_356) );
INVx5_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
AND2x2_ASAP7_75t_L g387 ( .A(n_293), .B(n_319), .Y(n_387) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_293), .Y(n_424) );
OR2x6_ASAP7_75t_L g293 ( .A(n_294), .B(n_304), .Y(n_293) );
AOI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_302), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g465 ( .A(n_307), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_307), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g498 ( .A(n_307), .B(n_364), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_307), .A2(n_421), .B(n_528), .C(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_319), .Y(n_307) );
BUFx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
INVx2_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_316), .Y(n_309) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_319), .B(n_352), .Y(n_361) );
AND2x2_ASAP7_75t_L g452 ( .A(n_319), .B(n_364), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI211x1_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_345), .B(n_358), .C(n_383), .Y(n_330) );
INVx1_ASAP7_75t_L g449 ( .A(n_331), .Y(n_449) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_344), .Y(n_331) );
INVx5_ASAP7_75t_SL g369 ( .A(n_333), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_333), .B(n_439), .Y(n_438) );
AOI311xp33_ASAP7_75t_L g457 ( .A1(n_333), .A2(n_458), .A3(n_460), .B(n_461), .C(n_467), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_333), .A2(n_405), .B(n_493), .C(n_496), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_337), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVxp67_ASAP7_75t_L g412 ( .A(n_344), .Y(n_412) );
NAND4xp25_ASAP7_75t_SL g345 ( .A(n_346), .B(n_349), .C(n_355), .D(n_357), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_346), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g403 ( .A(n_347), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_350), .B(n_356), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_350), .B(n_363), .Y(n_483) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_351), .B(n_364), .Y(n_501) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g376 ( .A(n_352), .Y(n_376) );
INVxp67_ASAP7_75t_L g411 ( .A(n_353), .Y(n_411) );
AND2x4_ASAP7_75t_L g363 ( .A(n_354), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g437 ( .A(n_354), .B(n_376), .Y(n_437) );
INVx1_ASAP7_75t_L g464 ( .A(n_354), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_354), .B(n_451), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_355), .B(n_425), .Y(n_445) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_356), .B(n_378), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_356), .B(n_425), .Y(n_524) );
INVx1_ASAP7_75t_L g535 ( .A(n_357), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_365), .C(n_373), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g377 ( .A(n_361), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g415 ( .A(n_361), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
AND2x2_ASAP7_75t_L g374 ( .A(n_363), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_363), .B(n_425), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_363), .B(n_444), .Y(n_468) );
OR2x2_ASAP7_75t_L g384 ( .A(n_364), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g416 ( .A(n_364), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_364), .B(n_376), .Y(n_431) );
AND2x2_ASAP7_75t_L g488 ( .A(n_364), .B(n_444), .Y(n_488) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_364), .Y(n_495) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_366), .A2(n_378), .B1(n_500), .B2(n_502), .C(n_505), .Y(n_499) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g389 ( .A(n_369), .B(n_372), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_369), .B(n_439), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_369), .B(n_396), .Y(n_504) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g489 ( .A(n_371), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g503 ( .A(n_371), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_372), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_372), .B(n_393), .Y(n_400) );
AND2x2_ASAP7_75t_L g470 ( .A(n_372), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_372), .B(n_419), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_372), .B(n_520), .Y(n_519) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_377), .B(n_379), .Y(n_373) );
INVx2_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
OR2x2_ASAP7_75t_L g430 ( .A(n_378), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g533 ( .A(n_378), .B(n_501), .Y(n_533) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g537 ( .A(n_384), .Y(n_537) );
INVx2_ASAP7_75t_SL g451 ( .A(n_385), .Y(n_451) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_388), .A2(n_469), .B(n_533), .C(n_534), .Y(n_532) );
OAI322xp33_ASAP7_75t_SL g401 ( .A1(n_389), .A2(n_402), .A3(n_405), .B1(n_406), .B2(n_407), .C1(n_409), .C2(n_412), .Y(n_401) );
INVx2_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_401), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI22xp33_ASAP7_75t_SL g467 ( .A1(n_392), .A2(n_468), .B1(n_469), .B2(n_472), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_393), .B(n_396), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_393), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g466 ( .A(n_395), .B(n_428), .Y(n_466) );
INVx1_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_400), .A2(n_510), .B(n_512), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_402), .A2(n_435), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp67_ASAP7_75t_SL g463 ( .A(n_404), .B(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_404), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g520 ( .A(n_405), .Y(n_520) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_441), .C(n_457), .D(n_473), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_422), .C(n_434), .Y(n_414) );
INVx1_ASAP7_75t_L g506 ( .A(n_415), .Y(n_506) );
AND2x2_ASAP7_75t_L g454 ( .A(n_416), .B(n_437), .Y(n_454) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_421), .B(n_456), .Y(n_455) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B1(n_430), .B2(n_432), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_424), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_425), .A2(n_464), .B(n_487), .C(n_489), .Y(n_486) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
INVx1_ASAP7_75t_L g531 ( .A(n_429), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g521 ( .A(n_430), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g460 ( .A(n_439), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B(n_446), .C(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_453), .B2(n_455), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_451), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_456), .B(n_477), .Y(n_539) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI21xp33_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_465), .B(n_466), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_479), .B1(n_482), .B2(n_484), .C(n_486), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_489), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_505) );
NAND3xp33_ASAP7_75t_SL g491 ( .A(n_492), .B(n_499), .C(n_509), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI211xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .C(n_527), .Y(n_515) );
INVx1_ASAP7_75t_L g536 ( .A(n_516), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .B1(n_523), .B2(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_537), .B2(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .A3(n_546), .B1(n_550), .B2(n_551), .C1(n_554), .C2(n_556), .Y(n_543) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
endmodule