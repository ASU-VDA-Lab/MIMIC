module fake_jpeg_7330_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.C(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_1),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_20),
.B1(n_17),
.B2(n_11),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_28),
.B1(n_15),
.B2(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_12),
.B1(n_15),
.B2(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_27),
.B(n_23),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_1),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_24),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_9),
.B(n_25),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_9),
.B1(n_16),
.B2(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_47),
.Y(n_54)
);

XOR2x2_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_31),
.Y(n_44)
);

A2O1A1O1Ixp25_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_2),
.B(n_3),
.C(n_5),
.D(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_49),
.B1(n_42),
.B2(n_41),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_44),
.B(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_37),
.C(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

NAND4xp25_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_9),
.C(n_16),
.D(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_2),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_62),
.B(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_57),
.B(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_55),
.B2(n_3),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_16),
.Y(n_69)
);


endmodule