module fake_netlist_5_80_n_1102 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1102);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1102;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_969;
wire n_866;
wire n_236;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_1094;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_639;
wire n_914;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_110),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_128),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_6),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_16),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_36),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_95),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_49),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_77),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_59),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_101),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_32),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_113),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_71),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_75),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_33),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_108),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_142),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_124),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_125),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_15),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_105),
.Y(n_251)
);

HB1xp67_ASAP7_75t_SL g252 ( 
.A(n_147),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_12),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_149),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_67),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_157),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_23),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

CKINVDCx6p67_ASAP7_75t_R g267 ( 
.A(n_104),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_215),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_231),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_240),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_235),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_260),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_260),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_207),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_224),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_207),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_207),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_210),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_259),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_196),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_223),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_267),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_248),
.B(n_223),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_312),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_271),
.A2(n_227),
.B1(n_211),
.B2(n_222),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_223),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_271),
.A2(n_200),
.B1(n_221),
.B2(n_263),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_276),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

AOI22x1_ASAP7_75t_SL g346 ( 
.A1(n_282),
.A2(n_265),
.B1(n_264),
.B2(n_257),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_198),
.B(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_280),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_248),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_199),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_286),
.B(n_201),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_272),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_273),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_202),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_293),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_292),
.B(n_223),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_208),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_294),
.B(n_248),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_209),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_R g373 ( 
.A(n_334),
.B(n_296),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_342),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_212),
.Y(n_375)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_310),
.B(n_297),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_R g378 ( 
.A(n_334),
.B(n_306),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_364),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_R g382 ( 
.A(n_358),
.B(n_306),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_358),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_336),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_328),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_328),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_329),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_329),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_350),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_346),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

OA22x2_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_314),
.B1(n_237),
.B2(n_246),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_346),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_320),
.B(n_287),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_339),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_341),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_332),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_351),
.B(n_293),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

AND3x2_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_0),
.C(n_1),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_357),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_363),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_370),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_322),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_327),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_327),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_327),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_349),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_365),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_359),
.B(n_300),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_365),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_337),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_337),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_337),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_319),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_367),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_R g438 ( 
.A(n_359),
.B(n_300),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_367),
.B(n_214),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_347),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_353),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_367),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_367),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_369),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_345),
.B(n_219),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_347),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_347),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_347),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_248),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_302),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_226),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_229),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_383),
.B(n_302),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_371),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_413),
.B(n_319),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_359),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_418),
.B(n_230),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_L g469 ( 
.A1(n_397),
.A2(n_371),
.B1(n_369),
.B2(n_348),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_368),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_434),
.B(n_325),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_374),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_421),
.B(n_232),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_415),
.B(n_236),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_419),
.B(n_238),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_431),
.B(n_239),
.Y(n_482)
);

AND2x2_ASAP7_75t_SL g483 ( 
.A(n_410),
.B(n_325),
.Y(n_483)
);

NOR2x1p5_ASAP7_75t_L g484 ( 
.A(n_422),
.B(n_241),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_412),
.B(n_333),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_438),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_375),
.B(n_368),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_321),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_392),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_368),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_403),
.B(n_279),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_318),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_403),
.B(n_385),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_373),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_433),
.B(n_344),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_321),
.Y(n_504)
);

CKINVDCx11_ASAP7_75t_R g505 ( 
.A(n_374),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_437),
.B(n_442),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_423),
.B(n_318),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_376),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_380),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_440),
.B(n_242),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_386),
.B(n_279),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_387),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_440),
.B(n_447),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_445),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_447),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_439),
.B(n_344),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_384),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_384),
.B(n_244),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_446),
.B(n_318),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_378),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_382),
.B(n_348),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_461),
.B(n_325),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_524),
.A2(n_521),
.B1(n_523),
.B2(n_483),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_461),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_449),
.A2(n_395),
.B(n_391),
.C(n_338),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

BUFx8_ASAP7_75t_L g538 ( 
.A(n_531),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_503),
.B(n_390),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_505),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_338),
.B1(n_343),
.B2(n_331),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_511),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_483),
.B(n_345),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_511),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_472),
.B(n_345),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_343),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

BUFx8_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_466),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_490),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_472),
.B(n_345),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_490),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_503),
.B(n_34),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_449),
.B(n_345),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_476),
.B(n_35),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_478),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_2),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_497),
.B(n_40),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_497),
.B(n_41),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_493),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_331),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_456),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_528),
.B(n_3),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_513),
.A2(n_331),
.B1(n_330),
.B2(n_345),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_462),
.B(n_352),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_471),
.B(n_333),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_508),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_473),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_498),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_43),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_520),
.B(n_330),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_499),
.Y(n_587)
);

AOI211xp5_ASAP7_75t_L g588 ( 
.A1(n_527),
.A2(n_479),
.B(n_453),
.C(n_516),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_514),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_512),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_519),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_522),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_509),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_352),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_588),
.B(n_458),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_479),
.Y(n_601)
);

INVx11_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_556),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_572),
.B(n_453),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_571),
.A2(n_487),
.B(n_492),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_571),
.A2(n_510),
.B(n_529),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_560),
.A2(n_510),
.B(n_513),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_541),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_480),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_555),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_566),
.B(n_480),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_535),
.A2(n_560),
.B(n_546),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_553),
.B(n_517),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_566),
.B(n_458),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_543),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_SL g620 ( 
.A(n_598),
.B(n_515),
.Y(n_620)
);

AOI21xp33_ASAP7_75t_L g621 ( 
.A1(n_573),
.A2(n_454),
.B(n_482),
.Y(n_621)
);

O2A1O1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_573),
.A2(n_536),
.B(n_534),
.C(n_450),
.Y(n_622)
);

AO32x2_ASAP7_75t_L g623 ( 
.A1(n_534),
.A2(n_518),
.A3(n_486),
.B1(n_469),
.B2(n_450),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_591),
.Y(n_624)
);

AO22x1_ASAP7_75t_L g625 ( 
.A1(n_539),
.A2(n_526),
.B1(n_530),
.B2(n_502),
.Y(n_625)
);

NOR2x1_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_452),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_559),
.B(n_525),
.Y(n_627)
);

OAI321xp33_ASAP7_75t_L g628 ( 
.A1(n_547),
.A2(n_482),
.A3(n_467),
.B1(n_477),
.B2(n_485),
.C(n_7),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_535),
.A2(n_520),
.B1(n_525),
.B2(n_467),
.Y(n_629)
);

O2A1O1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_536),
.A2(n_477),
.B(n_507),
.C(n_484),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_543),
.B(n_520),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_569),
.Y(n_632)
);

CKINVDCx10_ASAP7_75t_R g633 ( 
.A(n_538),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_457),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_592),
.B(n_455),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_457),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_546),
.A2(n_468),
.B(n_330),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_565),
.A2(n_518),
.B(n_457),
.C(n_5),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_578),
.A2(n_468),
.B(n_330),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_567),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_539),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_587),
.B(n_505),
.Y(n_644)
);

O2A1O1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_594),
.A2(n_457),
.B(n_4),
.C(n_5),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_568),
.B(n_457),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_468),
.Y(n_647)
);

AOI22x1_ASAP7_75t_L g648 ( 
.A1(n_597),
.A2(n_504),
.B1(n_488),
.B2(n_330),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_568),
.B(n_468),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_548),
.B(n_488),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_SL g651 ( 
.A1(n_599),
.A2(n_504),
.B(n_488),
.C(n_102),
.Y(n_651)
);

OAI21xp33_ASAP7_75t_L g652 ( 
.A1(n_582),
.A2(n_3),
.B(n_4),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_595),
.B(n_488),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_550),
.B(n_488),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_504),
.C(n_6),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_578),
.A2(n_352),
.B(n_504),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_599),
.A2(n_504),
.B(n_352),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_641),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_615),
.A2(n_557),
.B1(n_548),
.B2(n_563),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_605),
.A2(n_576),
.B(n_533),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_601),
.B(n_552),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_611),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_614),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_617),
.B(n_563),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_641),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_631),
.B(n_593),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_604),
.B(n_552),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_641),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_612),
.B(n_577),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_627),
.A2(n_557),
.B1(n_581),
.B2(n_583),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_622),
.A2(n_586),
.B(n_576),
.C(n_589),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_SL g673 ( 
.A1(n_642),
.A2(n_550),
.B1(n_537),
.B2(n_540),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_606),
.A2(n_533),
.B(n_585),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_642),
.A2(n_550),
.B1(n_542),
.B2(n_584),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_550),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_621),
.A2(n_590),
.B(n_580),
.C(n_545),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_643),
.B(n_618),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_619),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_624),
.B(n_549),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_628),
.B(n_570),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_616),
.A2(n_585),
.B(n_579),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_643),
.B(n_550),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_607),
.A2(n_574),
.B(n_542),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_603),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_628),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_630),
.A2(n_575),
.B(n_352),
.C(n_10),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_610),
.B(n_44),
.Y(n_689)
);

AOI21x1_ASAP7_75t_L g690 ( 
.A1(n_640),
.A2(n_352),
.B(n_46),
.Y(n_690)
);

AO21x2_ASAP7_75t_L g691 ( 
.A1(n_607),
.A2(n_47),
.B(n_45),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_644),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_600),
.B(n_8),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_609),
.B(n_50),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_636),
.B(n_9),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_652),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_639),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_629),
.B(n_14),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_609),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_609),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_SL g702 ( 
.A(n_646),
.B(n_18),
.Y(n_702)
);

AO21x2_ASAP7_75t_L g703 ( 
.A1(n_657),
.A2(n_120),
.B(n_195),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_625),
.B(n_19),
.C(n_20),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_SL g705 ( 
.A(n_655),
.B(n_19),
.C(n_20),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_602),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_650),
.A2(n_122),
.B(n_194),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_632),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_623),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_626),
.B(n_647),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_649),
.B(n_21),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_634),
.A2(n_637),
.B1(n_653),
.B2(n_654),
.Y(n_712)
);

XNOR2xp5_ASAP7_75t_L g713 ( 
.A(n_633),
.B(n_52),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_620),
.B(n_21),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_648),
.B(n_53),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_SL g716 ( 
.A1(n_696),
.A2(n_650),
.B1(n_657),
.B2(n_623),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_700),
.Y(n_717)
);

BUFx2_ASAP7_75t_SL g718 ( 
.A(n_700),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_689),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_713),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_700),
.Y(n_721)
);

CKINVDCx8_ASAP7_75t_R g722 ( 
.A(n_669),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_677),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_670),
.B(n_645),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_680),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_669),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_706),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_695),
.Y(n_729)
);

BUFx4f_ASAP7_75t_SL g730 ( 
.A(n_668),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_667),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_661),
.A2(n_651),
.B1(n_656),
.B2(n_638),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_658),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_682),
.B(n_623),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_666),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_662),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_681),
.B(n_22),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_686),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_663),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_694),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_665),
.B(n_22),
.Y(n_742)
);

BUFx10_ASAP7_75t_L g743 ( 
.A(n_693),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_664),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_658),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_666),
.Y(n_746)
);

BUFx2_ASAP7_75t_SL g747 ( 
.A(n_692),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_659),
.B(n_23),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_687),
.B(n_24),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_699),
.B(n_54),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_679),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_675),
.B(n_55),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_708),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_676),
.B(n_56),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_714),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_709),
.Y(n_757)
);

BUFx12f_ASAP7_75t_L g758 ( 
.A(n_715),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_674),
.B(n_707),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_702),
.Y(n_760)
);

INVx6_ASAP7_75t_L g761 ( 
.A(n_673),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_691),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_57),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_711),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_691),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_688),
.B(n_25),
.Y(n_767)
);

BUFx12f_ASAP7_75t_L g768 ( 
.A(n_704),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_703),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_701),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_703),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_690),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_671),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_672),
.B(n_26),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_678),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_712),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_737),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_762),
.A2(n_698),
.B1(n_685),
.B2(n_683),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_759),
.A2(n_660),
.B(n_133),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_755),
.B(n_58),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_740),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_736),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_725),
.A2(n_27),
.B(n_28),
.Y(n_783)
);

OAI211xp5_ASAP7_75t_L g784 ( 
.A1(n_725),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_756),
.B(n_751),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_741),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_776),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_736),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_759),
.A2(n_138),
.B(n_193),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_772),
.A2(n_135),
.B(n_192),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_735),
.A2(n_30),
.B(n_31),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_772),
.A2(n_763),
.B(n_732),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_749),
.A2(n_132),
.B(n_191),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_735),
.A2(n_30),
.B(n_31),
.Y(n_794)
);

OA21x2_ASAP7_75t_L g795 ( 
.A1(n_774),
.A2(n_60),
.B(n_62),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_736),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_755),
.B(n_63),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_751),
.B(n_64),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_736),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_723),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_765),
.B(n_731),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_726),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_66),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_747),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_749),
.A2(n_68),
.B(n_70),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_764),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_763),
.A2(n_76),
.B(n_78),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_775),
.A2(n_79),
.B(n_80),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_720),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_753),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_764),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_757),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_774),
.A2(n_84),
.B(n_85),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_757),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_771),
.Y(n_815)
);

CKINVDCx6p67_ASAP7_75t_R g816 ( 
.A(n_728),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_719),
.B(n_86),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_748),
.A2(n_88),
.B(n_89),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_748),
.A2(n_90),
.B(n_92),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_771),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_729),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_729),
.B(n_93),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_761),
.A2(n_730),
.B1(n_764),
.B2(n_770),
.Y(n_823)
);

OA21x2_ASAP7_75t_L g824 ( 
.A1(n_767),
.A2(n_94),
.B(n_96),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_767),
.A2(n_97),
.B(n_98),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_750),
.A2(n_99),
.B(n_100),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_752),
.A2(n_106),
.B(n_107),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_744),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_757),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_753),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_742),
.B(n_109),
.Y(n_831)
);

OAI21x1_ASAP7_75t_SL g832 ( 
.A1(n_766),
.A2(n_112),
.B(n_115),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_769),
.A2(n_771),
.B(n_766),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_785),
.B(n_773),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_777),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_777),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_792),
.A2(n_752),
.B(n_754),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_802),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_781),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_815),
.B(n_757),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_821),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_787),
.B(n_716),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_787),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_823),
.A2(n_768),
.B1(n_760),
.B2(n_730),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_786),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_SL g846 ( 
.A1(n_783),
.A2(n_761),
.B1(n_743),
.B2(n_773),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_800),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_779),
.A2(n_754),
.B(n_750),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_810),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_784),
.A2(n_761),
.B1(n_743),
.B2(n_769),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_830),
.B(n_738),
.Y(n_851)
);

BUFx2_ASAP7_75t_SL g852 ( 
.A(n_804),
.Y(n_852)
);

AOI21x1_ASAP7_75t_L g853 ( 
.A1(n_833),
.A2(n_739),
.B(n_758),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_791),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_812),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_801),
.B(n_746),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_812),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_815),
.B(n_771),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_814),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_821),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_779),
.A2(n_746),
.B(n_724),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_811),
.A2(n_716),
.B1(n_722),
.B2(n_733),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_809),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_814),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_829),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_778),
.A2(n_733),
.B(n_729),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_829),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_821),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_816),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_821),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_778),
.A2(n_718),
.B(n_717),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_791),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_828),
.Y(n_873)
);

OAI222xp33_ASAP7_75t_L g874 ( 
.A1(n_811),
.A2(n_724),
.B1(n_720),
.B2(n_745),
.C1(n_734),
.C2(n_727),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_824),
.B(n_727),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_793),
.A2(n_733),
.B1(n_729),
.B2(n_721),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_838),
.B(n_834),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_863),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_873),
.B(n_836),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_854),
.Y(n_880)
);

NOR2x1p5_ASAP7_75t_L g881 ( 
.A(n_869),
.B(n_803),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_863),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_839),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_846),
.A2(n_805),
.B1(n_826),
.B2(n_824),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_852),
.B(n_820),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_849),
.B(n_820),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_842),
.B(n_791),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_836),
.B(n_794),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_842),
.B(n_794),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_R g890 ( 
.A(n_869),
.B(n_782),
.Y(n_890)
);

AOI222xp33_ASAP7_75t_L g891 ( 
.A1(n_862),
.A2(n_831),
.B1(n_818),
.B2(n_819),
.C1(n_832),
.C2(n_798),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_844),
.B(n_798),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_853),
.B(n_782),
.Y(n_893)
);

CKINVDCx11_ASAP7_75t_R g894 ( 
.A(n_860),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_872),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_860),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_856),
.B(n_788),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_865),
.B(n_788),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_SL g899 ( 
.A(n_874),
.B(n_806),
.C(n_817),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_850),
.A2(n_827),
.B(n_818),
.C(n_819),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_857),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_870),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_865),
.B(n_796),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_845),
.B(n_794),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_R g905 ( 
.A(n_865),
.B(n_798),
.Y(n_905)
);

AO32x2_ASAP7_75t_L g906 ( 
.A1(n_855),
.A2(n_795),
.A3(n_825),
.B1(n_824),
.B2(n_734),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_880),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_880),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_895),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_895),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_887),
.B(n_858),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_894),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_877),
.B(n_879),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_888),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_857),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_904),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_883),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_886),
.B(n_835),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_898),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_896),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_906),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_898),
.B(n_867),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_896),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_885),
.B(n_903),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_903),
.B(n_858),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_896),
.B(n_867),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_896),
.B(n_867),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_906),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_925),
.B(n_897),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_908),
.Y(n_931)
);

OA21x2_ASAP7_75t_L g932 ( 
.A1(n_922),
.A2(n_929),
.B(n_907),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_908),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_924),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_925),
.B(n_906),
.Y(n_935)
);

INVxp67_ASAP7_75t_SL g936 ( 
.A(n_917),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_916),
.B(n_855),
.Y(n_937)
);

OAI211xp5_ASAP7_75t_L g938 ( 
.A1(n_922),
.A2(n_884),
.B(n_891),
.C(n_900),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_913),
.B(n_871),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_SL g940 ( 
.A1(n_912),
.A2(n_871),
.B1(n_878),
.B2(n_882),
.Y(n_940)
);

AO31x2_ASAP7_75t_L g941 ( 
.A1(n_929),
.A2(n_843),
.A3(n_845),
.B(n_847),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_912),
.A2(n_899),
.B(n_884),
.C(n_881),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_924),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_910),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_907),
.Y(n_945)
);

AOI222xp33_ASAP7_75t_L g946 ( 
.A1(n_938),
.A2(n_892),
.B1(n_912),
.B2(n_851),
.C1(n_914),
.C2(n_918),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_934),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_941),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_935),
.B(n_923),
.Y(n_949)
);

NOR2x1_ASAP7_75t_R g950 ( 
.A(n_942),
.B(n_912),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_934),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_945),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_932),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_936),
.B(n_911),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_935),
.B(n_923),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_934),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_934),
.B(n_923),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_957),
.B(n_943),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_957),
.B(n_943),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_952),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_953),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_950),
.B(n_912),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_954),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_947),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_949),
.B(n_930),
.Y(n_965)
);

NOR2x1_ASAP7_75t_R g966 ( 
.A(n_962),
.B(n_717),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_962),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_963),
.B(n_965),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_960),
.B(n_939),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_961),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_958),
.B(n_949),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_958),
.B(n_946),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_959),
.B(n_955),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_967),
.B(n_959),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_970),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_968),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_972),
.B(n_964),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_971),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_973),
.B(n_956),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_966),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_966),
.B(n_955),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_969),
.B(n_956),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_967),
.B(n_930),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_971),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_983),
.B(n_951),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_947),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_976),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_977),
.B(n_890),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_979),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_951),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_984),
.B(n_951),
.Y(n_992)
);

AND2x4_ASAP7_75t_SL g993 ( 
.A(n_979),
.B(n_951),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_985),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_989),
.A2(n_980),
.B1(n_981),
.B2(n_940),
.Y(n_995)
);

INVxp67_ASAP7_75t_SL g996 ( 
.A(n_990),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_986),
.A2(n_992),
.B(n_991),
.Y(n_997)
);

OAI211xp5_ASAP7_75t_SL g998 ( 
.A1(n_988),
.A2(n_975),
.B(n_982),
.C(n_943),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_993),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_987),
.A2(n_975),
.B(n_943),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_SL g1001 ( 
.A1(n_987),
.A2(n_945),
.B(n_951),
.C(n_937),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_985),
.B(n_933),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_994),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_999),
.B(n_924),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1002),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_933),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_997),
.B(n_995),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1000),
.B(n_933),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_1001),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_996),
.B(n_931),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_931),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_944),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1003),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_944),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1011),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_1006),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1005),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_SL g1019 ( 
.A(n_1009),
.B(n_893),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_1007),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1004),
.B(n_932),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_1014),
.B(n_924),
.Y(n_1022)
);

AOI211x1_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_909),
.B(n_914),
.C(n_920),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1021),
.Y(n_1024)
);

AOI221x1_ASAP7_75t_L g1025 ( 
.A1(n_1018),
.A2(n_1016),
.B1(n_1019),
.B2(n_1013),
.C(n_1012),
.Y(n_1025)
);

OAI221xp5_ASAP7_75t_SL g1026 ( 
.A1(n_1020),
.A2(n_921),
.B1(n_876),
.B2(n_948),
.C(n_937),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_1017),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_1020),
.B(n_924),
.Y(n_1028)
);

NOR2x1p5_ASAP7_75t_SL g1029 ( 
.A(n_1014),
.B(n_948),
.Y(n_1029)
);

AOI222xp33_ASAP7_75t_L g1030 ( 
.A1(n_1027),
.A2(n_921),
.B1(n_876),
.B2(n_910),
.C1(n_797),
.C2(n_780),
.Y(n_1030)
);

AOI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_1022),
.A2(n_899),
.B1(n_797),
.B2(n_780),
.C(n_822),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_932),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_R g1033 ( 
.A(n_1025),
.B(n_116),
.Y(n_1033)
);

XNOR2xp5_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_780),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_932),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_1026),
.A2(n_902),
.B(n_927),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_1032),
.B(n_1029),
.C(n_745),
.Y(n_1037)
);

AOI321xp33_ASAP7_75t_L g1038 ( 
.A1(n_1036),
.A2(n_822),
.A3(n_797),
.B1(n_866),
.B2(n_721),
.C(n_927),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_SL g1039 ( 
.A1(n_1034),
.A2(n_822),
.B(n_118),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1035),
.A2(n_928),
.B1(n_927),
.B2(n_915),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_1031),
.A2(n_827),
.B(n_789),
.C(n_790),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_SL g1042 ( 
.A1(n_1030),
.A2(n_875),
.B(n_928),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_1033),
.A2(n_825),
.B(n_790),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1033),
.A2(n_789),
.B(n_808),
.C(n_807),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1035),
.A2(n_813),
.B(n_825),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1032),
.B(n_795),
.C(n_905),
.Y(n_1046)
);

AOI222xp33_ASAP7_75t_L g1047 ( 
.A1(n_1037),
.A2(n_807),
.B1(n_911),
.B2(n_808),
.C1(n_733),
.C2(n_926),
.Y(n_1047)
);

NAND4xp25_ASAP7_75t_L g1048 ( 
.A(n_1038),
.B(n_841),
.C(n_868),
.D(n_926),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_941),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_1043),
.B(n_915),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_1042),
.A2(n_1044),
.B(n_1041),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1040),
.B(n_1045),
.C(n_1046),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1039),
.B(n_919),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_1037),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_1039),
.B(n_868),
.C(n_841),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_1037),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1055),
.B(n_1056),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1049),
.B(n_941),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1052),
.B(n_795),
.C(n_868),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

AND3x4_ASAP7_75t_L g1062 ( 
.A(n_1050),
.B(n_840),
.C(n_858),
.Y(n_1062)
);

AOI22x1_ASAP7_75t_L g1063 ( 
.A1(n_1047),
.A2(n_875),
.B1(n_841),
.B2(n_799),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1051),
.B(n_870),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_1048),
.B(n_941),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1055),
.B(n_941),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1056),
.A2(n_813),
.B1(n_799),
.B2(n_796),
.C(n_864),
.Y(n_1067)
);

OAI211xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1056),
.A2(n_117),
.B(n_123),
.C(n_127),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_1056),
.B(n_848),
.C(n_837),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1057),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1064),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1061),
.B(n_129),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_1058),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_SL g1074 ( 
.A(n_1062),
.B(n_864),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_1059),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1065),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1066),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_1063),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_1060),
.B1(n_1067),
.B2(n_1069),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1073),
.A2(n_1068),
.B1(n_919),
.B2(n_859),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_130),
.C(n_131),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1077),
.Y(n_1082)
);

AND3x2_ASAP7_75t_L g1083 ( 
.A(n_1072),
.B(n_139),
.C(n_141),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1076),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1078),
.Y(n_1085)
);

OAI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1075),
.A2(n_859),
.B1(n_847),
.B2(n_840),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1082),
.A2(n_1074),
.B1(n_840),
.B2(n_154),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1083),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1084),
.B(n_861),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1087),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_1085),
.B(n_1088),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_1079),
.B1(n_1080),
.B2(n_1081),
.Y(n_1092)
);

OAI222xp33_ASAP7_75t_L g1093 ( 
.A1(n_1092),
.A2(n_1086),
.B1(n_1089),
.B2(n_155),
.C1(n_156),
.C2(n_158),
.Y(n_1093)
);

XNOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_146),
.Y(n_1094)
);

AOI32xp33_ASAP7_75t_L g1095 ( 
.A1(n_1093),
.A2(n_1094),
.A3(n_861),
.B1(n_848),
.B2(n_162),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1094),
.Y(n_1096)
);

AOI222xp33_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_152),
.B1(n_159),
.B2(n_160),
.C1(n_163),
.C2(n_165),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1095),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_1098)
);

OA22x2_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_174),
.B(n_176),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1100),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.C(n_181),
.Y(n_1101)
);

AOI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_1099),
.B(n_184),
.C(n_185),
.Y(n_1102)
);


endmodule