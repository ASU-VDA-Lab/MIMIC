module fake_jpeg_10613_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_17),
.B1(n_19),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_43),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_22),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_60),
.B1(n_40),
.B2(n_19),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_19),
.Y(n_50)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_53),
.A3(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_63),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_30),
.B(n_27),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_20),
.C(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_17),
.B1(n_23),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_40),
.B1(n_32),
.B2(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_75),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_94),
.B1(n_23),
.B2(n_33),
.Y(n_101)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_76),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_53),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_116)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_82),
.B(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_18),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_88),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_39),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_78),
.B1(n_72),
.B2(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx9p33_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_23),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_36),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_32),
.B1(n_21),
.B2(n_28),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_18),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_0),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_114),
.B1(n_117),
.B2(n_72),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_103),
.A2(n_92),
.B(n_82),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_120),
.B1(n_86),
.B2(n_70),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_34),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_109),
.B(n_113),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_38),
.B1(n_39),
.B2(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_85),
.B1(n_68),
.B2(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_133),
.B1(n_142),
.B2(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_143),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_136),
.B1(n_100),
.B2(n_124),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_79),
.B1(n_71),
.B2(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_137),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_149),
.B(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_82),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_106),
.B(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_74),
.B1(n_82),
.B2(n_95),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_93),
.B1(n_65),
.B2(n_33),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_26),
.B1(n_25),
.B2(n_65),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_154),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_149)
);

AO21x2_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_26),
.B(n_25),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_25),
.B1(n_7),
.B2(n_8),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_103),
.C(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_7),
.C(n_12),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_168),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_165),
.B(n_166),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_100),
.B1(n_118),
.B2(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_155),
.B1(n_150),
.B2(n_137),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_104),
.B(n_117),
.C(n_100),
.D(n_114),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_164),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_149),
.B(n_126),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_102),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_184),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_118),
.C(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_179),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_185),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_118),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_6),
.C(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_111),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_152),
.CI(n_150),
.CON(n_192),
.SN(n_192)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_2),
.C(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_2),
.C(n_4),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_4),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_2),
.B1(n_14),
.B2(n_5),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_194),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_184),
.B1(n_175),
.B2(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_132),
.B1(n_136),
.B2(n_147),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_195),
.B(n_190),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_206),
.Y(n_221)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_178),
.B(n_151),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_217),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_166),
.B1(n_169),
.B2(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_161),
.B(n_165),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_158),
.B(n_177),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_188),
.B(n_192),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_6),
.B(n_10),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_189),
.A3(n_209),
.B1(n_192),
.B2(n_207),
.C1(n_205),
.C2(n_204),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_182),
.B1(n_169),
.B2(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_193),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_183),
.C(n_168),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_198),
.C(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_182),
.B1(n_165),
.B2(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_189),
.B1(n_206),
.B2(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_167),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_135),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_228),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_247),
.B1(n_225),
.B2(n_219),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_248),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_204),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_236),
.C(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_245),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_249),
.B1(n_237),
.B2(n_243),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_222),
.A2(n_196),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_251),
.C(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_226),
.C(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_226),
.C(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_227),
.C(n_218),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_242),
.C(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_256),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_234),
.B1(n_249),
.B2(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_217),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_255),
.A2(n_246),
.B(n_248),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_234),
.B1(n_224),
.B2(n_225),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_273),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.C(n_252),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_215),
.B(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_220),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_245),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_251),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_278),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_263),
.C(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_213),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_213),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_281),
.A2(n_270),
.B1(n_265),
.B2(n_273),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_284),
.B(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_268),
.B1(n_266),
.B2(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_287),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_223),
.B(n_231),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_6),
.A3(n_11),
.B1(n_12),
.B2(n_258),
.C1(n_277),
.C2(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.Y(n_296)
);


endmodule