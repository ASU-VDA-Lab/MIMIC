module fake_ariane_3361_n_107 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_107);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_107;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_5),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_5),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_7),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_26),
.B1(n_32),
.B2(n_28),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

OAI221xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_20),
.B1(n_25),
.B2(n_31),
.C(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_46),
.B1(n_40),
.B2(n_45),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_44),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_52),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_51),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_57),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AO32x1_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_46),
.A3(n_43),
.B1(n_38),
.B2(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI211xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_36),
.B(n_51),
.C(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_66),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_66),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_71),
.B(n_42),
.C(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_74),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_42),
.B1(n_41),
.B2(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_83),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_84),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_48),
.Y(n_95)
);

HAxp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_68),
.CON(n_96),
.SN(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_47),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_92),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_93),
.C(n_96),
.Y(n_101)
);

OR3x1_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_47),
.C(n_33),
.Y(n_102)
);

AOI222xp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_99),
.B1(n_29),
.B2(n_98),
.C1(n_102),
.C2(n_42),
.Y(n_103)
);

NAND4xp25_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_8),
.C(n_38),
.D(n_82),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_82),
.B1(n_64),
.B2(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_9),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_70),
.B1(n_12),
.B2(n_16),
.C(n_10),
.Y(n_107)
);


endmodule