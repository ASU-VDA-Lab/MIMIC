module fake_ibex_2003_n_1539 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_331, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1539);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1539;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1521;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_590;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1460;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1369;
wire n_1297;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g334 ( 
.A(n_190),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_108),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_5),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_158),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_315),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_58),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_332),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_279),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_43),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_196),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_144),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_22),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_115),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_23),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_3),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_74),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_160),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_75),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_134),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_23),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_199),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_241),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_283),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_324),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_12),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_325),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_233),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_90),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_179),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_244),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_310),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_67),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_282),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_0),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_27),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_114),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_58),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_85),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_205),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_189),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_14),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_148),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_150),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_316),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_226),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_224),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_157),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_293),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_198),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_35),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_289),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_103),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_70),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_168),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_84),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_299),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_237),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_15),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_30),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_53),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_94),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_106),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_111),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_25),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_292),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_222),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_209),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_60),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_323),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_246),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_130),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_240),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_284),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_73),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_81),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_156),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_254),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_277),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_197),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_11),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_65),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_29),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_37),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_122),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_220),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_92),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_268),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_255),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_213),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_70),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_275),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_164),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_307),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_153),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_82),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_88),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_173),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_300),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_230),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_296),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_178),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_140),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_232),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_193),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_172),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_118),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_102),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_80),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_231),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_326),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_281),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_313),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_312),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_305),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_314),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_175),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_311),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_171),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_273),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_124),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_21),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_136),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_16),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_303),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_12),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_218),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_110),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_319),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_72),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_306),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_0),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_261),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_72),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_192),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_260),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_290),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_276),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_184),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_288),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_186),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_256),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_98),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_30),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_60),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_128),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_322),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_216),
.Y(n_500)
);

BUFx2_ASAP7_75t_SL g501 ( 
.A(n_129),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_330),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_34),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_304),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_48),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_297),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_112),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_269),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_63),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_225),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_137),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_16),
.Y(n_512)
);

BUFx5_ASAP7_75t_L g513 ( 
.A(n_75),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_161),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_214),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_105),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_79),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_278),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_117),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_42),
.Y(n_520)
);

BUFx8_ASAP7_75t_SL g521 ( 
.A(n_272),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_3),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_113),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_104),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_274),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_20),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_321),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_138),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_257),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_280),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_191),
.Y(n_531)
);

CKINVDCx11_ASAP7_75t_R g532 ( 
.A(n_28),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_93),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_1),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_195),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_100),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_259),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_177),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_309),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_286),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_2),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_185),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_38),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_119),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_221),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_46),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_10),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_363),
.B(n_1),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_534),
.B(n_2),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_391),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_410),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_521),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_532),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_485),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_379),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_339),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_379),
.Y(n_559)
);

BUFx6f_ASAP7_75t_SL g560 ( 
.A(n_380),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_340),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_363),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_368),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_374),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_389),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_425),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_404),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_447),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_353),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_404),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_432),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_341),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_486),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_445),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_354),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_451),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_357),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_480),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_507),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_357),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_436),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_357),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_416),
.B(n_4),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_357),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_L g586 ( 
.A(n_358),
.B(n_4),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_336),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_536),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_357),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_428),
.B(n_5),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_402),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_364),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_407),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_513),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_440),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_359),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_513),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_440),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_513),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_372),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_362),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_349),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_385),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_381),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_349),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_409),
.B(n_6),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_411),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_415),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_419),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_390),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_401),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_427),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_435),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_433),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_443),
.B(n_6),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_434),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_547),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_429),
.B(n_7),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_578),
.B(n_384),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_571),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_581),
.B(n_384),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_600),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_583),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_590),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_570),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_595),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_559),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_557),
.B(n_474),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_551),
.B(n_334),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_559),
.B(n_401),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_598),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_601),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_603),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_609),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_584),
.B(n_384),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_568),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_553),
.B(n_476),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_493),
.Y(n_648)
);

INVxp33_ASAP7_75t_SL g649 ( 
.A(n_594),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_618),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_611),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_597),
.B(n_617),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_612),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_619),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_613),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_548),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_622),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_SL g660 ( 
.A(n_597),
.B(n_382),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_576),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_604),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_596),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_586),
.Y(n_665)
);

OA21x2_ASAP7_75t_L g666 ( 
.A1(n_591),
.A2(n_346),
.B(n_338),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_599),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_552),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_607),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_610),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_564),
.B(n_496),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_617),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_567),
.B(n_542),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_569),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_593),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_621),
.B(n_342),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_602),
.B(n_384),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_606),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_560),
.B(n_365),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_614),
.A2(n_371),
.B(n_367),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_560),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_616),
.B(n_350),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_620),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_605),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_605),
.A2(n_483),
.B(n_414),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_608),
.B(n_508),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_615),
.B(n_380),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_589),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_561),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_565),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_566),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_572),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_577),
.B(n_539),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_580),
.A2(n_386),
.B(n_376),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_588),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_555),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_575),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_575),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_579),
.Y(n_704)
);

OA21x2_ASAP7_75t_L g705 ( 
.A1(n_579),
.A2(n_388),
.B(n_387),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_573),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_574),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_600),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_557),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_559),
.B(n_456),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_571),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_557),
.B(n_517),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_559),
.B(n_456),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_600),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_600),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_578),
.A2(n_393),
.B(n_392),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_600),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_570),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_570),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_557),
.B(n_523),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_571),
.Y(n_724)
);

CKINVDCx16_ASAP7_75t_R g725 ( 
.A(n_550),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_557),
.B(n_523),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_600),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_571),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_571),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_557),
.B(n_396),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_557),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_564),
.B(n_444),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_557),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_559),
.B(n_382),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_600),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_600),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_571),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_600),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_557),
.B(n_408),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_600),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_570),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_602),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_578),
.B(n_384),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_571),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_571),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_571),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_602),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_571),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_557),
.B(n_413),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_559),
.B(n_472),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_571),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_571),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_552),
.A2(n_478),
.B1(n_484),
.B2(n_482),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_570),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_709),
.B(n_472),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_716),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_672),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_653),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_635),
.B(n_497),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_634),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_679),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_629),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_624),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_692),
.B(n_501),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_725),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_635),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_645),
.B(n_335),
.Y(n_772)
);

AO21x2_ASAP7_75t_L g773 ( 
.A1(n_623),
.A2(n_418),
.B(n_417),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_711),
.Y(n_774)
);

OR2x2_ASAP7_75t_SL g775 ( 
.A(n_668),
.B(n_382),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_719),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_661),
.B(n_337),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_651),
.A2(n_382),
.B1(n_522),
.B2(n_431),
.Y(n_778)
);

XNOR2x2_ASAP7_75t_L g779 ( 
.A(n_650),
.B(n_686),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_661),
.B(n_343),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_645),
.B(n_651),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_628),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_709),
.B(n_731),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_722),
.B(n_344),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_668),
.B(n_503),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_679),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_731),
.B(n_345),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_679),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_654),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_654),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_656),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_628),
.Y(n_792)
);

INVxp33_ASAP7_75t_L g793 ( 
.A(n_638),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_723),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_669),
.B(n_655),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_636),
.B(n_520),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_724),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_722),
.B(n_347),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_744),
.B(n_522),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_728),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_655),
.B(n_505),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_729),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_636),
.B(n_509),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_628),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_742),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_751),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_683),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_679),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_734),
.B(n_659),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_721),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_683),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_738),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_721),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_657),
.B(n_512),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_746),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_721),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_683),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_726),
.B(n_348),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_644),
.B(n_351),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_683),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_634),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_747),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_721),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_736),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_726),
.B(n_352),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_710),
.B(n_526),
.Y(n_831)
);

NOR2x1_ASAP7_75t_L g832 ( 
.A(n_681),
.B(n_421),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_649),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_742),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_730),
.B(n_355),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_662),
.B(n_400),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_356),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_750),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_736),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_752),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_712),
.B(n_541),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_713),
.B(n_543),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_692),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_736),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_678),
.B(n_658),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_755),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_736),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_647),
.B(n_463),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_704),
.A2(n_546),
.B1(n_438),
.B2(n_439),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_756),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_754),
.B(n_522),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_649),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_703),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_712),
.B(n_522),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_737),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_740),
.B(n_360),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_757),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_737),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_656),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_758),
.B(n_674),
.Y(n_861)
);

INVx8_ASAP7_75t_L g862 ( 
.A(n_678),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_637),
.A2(n_448),
.B1(n_457),
.B2(n_453),
.Y(n_863)
);

BUFx8_ASAP7_75t_SL g864 ( 
.A(n_701),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_633),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_633),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_652),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_685),
.B(n_460),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_737),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_688),
.B(n_464),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_740),
.B(n_753),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_671),
.B(n_465),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_646),
.B(n_494),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_637),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_646),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_753),
.B(n_361),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_671),
.B(n_366),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_687),
.B(n_7),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_676),
.B(n_682),
.Y(n_879)
);

AND2x2_ASAP7_75t_SL g880 ( 
.A(n_689),
.B(n_466),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_718),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_720),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_720),
.B(n_369),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_634),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_637),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_634),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_727),
.Y(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_637),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_703),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_664),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_665),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_680),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_648),
.B(n_370),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_676),
.B(n_373),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_664),
.B(n_467),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_666),
.A2(n_479),
.B1(n_488),
.B2(n_481),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_667),
.B(n_489),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_682),
.B(n_375),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_666),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_667),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_675),
.B(n_544),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_687),
.B(n_377),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_670),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_663),
.B(n_378),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_680),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_632),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_627),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_697),
.B(n_383),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_690),
.B(n_490),
.Y(n_909)
);

AO22x2_ASAP7_75t_L g910 ( 
.A1(n_704),
.A2(n_702),
.B1(n_707),
.B2(n_706),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_673),
.B(n_394),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_708),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_714),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_660),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_698),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_732),
.B(n_395),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_698),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_707),
.B(n_8),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_691),
.B(n_491),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_735),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_715),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_693),
.B(n_492),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_735),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_660),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_697),
.B(n_540),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_643),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_703),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_630),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_677),
.B(n_397),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_684),
.B(n_8),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_696),
.B(n_495),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_643),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_677),
.B(n_398),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_741),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_743),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_623),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_639),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_694),
.B(n_500),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_703),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_705),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_640),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_625),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_631),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_625),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_695),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_641),
.B(n_399),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_642),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_745),
.Y(n_950)
);

INVx4_ASAP7_75t_SL g951 ( 
.A(n_699),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_705),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_745),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_702),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_700),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_626),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_L g957 ( 
.A(n_786),
.B(n_384),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_888),
.B(n_538),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_951),
.B(n_502),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_871),
.A2(n_510),
.B1(n_511),
.B2(n_506),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_783),
.B(n_403),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_808),
.B(n_514),
.Y(n_962)
);

AO22x2_ASAP7_75t_L g963 ( 
.A1(n_942),
.A2(n_528),
.B1(n_529),
.B2(n_515),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_855),
.Y(n_964)
);

AND2x2_ASAP7_75t_SL g965 ( 
.A(n_844),
.B(n_504),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_952),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_855),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_852),
.Y(n_968)
);

OAI221xp5_ASAP7_75t_L g969 ( 
.A1(n_762),
.A2(n_412),
.B1(n_420),
.B2(n_406),
.C(n_405),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_825),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_951),
.B(n_9),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_888),
.B(n_537),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_811),
.B(n_422),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_928),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_761),
.B(n_423),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_928),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_945),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_945),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_768),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_902),
.B(n_424),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_774),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_949),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_776),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_949),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_771),
.Y(n_985)
);

AO22x2_ASAP7_75t_L g986 ( 
.A1(n_915),
.A2(n_917),
.B1(n_892),
.B2(n_878),
.Y(n_986)
);

AO22x2_ASAP7_75t_L g987 ( 
.A1(n_892),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_925),
.B(n_426),
.Y(n_988)
);

AO22x2_ASAP7_75t_L g989 ( 
.A1(n_796),
.A2(n_18),
.B1(n_13),
.B2(n_17),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_794),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_797),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_890),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_801),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_781),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_816),
.B(n_17),
.Y(n_995)
);

CKINVDCx14_ASAP7_75t_R g996 ( 
.A(n_834),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_803),
.Y(n_997)
);

AO22x2_ASAP7_75t_L g998 ( 
.A1(n_796),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_804),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_853),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_769),
.B(n_19),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_814),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_781),
.B(n_430),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_817),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_826),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_827),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_793),
.A2(n_441),
.B(n_437),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_802),
.B(n_785),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_805),
.A2(n_446),
.B1(n_449),
.B2(n_442),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_947),
.B(n_900),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_769),
.B(n_21),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_795),
.B(n_450),
.Y(n_1012)
);

AO22x2_ASAP7_75t_L g1013 ( 
.A1(n_918),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_805),
.B(n_842),
.Y(n_1014)
);

OAI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_850),
.A2(n_487),
.B1(n_533),
.B2(n_531),
.C(n_530),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_879),
.B(n_452),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_833),
.Y(n_1017)
);

BUFx8_ASAP7_75t_L g1018 ( 
.A(n_955),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_831),
.B(n_24),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_836),
.B(n_454),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_763),
.B(n_26),
.Y(n_1021)
);

AO22x2_ASAP7_75t_L g1022 ( 
.A1(n_775),
.A2(n_842),
.B1(n_927),
.B2(n_930),
.Y(n_1022)
);

OAI221xp5_ASAP7_75t_L g1023 ( 
.A1(n_868),
.A2(n_535),
.B1(n_527),
.B2(n_525),
.C(n_524),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_839),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_843),
.B(n_455),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_880),
.A2(n_461),
.B1(n_462),
.B2(n_458),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_841),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_900),
.B(n_504),
.Y(n_1028)
);

AND2x6_ASAP7_75t_SL g1029 ( 
.A(n_909),
.B(n_29),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_847),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_824),
.B(n_866),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_851),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_907),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_858),
.A2(n_469),
.B1(n_470),
.B2(n_468),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_838),
.B(n_471),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_789),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_867),
.Y(n_1037)
);

AO22x2_ASAP7_75t_L g1038 ( 
.A1(n_872),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1038)
);

OR2x6_ASAP7_75t_SL g1039 ( 
.A(n_770),
.B(n_519),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_790),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_790),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_791),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_791),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_864),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_857),
.B(n_473),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_518),
.B1(n_475),
.B2(n_477),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_765),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_866),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_875),
.B(n_504),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_860),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_767),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_854),
.Y(n_1052)
);

AO22x2_ASAP7_75t_L g1053 ( 
.A1(n_895),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_1053)
);

AO22x2_ASAP7_75t_L g1054 ( 
.A1(n_895),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_956),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_903),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_940),
.A2(n_499),
.B1(n_516),
.B2(n_498),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_881),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_901),
.B(n_39),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_882),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_865),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_865),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_906),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_887),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_939),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_889),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_911),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_943),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_870),
.A2(n_830),
.B1(n_837),
.B2(n_849),
.C(n_922),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_941),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_912),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_898),
.B(n_39),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_861),
.Y(n_1074)
);

AO22x2_ASAP7_75t_L g1075 ( 
.A1(n_897),
.A2(n_779),
.B1(n_910),
.B2(n_920),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_923),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_954),
.B(n_40),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_832),
.B(n_40),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_954),
.B(n_41),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_875),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_807),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_835),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_835),
.Y(n_1083)
);

AO22x2_ASAP7_75t_L g1084 ( 
.A1(n_897),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_862),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_870),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_954),
.B(n_45),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_910),
.Y(n_1088)
);

AO22x2_ASAP7_75t_L g1089 ( 
.A1(n_784),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_913),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_921),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_905),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_931),
.Y(n_1093)
);

AO22x2_ASAP7_75t_L g1094 ( 
.A1(n_798),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_862),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_799),
.Y(n_1096)
);

AO22x2_ASAP7_75t_L g1097 ( 
.A1(n_820),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_934),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_936),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_877),
.B(n_57),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_893),
.B(n_57),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_916),
.B(n_59),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_759),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_821),
.B(n_61),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_937),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_899),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_926),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_777),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1008),
.B(n_772),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_965),
.B(n_885),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_985),
.B(n_885),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_970),
.B(n_873),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_962),
.B(n_885),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1010),
.B(n_788),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1010),
.B(n_788),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_971),
.B(n_810),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_SL g1117 ( 
.A(n_971),
.B(n_810),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_SL g1118 ( 
.A(n_1096),
.B(n_905),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_SL g1119 ( 
.A(n_1068),
.B(n_1064),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1018),
.B(n_766),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_SL g1121 ( 
.A(n_1001),
.B(n_1011),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_995),
.B(n_905),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_SL g1123 ( 
.A(n_1052),
.B(n_760),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1071),
.B(n_766),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1085),
.B(n_819),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1095),
.B(n_819),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1014),
.B(n_787),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1067),
.B(n_883),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1046),
.B(n_760),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1058),
.B(n_863),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1009),
.B(n_1034),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1019),
.B(n_809),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1000),
.B(n_813),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1026),
.B(n_822),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_979),
.B(n_919),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_992),
.B(n_780),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_981),
.B(n_932),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_983),
.B(n_932),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1025),
.B(n_764),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1036),
.B(n_764),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1040),
.B(n_764),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1087),
.B(n_823),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1087),
.B(n_823),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_SL g1144 ( 
.A(n_1060),
.B(n_899),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1088),
.B(n_899),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1048),
.B(n_823),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_990),
.B(n_932),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1108),
.B(n_948),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1031),
.B(n_896),
.Y(n_1149)
);

NAND2xp33_ASAP7_75t_SL g1150 ( 
.A(n_1021),
.B(n_894),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_982),
.B(n_914),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_908),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_984),
.B(n_924),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1007),
.B(n_929),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_993),
.B(n_846),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_988),
.B(n_935),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_SL g1157 ( 
.A(n_974),
.B(n_950),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_959),
.B(n_950),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_959),
.B(n_950),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_SL g1160 ( 
.A(n_976),
.B(n_933),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_994),
.B(n_904),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_980),
.B(n_1079),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1003),
.B(n_778),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_989),
.B(n_932),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_977),
.B(n_938),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_978),
.B(n_944),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_997),
.B(n_846),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_989),
.B(n_846),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1074),
.B(n_946),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1012),
.B(n_953),
.Y(n_1170)
);

NAND2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1102),
.B(n_829),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1078),
.B(n_829),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1104),
.B(n_829),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1078),
.B(n_845),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1041),
.B(n_1042),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1043),
.B(n_845),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1047),
.B(n_845),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1055),
.B(n_856),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_999),
.B(n_846),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1051),
.B(n_856),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1073),
.B(n_884),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1080),
.B(n_1077),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1002),
.B(n_886),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_SL g1184 ( 
.A(n_1004),
.B(n_773),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1005),
.B(n_782),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1006),
.B(n_1017),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1024),
.B(n_792),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1027),
.B(n_800),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1020),
.B(n_806),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1035),
.B(n_812),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1045),
.B(n_815),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1100),
.B(n_818),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1050),
.B(n_828),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1037),
.B(n_840),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1056),
.B(n_848),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1057),
.B(n_869),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1065),
.B(n_859),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_975),
.B(n_66),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_961),
.B(n_66),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_960),
.B(n_67),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_968),
.B(n_68),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_SL g1203 ( 
.A(n_1101),
.B(n_68),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1070),
.B(n_69),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_973),
.B(n_71),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1072),
.B(n_71),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1066),
.B(n_74),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1099),
.B(n_76),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1105),
.B(n_76),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1049),
.B(n_77),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1090),
.B(n_77),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1091),
.B(n_78),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1093),
.B(n_78),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1015),
.B(n_79),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1098),
.B(n_83),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1069),
.B(n_1028),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1059),
.B(n_86),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1016),
.B(n_87),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1103),
.B(n_89),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1061),
.B(n_91),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_964),
.B(n_967),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_963),
.B(n_95),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1063),
.B(n_96),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_998),
.B(n_97),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1033),
.B(n_99),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1081),
.B(n_101),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1062),
.B(n_1076),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1228)
);

BUFx8_ASAP7_75t_L g1229 ( 
.A(n_1224),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1222),
.A2(n_1106),
.A3(n_1075),
.B(n_986),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1202),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1202),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1120),
.B(n_1044),
.Y(n_1233)
);

NAND2x1_ASAP7_75t_L g1234 ( 
.A(n_1217),
.B(n_1220),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1119),
.B(n_1217),
.Y(n_1235)
);

NOR4xp25_ASAP7_75t_L g1236 ( 
.A(n_1164),
.B(n_1086),
.C(n_1092),
.D(n_998),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1204),
.A2(n_1075),
.A3(n_986),
.B(n_963),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1189),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1184),
.A2(n_957),
.B(n_1022),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_SL g1240 ( 
.A(n_1110),
.B(n_1039),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1177),
.A2(n_972),
.B(n_958),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1178),
.A2(n_987),
.B(n_966),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1181),
.A2(n_1185),
.B(n_1190),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1191),
.A2(n_1022),
.B(n_987),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1121),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1129),
.A2(n_1176),
.B(n_1180),
.Y(n_1246)
);

AO32x2_ASAP7_75t_L g1247 ( 
.A1(n_1145),
.A2(n_966),
.A3(n_1013),
.B1(n_1107),
.B2(n_1089),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1112),
.B(n_1023),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1127),
.B(n_1053),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1220),
.A2(n_1013),
.B1(n_1084),
.B2(n_1053),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1155),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1152),
.B(n_1113),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1192),
.A2(n_1094),
.B(n_1089),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1109),
.B(n_1054),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1131),
.B(n_996),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1133),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1142),
.A2(n_1084),
.B(n_1054),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1214),
.A2(n_1029),
.B1(n_969),
.B2(n_1038),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1152),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1186),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1163),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1182),
.A2(n_1107),
.B(n_1097),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1219),
.A2(n_1097),
.B(n_1094),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1128),
.B(n_1038),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1215),
.A2(n_107),
.B(n_109),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1227),
.B(n_116),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1156),
.A2(n_120),
.B(n_121),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1207),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1155),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1161),
.B(n_333),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1167),
.A2(n_123),
.A3(n_125),
.B(n_126),
.Y(n_1271)
);

AO22x2_ASAP7_75t_L g1272 ( 
.A1(n_1168),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1175),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1179),
.A2(n_133),
.A3(n_135),
.B(n_139),
.Y(n_1274)
);

OAI21xp33_ASAP7_75t_L g1275 ( 
.A1(n_1201),
.A2(n_141),
.B(n_142),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1160),
.A2(n_1195),
.B(n_1154),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1216),
.A2(n_143),
.B(n_145),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1135),
.A2(n_146),
.A3(n_147),
.B(n_149),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1225),
.A2(n_1223),
.B(n_1226),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1162),
.B(n_151),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1143),
.A2(n_1174),
.B1(n_1172),
.B2(n_1138),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1196),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1136),
.B(n_152),
.Y(n_1283)
);

AOI211x1_ASAP7_75t_L g1284 ( 
.A1(n_1199),
.A2(n_154),
.B(n_155),
.C(n_159),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1137),
.A2(n_162),
.B(n_163),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1147),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1197),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1169),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1123),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1132),
.B(n_165),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1144),
.A2(n_166),
.A3(n_167),
.B(n_169),
.Y(n_1291)
);

AOI221x1_ASAP7_75t_L g1292 ( 
.A1(n_1122),
.A2(n_170),
.B1(n_174),
.B2(n_181),
.C(n_183),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1158),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1203),
.A2(n_187),
.B1(n_188),
.B2(n_194),
.Y(n_1294)
);

AOI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1149),
.A2(n_331),
.B(n_201),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_1200),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1210),
.A2(n_204),
.B(n_206),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1150),
.A2(n_207),
.B(n_208),
.C(n_210),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1170),
.A2(n_211),
.B(n_212),
.Y(n_1299)
);

BUFx2_ASAP7_75t_R g1300 ( 
.A(n_1124),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1205),
.A2(n_215),
.B(n_217),
.C(n_219),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1193),
.A2(n_223),
.B(n_227),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1116),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1159),
.B(n_228),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1117),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1198),
.A2(n_229),
.B(n_234),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1234),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1239),
.A2(n_1218),
.B(n_1206),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1244),
.A2(n_1118),
.A3(n_1171),
.B(n_1173),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1282),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1229),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1250),
.A2(n_1212),
.B1(n_1213),
.B2(n_1211),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1287),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1260),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1242),
.A2(n_1208),
.B(n_1209),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1246),
.A2(n_1194),
.B(n_1188),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1247),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1279),
.A2(n_1187),
.B(n_1153),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1236),
.A2(n_1139),
.B(n_1134),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1273),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1269),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1231),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1278),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1247),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1251),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1266),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1266),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1264),
.A2(n_1228),
.B1(n_1157),
.B2(n_1165),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1235),
.A2(n_1114),
.B1(n_1115),
.B2(n_1166),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1247),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1253),
.A2(n_1151),
.B(n_1183),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1278),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1262),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1259),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1245),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1303),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1268),
.A2(n_1111),
.B(n_1141),
.C(n_1140),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1277),
.A2(n_1146),
.B(n_1221),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1263),
.A2(n_1276),
.B(n_1261),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1252),
.B(n_1125),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1238),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1292),
.A2(n_1126),
.B(n_236),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1249),
.B(n_235),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_L g1344 ( 
.A(n_1255),
.B(n_238),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1272),
.B(n_239),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1291),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1243),
.A2(n_327),
.A3(n_243),
.B(n_245),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1258),
.B(n_1248),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1291),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1265),
.A2(n_242),
.B(n_247),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1272),
.B(n_248),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1313),
.B(n_1254),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1345),
.A2(n_1252),
.B1(n_1240),
.B2(n_1232),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1322),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1313),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1320),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1326),
.B(n_1230),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1320),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1326),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1333),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1333),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1341),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1341),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1314),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1317),
.B(n_1230),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1345),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1351),
.B(n_1257),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1317),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1346),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1346),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1310),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1334),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1342),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1307),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1311),
.A2(n_1256),
.B1(n_1305),
.B2(n_1289),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1324),
.B(n_1237),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1311),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1349),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1349),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1324),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1348),
.B(n_1288),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1377),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1376),
.B(n_1330),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1354),
.B(n_1330),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_R g1385 ( 
.A(n_1367),
.B(n_1351),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1364),
.B(n_1307),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_R g1387 ( 
.A(n_1359),
.B(n_1321),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1359),
.B(n_1321),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_R g1389 ( 
.A(n_1359),
.B(n_1336),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1353),
.B(n_1327),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1364),
.B(n_1327),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1374),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1375),
.Y(n_1393)
);

XNOR2xp5_ASAP7_75t_L g1394 ( 
.A(n_1367),
.B(n_1233),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1372),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1355),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1367),
.B(n_1309),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_R g1399 ( 
.A(n_1376),
.B(n_1283),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1362),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_R g1401 ( 
.A(n_1357),
.B(n_1283),
.Y(n_1401)
);

XNOR2xp5_ASAP7_75t_L g1402 ( 
.A(n_1381),
.B(n_1344),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1362),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1363),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1352),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1395),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1383),
.B(n_1368),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1396),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1383),
.B(n_1365),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1405),
.A2(n_1312),
.B1(n_1319),
.B2(n_1340),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1400),
.Y(n_1411)
);

AOI222xp33_ASAP7_75t_L g1412 ( 
.A1(n_1390),
.A2(n_1380),
.B1(n_1368),
.B2(n_1335),
.C1(n_1357),
.C2(n_1360),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1384),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1403),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1402),
.B(n_1380),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1404),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1398),
.B(n_1369),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1392),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1392),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1393),
.A2(n_1340),
.B1(n_1296),
.B2(n_1325),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1398),
.B(n_1369),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1391),
.B(n_1371),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1382),
.B(n_1340),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1420),
.A2(n_1385),
.B1(n_1399),
.B2(n_1401),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1406),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1409),
.B(n_1386),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1413),
.B(n_1360),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1414),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1419),
.A2(n_1332),
.B(n_1323),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1415),
.A2(n_1397),
.A3(n_1361),
.B(n_1370),
.Y(n_1431)
);

OAI31xp33_ASAP7_75t_L g1432 ( 
.A1(n_1420),
.A2(n_1394),
.A3(n_1296),
.B(n_1387),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1418),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1418),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1425),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1434),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1428),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1429),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1433),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1427),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1426),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1427),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1431),
.B(n_1417),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1430),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1430),
.Y(n_1445)
);

NAND2xp33_ASAP7_75t_SL g1446 ( 
.A(n_1439),
.B(n_1388),
.Y(n_1446)
);

AND2x4_ASAP7_75t_SL g1447 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1447)
);

AND2x4_ASAP7_75t_SL g1448 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1436),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1441),
.A2(n_1424),
.B1(n_1410),
.B2(n_1432),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1449),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1446),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1450),
.A2(n_1424),
.B1(n_1415),
.B2(n_1443),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1451),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1454),
.B(n_1452),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1454),
.B(n_1453),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1454),
.B(n_1442),
.Y(n_1457)
);

XNOR2x1_ASAP7_75t_L g1458 ( 
.A(n_1455),
.B(n_1438),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1457),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1456),
.B(n_1440),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1457),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1457),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1455),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1463),
.B(n_1461),
.C(n_1459),
.Y(n_1464)
);

NAND4xp25_ASAP7_75t_SL g1465 ( 
.A(n_1462),
.B(n_1412),
.C(n_1410),
.D(n_1435),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1458),
.A2(n_1448),
.B1(n_1447),
.B2(n_1442),
.Y(n_1466)
);

O2A1O1Ixp5_ASAP7_75t_SL g1467 ( 
.A1(n_1460),
.A2(n_1435),
.B(n_1270),
.C(n_1295),
.Y(n_1467)
);

NOR3x1_ASAP7_75t_L g1468 ( 
.A(n_1460),
.B(n_1343),
.C(n_1389),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_L g1469 ( 
.A(n_1463),
.B(n_1444),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_SL g1470 ( 
.A(n_1463),
.B(n_1294),
.C(n_1298),
.Y(n_1470)
);

NOR4xp25_ASAP7_75t_L g1471 ( 
.A(n_1463),
.B(n_1445),
.C(n_1444),
.D(n_1301),
.Y(n_1471)
);

NAND4xp25_ASAP7_75t_SL g1472 ( 
.A(n_1463),
.B(n_1445),
.C(n_1437),
.D(n_1328),
.Y(n_1472)
);

AOI211xp5_ASAP7_75t_L g1473 ( 
.A1(n_1463),
.A2(n_1329),
.B(n_1337),
.C(n_1281),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1464),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_SL g1475 ( 
.A(n_1471),
.B(n_1267),
.C(n_1299),
.Y(n_1475)
);

OAI211xp5_ASAP7_75t_L g1476 ( 
.A1(n_1469),
.A2(n_1284),
.B(n_1297),
.C(n_1275),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1466),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1465),
.B(n_1300),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1467),
.B(n_1290),
.C(n_1280),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1472),
.A2(n_1421),
.B1(n_1417),
.B2(n_1339),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1468),
.Y(n_1481)
);

AND3x2_ASAP7_75t_L g1482 ( 
.A(n_1473),
.B(n_1304),
.C(n_1293),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1470),
.A2(n_1421),
.B1(n_1339),
.B2(n_1422),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1464),
.A2(n_1407),
.B1(n_1416),
.B2(n_1411),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_1477),
.Y(n_1485)
);

XNOR2x1_ASAP7_75t_L g1486 ( 
.A(n_1474),
.B(n_1304),
.Y(n_1486)
);

XOR2xp5_ASAP7_75t_L g1487 ( 
.A(n_1481),
.B(n_1479),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1482),
.B(n_1431),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1484),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1483),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1478),
.B(n_1411),
.Y(n_1491)
);

NAND3x1_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1285),
.C(n_1302),
.Y(n_1492)
);

OR3x2_ASAP7_75t_L g1493 ( 
.A(n_1475),
.B(n_1347),
.C(n_1291),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1476),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1481),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1481),
.B(n_1416),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1485),
.B(n_1361),
.Y(n_1497)
);

NAND2x1_ASAP7_75t_SL g1498 ( 
.A(n_1495),
.B(n_1342),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1494),
.B(n_249),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_SL g1500 ( 
.A(n_1487),
.B(n_1306),
.C(n_1347),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1489),
.B(n_1286),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_R g1502 ( 
.A(n_1490),
.B(n_250),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_R g1503 ( 
.A(n_1496),
.B(n_1491),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_R g1504 ( 
.A(n_1496),
.B(n_251),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_SL g1505 ( 
.A(n_1486),
.B(n_1373),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1488),
.B(n_1373),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1492),
.B(n_1339),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_SL g1508 ( 
.A(n_1493),
.B(n_252),
.C(n_253),
.Y(n_1508)
);

XNOR2xp5_ASAP7_75t_L g1509 ( 
.A(n_1486),
.B(n_1315),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_SL g1510 ( 
.A(n_1494),
.B(n_1373),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1497),
.B(n_1315),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1508),
.B(n_1347),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1501),
.B(n_1347),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1500),
.A2(n_1331),
.B1(n_1373),
.B2(n_1358),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1499),
.B(n_1241),
.Y(n_1515)
);

OAI22x1_ASAP7_75t_L g1516 ( 
.A1(n_1502),
.A2(n_1342),
.B1(n_1315),
.B2(n_1347),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1505),
.A2(n_1331),
.B1(n_1358),
.B2(n_1356),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1503),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1498),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1507),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_SL g1521 ( 
.A(n_1518),
.B(n_1504),
.C(n_1510),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1519),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_SL g1523 ( 
.A1(n_1512),
.A2(n_1509),
.B(n_1506),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1515),
.Y(n_1524)
);

AO221x2_ASAP7_75t_L g1525 ( 
.A1(n_1513),
.A2(n_1516),
.B1(n_1514),
.B2(n_1511),
.C(n_1517),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1518),
.B(n_1309),
.Y(n_1526)
);

OAI321xp33_ASAP7_75t_L g1527 ( 
.A1(n_1520),
.A2(n_1356),
.A3(n_1378),
.B1(n_1379),
.B2(n_1271),
.C(n_1274),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1522),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1521),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1526),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1524),
.B(n_1350),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1523),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1528),
.A2(n_1525),
.B1(n_1527),
.B2(n_1308),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1529),
.A2(n_1350),
.B1(n_1338),
.B2(n_1308),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1533),
.A2(n_1532),
.B1(n_1530),
.B2(n_1531),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1534),
.B1(n_1338),
.B2(n_1378),
.C1(n_1318),
.C2(n_1316),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1536),
.Y(n_1537)
);

AOI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.C(n_266),
.Y(n_1538)
);

AOI211xp5_ASAP7_75t_L g1539 ( 
.A1(n_1538),
.A2(n_267),
.B(n_270),
.C(n_271),
.Y(n_1539)
);


endmodule