module real_jpeg_10898_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_44),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_1),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_1),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_31),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_35),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_3),
.B(n_32),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_109),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_2),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_96),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_96),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_96),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_7),
.A2(n_31),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_9),
.A2(n_23),
.B1(n_60),
.B2(n_61),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_9),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_10),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_125),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_125),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_144),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_144),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_144),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_84),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_84),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_84),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_14),
.A2(n_34),
.B1(n_60),
.B2(n_61),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_15),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_16),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_89),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_329),
.B(n_332),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_71),
.B(n_328),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_21),
.B(n_36),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_21),
.B(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_21),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_22),
.A2(n_26),
.B1(n_35),
.B2(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_24),
.A2(n_28),
.B(n_109),
.C(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_26),
.A2(n_35),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_331)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_30),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_27),
.A2(n_30),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_27),
.A2(n_30),
.B1(n_207),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_27),
.A2(n_30),
.B1(n_232),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_27),
.A2(n_30),
.B1(n_250),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_27),
.A2(n_30),
.B1(n_51),
.B2(n_276),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_64),
.C(n_66),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_37),
.A2(n_38),
.B1(n_323),
.B2(n_325),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_49),
.C(n_55),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_39),
.A2(n_40),
.B1(n_55),
.B2(n_303),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_41),
.A2(n_43),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_41),
.A2(n_43),
.B1(n_135),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_41),
.A2(n_43),
.B1(n_152),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_41),
.A2(n_43),
.B1(n_192),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_41),
.A2(n_43),
.B1(n_203),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_41),
.A2(n_43),
.B1(n_229),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_42),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_43),
.B(n_109),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_44),
.B(n_46),
.Y(n_139)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_45),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_49),
.A2(n_50),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_55),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_55),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_63),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_59),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_59),
.B1(n_95),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_59),
.B1(n_122),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_56),
.A2(n_59),
.B1(n_131),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_56),
.A2(n_59),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_56),
.A2(n_59),
.B1(n_215),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_56),
.A2(n_59),
.B1(n_224),
.B2(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_59),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_60),
.B(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_63),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_64),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_68),
.A2(n_69),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_321),
.B(n_327),
.Y(n_71)
);

OAI321xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_294),
.A3(n_314),
.B1(n_319),
.B2(n_320),
.C(n_336),
.Y(n_72)
);

AOI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_240),
.A3(n_282),
.B1(n_288),
.B2(n_293),
.C(n_337),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_197),
.C(n_236),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_167),
.B(n_196),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_146),
.B(n_166),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_127),
.B(n_145),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_116),
.B(n_126),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_102),
.B(n_115),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_81),
.B(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_85),
.A2(n_86),
.B1(n_143),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_106),
.B1(n_107),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_101),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_110),
.B(n_114),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_107),
.B1(n_124),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_106),
.A2(n_107),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_106),
.A2(n_107),
.B1(n_178),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_106),
.A2(n_107),
.B1(n_212),
.B2(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_106),
.A2(n_107),
.B(n_222),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_121),
.C(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.CI(n_136),
.CON(n_129),
.SN(n_129)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_160),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_162),
.C(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_158),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_161),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_181),
.C(n_182),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_190),
.C(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_187),
.A2(n_189),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_198),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_217),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_199),
.B(n_217),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.C(n_216),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_216),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_234),
.B2(n_235),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_225),
.C(n_235),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_223),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_230),
.C(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_228),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_238),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_259),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_241),
.B(n_259),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.C(n_258),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_242),
.A2(n_243),
.B1(n_252),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_248),
.C(n_251),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_254),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_253),
.A2(n_275),
.B(n_278),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_255),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_280),
.B2(n_281),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_272),
.C(n_281),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_267),
.B(n_270),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_270),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_270),
.A2(n_296),
.B1(n_305),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_278),
.B2(n_279),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_289),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_307),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_305),
.C(n_306),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_298),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_303),
.C(n_304),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_309),
.C(n_313),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_301),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_326),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_323),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule