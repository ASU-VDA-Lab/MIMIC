module fake_jpeg_10611_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_41),
.CON(n_63),
.SN(n_63)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_29),
.B1(n_30),
.B2(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_15),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_33),
.B1(n_18),
.B2(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_107)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_55),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_61),
.B(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_29),
.B1(n_21),
.B2(n_30),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_71),
.B(n_28),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_21),
.B1(n_30),
.B2(n_18),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_45),
.B1(n_36),
.B2(n_47),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_96)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_84),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_47),
.B1(n_44),
.B2(n_41),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_93),
.B1(n_94),
.B2(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_44),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_36),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_95),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_33),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_14),
.B(n_12),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_92),
.A2(n_97),
.B1(n_90),
.B2(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_38),
.B1(n_40),
.B2(n_20),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_27),
.B1(n_35),
.B2(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_103),
.B1(n_90),
.B2(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_32),
.B1(n_25),
.B2(n_35),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_0),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_31),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_52),
.A2(n_34),
.B1(n_16),
.B2(n_39),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_31),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_66),
.C(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_52),
.A2(n_34),
.B1(n_31),
.B2(n_2),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_0),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_34),
.B1(n_15),
.B2(n_14),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_68),
.B(n_62),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_116),
.A2(n_120),
.B(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_91),
.B(n_99),
.Y(n_155)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_128),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_14),
.A3(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_142),
.B1(n_130),
.B2(n_120),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_94),
.B1(n_105),
.B2(n_93),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_0),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_146),
.B1(n_111),
.B2(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_166),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_150),
.B(n_152),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_110),
.C(n_79),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_162),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_160),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_127),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_78),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_167),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_115),
.B(n_113),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_165),
.B(n_172),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_179),
.B1(n_119),
.B2(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_112),
.B1(n_98),
.B2(n_85),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_170),
.B1(n_176),
.B2(n_116),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_134),
.C(n_135),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_10),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_88),
.B1(n_86),
.B2(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_133),
.B1(n_123),
.B2(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_88),
.B1(n_106),
.B2(n_86),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_177),
.B1(n_137),
.B2(n_117),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_114),
.B1(n_83),
.B2(n_109),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_121),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_185),
.Y(n_219)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_200),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_189),
.B1(n_198),
.B2(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_196),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_116),
.B1(n_125),
.B2(n_121),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_201),
.B1(n_204),
.B2(n_210),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_139),
.B(n_89),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_203),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_150),
.B1(n_149),
.B2(n_166),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_102),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_179),
.B1(n_161),
.B2(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_102),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_165),
.C(n_151),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_153),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_181),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_226),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_220),
.B1(n_232),
.B2(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_230),
.C(n_242),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_152),
.B1(n_169),
.B2(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_155),
.C(n_180),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_207),
.B(n_213),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_209),
.C(n_162),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_193),
.A2(n_169),
.B1(n_174),
.B2(n_162),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_174),
.B1(n_175),
.B2(n_153),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_175),
.B1(n_163),
.B2(n_10),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_6),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_9),
.B1(n_190),
.B2(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_196),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_242),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_182),
.C(n_199),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_205),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_255),
.C(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_187),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_211),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_198),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_228),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_235),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_186),
.B(n_210),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_237),
.B(n_217),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_184),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_198),
.C(n_202),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_224),
.C(n_231),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_222),
.B(n_238),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_275),
.B(n_277),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_282),
.B1(n_271),
.B2(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_254),
.C(n_243),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_258),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_241),
.B1(n_238),
.B2(n_226),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_227),
.C(n_223),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_285),
.C(n_248),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_223),
.C(n_198),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_289),
.C(n_292),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_251),
.B1(n_265),
.B2(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_293),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_255),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_284),
.C(n_285),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_225),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_236),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_300),
.B1(n_280),
.B2(n_277),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_278),
.A2(n_253),
.B1(n_244),
.B2(n_250),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_311),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_266),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_309),
.C(n_310),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_266),
.C(n_267),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_289),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_267),
.C(n_270),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_286),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_319),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_293),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_322),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_269),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_326),
.B(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_312),
.B1(n_272),
.B2(n_287),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_307),
.C(n_310),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_291),
.B1(n_272),
.B2(n_250),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_225),
.B1(n_268),
.B2(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_306),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_328),
.C(n_327),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_328),
.B(n_336),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_332),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_329),
.Y(n_341)
);


endmodule