module fake_jpeg_22162_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_44),
.B1(n_49),
.B2(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_16),
.B2(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_60),
.Y(n_86)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_63),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_34),
.B1(n_29),
.B2(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_68),
.B1(n_70),
.B2(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_69),
.C(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_33),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_82),
.Y(n_105)
);

AO21x2_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_26),
.B(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_51),
.B1(n_37),
.B2(n_31),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_16),
.B1(n_27),
.B2(n_19),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_34),
.B(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_27),
.B1(n_19),
.B2(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_74),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_30),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_51),
.B1(n_31),
.B2(n_28),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_30),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_94),
.B1(n_106),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_100),
.B1(n_107),
.B2(n_57),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_28),
.B(n_20),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_104),
.B1(n_106),
.B2(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_81),
.B1(n_69),
.B2(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_31),
.B1(n_15),
.B2(n_14),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_118),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_123),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_125),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_129),
.C(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_85),
.Y(n_117)
);

NAND2x1_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_84),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_62),
.B(n_61),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_92),
.B(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_75),
.B(n_62),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_79),
.C(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_80),
.B1(n_73),
.B2(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_1),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_99),
.B(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_66),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_66),
.C(n_74),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_158),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_148),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_147),
.B(n_150),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_101),
.B(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_99),
.B(n_94),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_118),
.B(n_110),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_3),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_154),
.C(n_155),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_87),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_14),
.C(n_13),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_163),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_125),
.B(n_118),
.C(n_132),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_171),
.B1(n_176),
.B2(n_155),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_154),
.C(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_157),
.A2(n_113),
.B1(n_132),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_173),
.B1(n_149),
.B2(n_144),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_113),
.B1(n_112),
.B2(n_12),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_112),
.B1(n_12),
.B2(n_5),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_186),
.C(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_148),
.B1(n_139),
.B2(n_137),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_153),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_189),
.B1(n_160),
.B2(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_140),
.B1(n_156),
.B2(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_174),
.B1(n_164),
.B2(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_170),
.C(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_200),
.C(n_9),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_160),
.C(n_8),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_190),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_3),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_181),
.B(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_8),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_8),
.B(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_10),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_208),
.C(n_211),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_10),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_212),
.C(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_204),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_218),
.B(n_10),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_222),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_11),
.B(n_229),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_11),
.Y(n_233)
);


endmodule