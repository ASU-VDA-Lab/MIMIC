module fake_jpeg_18084_n_58 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_3),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_34),
.B(n_1),
.C(n_5),
.Y(n_43)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_6),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_11),
.B(n_12),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_13),
.B(n_14),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_15),
.C(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_22),
.Y(n_58)
);


endmodule