module fake_jpeg_7412_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_39),
.B1(n_49),
.B2(n_48),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_50),
.B1(n_46),
.B2(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_74),
.B1(n_76),
.B2(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_4),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_4),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_20),
.C(n_21),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_85),
.B(n_86),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_71),
.B(n_62),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_71),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_83),
.B(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_22),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_25),
.B(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_99),
.B1(n_84),
.B2(n_88),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_87),
.A3(n_91),
.B1(n_90),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_27),
.C(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_30),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_34),
.Y(n_106)
);


endmodule