module fake_jpeg_1357_n_168 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_61),
.Y(n_77)
);

BUFx12f_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_48),
.B1(n_50),
.B2(n_55),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_57),
.C(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_55),
.B1(n_47),
.B2(n_45),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_54),
.B1(n_51),
.B2(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_1),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_58),
.CI(n_2),
.CON(n_84),
.SN(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_59),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_116),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_4),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_113),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_8),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_10),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_20),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_92),
.B1(n_12),
.B2(n_11),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_137),
.B1(n_31),
.B2(n_34),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_29),
.C(n_14),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_12),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_16),
.B(n_19),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_108),
.B1(n_23),
.B2(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_42),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_124),
.C(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_35),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_132),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_156),
.B1(n_147),
.B2(n_150),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_142),
.B1(n_146),
.B2(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_159),
.B1(n_134),
.B2(n_125),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

NAND2x1p5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_158),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_157),
.B1(n_145),
.B2(n_144),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_162),
.C(n_134),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_37),
.C(n_38),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_41),
.Y(n_168)
);


endmodule