module fake_jpeg_3103_n_94 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_37),
.Y(n_40)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2x1_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_23),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_0),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_0),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_23),
.C(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_43),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_19),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_60),
.B1(n_57),
.B2(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_74),
.B1(n_16),
.B2(n_18),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_4),
.B(n_5),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_7),
.C(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_12),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_6),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_82),
.B(n_74),
.C(n_20),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_78),
.B1(n_67),
.B2(n_76),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_85),
.B1(n_86),
.B2(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_83),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_80),
.C(n_21),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_93),
.Y(n_94)
);


endmodule