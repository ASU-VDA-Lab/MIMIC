module fake_jpeg_5580_n_320 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_11),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_38),
.B(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_42),
.B(n_46),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_16),
.B(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_50),
.B1(n_27),
.B2(n_22),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_60),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_29),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_59),
.B(n_61),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_69),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_89),
.B1(n_93),
.B2(n_20),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_71),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_75),
.B(n_81),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_23),
.Y(n_77)
);

OAI222xp33_ASAP7_75t_L g127 ( 
.A1(n_77),
.A2(n_24),
.B1(n_31),
.B2(n_19),
.C1(n_8),
.C2(n_12),
.Y(n_127)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_34),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_27),
.B1(n_17),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_84),
.B1(n_92),
.B2(n_15),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_23),
.B1(n_30),
.B2(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_34),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_34),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_33),
.B1(n_25),
.B2(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_33),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_99),
.B1(n_22),
.B2(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_100),
.B1(n_20),
.B2(n_16),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_22),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_18),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_127),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_123),
.B(n_63),
.C(n_61),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_112),
.B1(n_117),
.B2(n_111),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_52),
.B1(n_62),
.B2(n_76),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_119),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_77),
.B(n_99),
.C(n_64),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_64),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_135),
.C(n_101),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_95),
.A3(n_72),
.B1(n_90),
.B2(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_57),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_139),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_137),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_59),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_24),
.Y(n_199)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_149),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_60),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_148),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_123),
.B1(n_127),
.B2(n_109),
.Y(n_143)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_53),
.B1(n_63),
.B2(n_67),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_113),
.B1(n_128),
.B2(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_58),
.B1(n_71),
.B2(n_69),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_31),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_52),
.B1(n_54),
.B2(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_78),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_153),
.Y(n_180)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_160),
.B1(n_161),
.B2(n_128),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_24),
.B(n_31),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_19),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_108),
.B1(n_114),
.B2(n_105),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_62),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_118),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_175),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_201),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_199),
.B1(n_149),
.B2(n_140),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_101),
.C(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_196),
.C(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_113),
.B1(n_128),
.B2(n_24),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_137),
.B(n_133),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_189),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_68),
.B1(n_65),
.B2(n_24),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_192),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_31),
.C(n_19),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_130),
.A2(n_31),
.B1(n_19),
.B2(n_8),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_31),
.C(n_122),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_218),
.B(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_139),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_134),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_210),
.B(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_187),
.B1(n_193),
.B2(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_155),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_138),
.C(n_131),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_151),
.B1(n_153),
.B2(n_152),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_151),
.C(n_162),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_151),
.B(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_0),
.C(n_2),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_2),
.C(n_3),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_186),
.C(n_196),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_185),
.B(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_7),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_172),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_247),
.C(n_208),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_250),
.Y(n_257)
);

OAI322xp33_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_172),
.A3(n_171),
.B1(n_190),
.B2(n_175),
.C1(n_191),
.C2(n_188),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_203),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_252),
.CI(n_216),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_202),
.C(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_214),
.A2(n_177),
.B1(n_184),
.B2(n_169),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_205),
.B1(n_206),
.B2(n_221),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_215),
.C(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_211),
.A2(n_195),
.B1(n_177),
.B2(n_169),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_253),
.A2(n_204),
.B1(n_220),
.B2(n_219),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_217),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_264),
.C(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_212),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_263),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_236),
.B1(n_243),
.B2(n_232),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_204),
.B1(n_167),
.B2(n_176),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_246),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_238),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_230),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_233),
.B(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_280),
.C(n_283),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_269),
.A2(n_250),
.B1(n_237),
.B2(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

FAx1_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_234),
.CI(n_229),
.CON(n_278),
.SN(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_234),
.C(n_240),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_238),
.B1(n_235),
.B2(n_231),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_266),
.Y(n_286)
);

NOR4xp25_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_256),
.C(n_259),
.D(n_270),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_3),
.C(n_4),
.Y(n_283)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_291),
.B(n_279),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_258),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_294),
.B(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_265),
.C(n_261),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_272),
.B(n_276),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_258),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_293),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_260),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_268),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_7),
.Y(n_309)
);

NAND2xp67_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_282),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_300),
.B(n_301),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_279),
.B(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_285),
.B(n_289),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_275),
.B1(n_283),
.B2(n_281),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_290),
.B1(n_5),
.B2(n_4),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_9),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_303),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_305),
.Y(n_317)
);

OAI211xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_310),
.B(n_308),
.C(n_302),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_313),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_12),
.Y(n_320)
);


endmodule