module fake_jpeg_13177_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_49),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_1),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_80),
.B1(n_33),
.B2(n_35),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_17),
.B1(n_23),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_77),
.B1(n_81),
.B2(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_16),
.B1(n_30),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_66),
.B1(n_20),
.B2(n_21),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_16),
.B1(n_30),
.B2(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_22),
.Y(n_101)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_23),
.B1(n_30),
.B2(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_23),
.B1(n_16),
.B2(n_33),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_86),
.Y(n_132)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_97),
.Y(n_119)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_90),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_143)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_55),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_104),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_22),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_65),
.B(n_41),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_42),
.C(n_53),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_22),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_79),
.B(n_73),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_114),
.B(n_86),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_66),
.B1(n_33),
.B2(n_34),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_87),
.B1(n_100),
.B2(n_92),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_76),
.A3(n_57),
.B1(n_53),
.B2(n_35),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_86),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_100),
.C(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_104),
.B1(n_94),
.B2(n_83),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_148),
.B(n_42),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_20),
.B1(n_29),
.B2(n_21),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_27),
.B1(n_41),
.B2(n_20),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_91),
.A2(n_109),
.B1(n_86),
.B2(n_103),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_91),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_150),
.B(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_152),
.A2(n_153),
.B1(n_166),
.B2(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_107),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_168),
.B(n_182),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_159),
.B(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_95),
.B1(n_112),
.B2(n_108),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_106),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_57),
.B1(n_89),
.B2(n_39),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_84),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_175),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_84),
.C(n_90),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_178),
.C(n_129),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_90),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_26),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_102),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_117),
.C(n_41),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_138),
.B1(n_142),
.B2(n_147),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_121),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_102),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_19),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_13),
.B(n_9),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_29),
.B(n_21),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_26),
.B(n_2),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_124),
.B(n_137),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_185),
.A2(n_186),
.B(n_165),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_140),
.B(n_145),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_212),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_202),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_118),
.B1(n_143),
.B2(n_134),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_204),
.B1(n_209),
.B2(n_189),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_152),
.A2(n_118),
.B1(n_138),
.B2(n_147),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_201),
.B1(n_206),
.B2(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_213),
.C(n_149),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_131),
.B1(n_122),
.B2(n_19),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

AOI211xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_27),
.B(n_122),
.C(n_131),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_129),
.B1(n_126),
.B2(n_28),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_208),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_153),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_26),
.C(n_19),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_19),
.B1(n_9),
.B2(n_15),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_216),
.B1(n_218),
.B2(n_10),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_163),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

AOI22x1_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_155),
.B1(n_183),
.B2(n_168),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_228),
.B1(n_236),
.B2(n_196),
.Y(n_248)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_156),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_167),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_157),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_230),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_176),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_240),
.B(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_149),
.C(n_170),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_160),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_241),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_151),
.B1(n_179),
.B2(n_177),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_181),
.B(n_175),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_214),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_213),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_10),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_10),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_32),
.C(n_2),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_255),
.B1(n_223),
.B2(n_240),
.Y(n_276)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_224),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_229),
.A2(n_202),
.B1(n_184),
.B2(n_194),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_198),
.B1(n_201),
.B2(n_184),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_260),
.B1(n_32),
.B2(n_3),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_190),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_187),
.B1(n_216),
.B2(n_186),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_208),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_233),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_217),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_241),
.Y(n_268)
);

XOR2x2_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_204),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_238),
.B1(n_239),
.B2(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_250),
.B1(n_268),
.B2(n_6),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_190),
.B(n_212),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_256),
.B(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_280),
.B(n_4),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_206),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_258),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_264),
.B(n_271),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_32),
.C(n_2),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_288),
.C(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_32),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_32),
.C(n_3),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_263),
.B1(n_253),
.B2(n_260),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_1),
.C(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_296),
.A2(n_306),
.B(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_304),
.C(n_301),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_309),
.B(n_277),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_250),
.B(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_4),
.C(n_5),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_5),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_322),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_291),
.B1(n_274),
.B2(n_283),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_316),
.B1(n_318),
.B2(n_295),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_298),
.B(n_279),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_310),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_296),
.A2(n_281),
.B1(n_292),
.B2(n_286),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_305),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_287),
.B(n_288),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_324),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_303),
.A2(n_5),
.B(n_6),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_297),
.B(n_308),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_327),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_318),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_329),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_332),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_297),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_321),
.B(n_300),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_336),
.A2(n_313),
.B(n_312),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_342),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_323),
.C(n_321),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_341),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_313),
.B(n_322),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_336),
.C(n_326),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_345),
.A2(n_344),
.B(n_340),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_325),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_349),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_304),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_347),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_352),
.B(n_350),
.CI(n_343),
.CON(n_353),
.SN(n_353)
);

OAI311xp33_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_7),
.A3(n_8),
.B1(n_346),
.C1(n_352),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_353),
.C(n_7),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_7),
.Y(n_356)
);


endmodule