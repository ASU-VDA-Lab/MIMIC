module real_jpeg_21419_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_21),
.A3(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_1),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_87)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_5),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_49),
.B(n_59),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_10),
.B(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_36),
.B1(n_40),
.B2(n_87),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

BUFx3_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_68),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_67),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_43),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_43),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_30),
.C(n_35),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_17),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_18),
.A2(n_23),
.B1(n_28),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_18),
.A2(n_23),
.B1(n_26),
.B2(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_21),
.A2(n_22),
.B(n_53),
.C(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_53),
.Y(n_85)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_25),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_34),
.B(n_50),
.C(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_50),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_35),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_36),
.A2(n_40),
.B1(n_74),
.B2(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_96),
.B(n_101),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_83),
.B(n_95),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_76),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_88),
.B(n_94),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);


endmodule