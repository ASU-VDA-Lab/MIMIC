module fake_jpeg_5862_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_52),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_30),
.B1(n_15),
.B2(n_19),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_52),
.B1(n_22),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_28),
.C(n_19),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_69),
.B1(n_81),
.B2(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_31),
.B1(n_20),
.B2(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_21),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_40),
.B(n_32),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_76),
.B(n_21),
.C(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_83),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_25),
.B1(n_16),
.B2(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_21),
.B1(n_6),
.B2(n_12),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_32),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_23),
.B1(n_29),
.B2(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_56),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_29),
.B1(n_23),
.B2(n_36),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_99),
.B1(n_75),
.B2(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_58),
.C(n_47),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_106),
.C(n_79),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_49),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_91),
.CI(n_95),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_0),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_102),
.B1(n_79),
.B2(n_74),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_40),
.B1(n_61),
.B2(n_36),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_78),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_81),
.Y(n_111)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_32),
.C(n_38),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_111),
.B1(n_114),
.B2(n_99),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_73),
.B1(n_82),
.B2(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_125),
.B1(n_70),
.B2(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_84),
.B1(n_76),
.B2(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_88),
.B(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_76),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_99),
.B1(n_97),
.B2(n_86),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_67),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_137),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_125),
.B1(n_110),
.B2(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_103),
.B1(n_70),
.B2(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_139),
.B1(n_111),
.B2(n_108),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_149),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_100),
.B(n_103),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_136),
.B(n_138),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_93),
.B(n_87),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_104),
.B1(n_43),
.B2(n_44),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_83),
.B(n_32),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_147),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_0),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_38),
.B(n_23),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_151),
.B(n_128),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_140),
.B1(n_144),
.B2(n_139),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_114),
.B1(n_111),
.B2(n_109),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_168),
.B(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_115),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_120),
.C(n_144),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_135),
.B(n_145),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_176),
.B(n_154),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_129),
.B(n_143),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_129),
.A3(n_137),
.B1(n_115),
.B2(n_143),
.C1(n_132),
.C2(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_188),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_115),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_160),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_150),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_138),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_151),
.C(n_148),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_189),
.C(n_162),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_108),
.C(n_147),
.Y(n_189)
);

BUFx12f_ASAP7_75t_SL g195 ( 
.A(n_182),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_196),
.B(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_157),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_152),
.B(n_166),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_203),
.C(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_172),
.B1(n_167),
.B2(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_172),
.B1(n_167),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_173),
.B1(n_185),
.B2(n_176),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_154),
.C(n_38),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_184),
.C(n_187),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_214),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_189),
.B(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_211),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_3),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_8),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_174),
.C(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_194),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_204),
.C(n_203),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_198),
.B1(n_202),
.B2(n_61),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_7),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_44),
.B(n_43),
.C(n_23),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_13),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_29),
.B1(n_4),
.B2(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_219),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_211),
.B(n_218),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_233),
.B(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_8),
.Y(n_241)
);

FAx1_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_219),
.CI(n_4),
.CON(n_233),
.SN(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_6),
.C(n_7),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_222),
.B(n_10),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_237),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_228),
.B1(n_227),
.B2(n_11),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_240),
.B(n_243),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_8),
.B(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_231),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_12),
.C(n_13),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_245),
.B1(n_233),
.B2(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_234),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_249),
.B(n_247),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_251),
.Y(n_252)
);


endmodule