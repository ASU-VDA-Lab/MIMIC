module real_aes_9149_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g511 ( .A1(n_0), .A2(n_171), .B(n_512), .C(n_515), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_1), .B(n_462), .Y(n_516) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
NAND3xp33_ASAP7_75t_SL g765 ( .A(n_2), .B(n_111), .C(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g183 ( .A(n_3), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_4), .B(n_143), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_5), .A2(n_435), .B(n_456), .Y(n_455) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_6), .A2(n_163), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_7), .A2(n_39), .B1(n_137), .B2(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_8), .B(n_163), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_9), .A2(n_727), .B1(n_733), .B2(n_734), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_9), .Y(n_733) );
AND2x6_ASAP7_75t_L g155 ( .A(n_10), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_11), .A2(n_155), .B(n_440), .C(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_12), .B(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g763 ( .A(n_12), .Y(n_763) );
INVx1_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
INVx1_ASAP7_75t_L g176 ( .A(n_14), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_15), .B(n_141), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_16), .B(n_143), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_17), .B(n_129), .Y(n_247) );
AO32x2_ASAP7_75t_L g189 ( .A1(n_18), .A2(n_128), .A3(n_154), .B1(n_163), .B2(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_19), .B(n_137), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_20), .B(n_129), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_21), .A2(n_55), .B1(n_137), .B2(n_192), .Y(n_193) );
AOI22xp33_ASAP7_75t_SL g231 ( .A1(n_22), .A2(n_82), .B1(n_137), .B2(n_141), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_23), .B(n_137), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_24), .A2(n_154), .B(n_440), .C(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_25), .A2(n_60), .B1(n_425), .B2(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_25), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_26), .A2(n_154), .B(n_440), .C(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_28), .B(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_29), .A2(n_435), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_30), .B(n_158), .Y(n_206) );
INVx2_ASAP7_75t_L g139 ( .A(n_31), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_32), .A2(n_438), .B(n_448), .C(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_33), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_34), .B(n_158), .Y(n_217) );
XNOR2x2_ASAP7_75t_SL g747 ( .A(n_35), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_36), .B(n_213), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_37), .A2(n_86), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_37), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_38), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_40), .B(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_41), .B(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_42), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_43), .B(n_143), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_44), .B(n_435), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_45), .A2(n_438), .B(n_442), .C(n_448), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_46), .A2(n_84), .B1(n_482), .B2(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_46), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_47), .B(n_137), .Y(n_166) );
INVx1_ASAP7_75t_L g513 ( .A(n_48), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_49), .A2(n_92), .B1(n_192), .B2(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g443 ( .A(n_50), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_51), .B(n_137), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_52), .B(n_137), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_53), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_54), .B(n_149), .Y(n_170) );
AOI22xp33_ASAP7_75t_SL g245 ( .A1(n_56), .A2(n_61), .B1(n_137), .B2(n_141), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_57), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_58), .B(n_137), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_59), .B(n_137), .Y(n_210) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_60), .A2(n_121), .B1(n_425), .B2(n_426), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_60), .Y(n_425) );
INVx1_ASAP7_75t_L g156 ( .A(n_62), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_63), .B(n_435), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_64), .B(n_462), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_65), .A2(n_149), .B(n_179), .C(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_66), .B(n_137), .Y(n_184) );
INVx1_ASAP7_75t_L g132 ( .A(n_67), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_68), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_69), .B(n_143), .Y(n_480) );
AO32x2_ASAP7_75t_L g227 ( .A1(n_70), .A2(n_154), .A3(n_163), .B1(n_228), .B2(n_232), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_71), .B(n_144), .Y(n_526) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g201 ( .A(n_73), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_74), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_75), .B(n_445), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_76), .A2(n_440), .B(n_448), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_77), .B(n_141), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_78), .Y(n_457) );
INVx1_ASAP7_75t_L g768 ( .A(n_79), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g105 ( .A1(n_80), .A2(n_106), .B1(n_758), .B2(n_769), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_81), .B(n_444), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_83), .B(n_192), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_84), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_85), .B(n_141), .Y(n_205) );
INVx1_ASAP7_75t_L g732 ( .A(n_86), .Y(n_732) );
INVx2_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_88), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_89), .B(n_153), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_90), .B(n_141), .Y(n_167) );
INVx2_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
OR2x2_ASAP7_75t_L g743 ( .A(n_91), .B(n_112), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_93), .A2(n_104), .B1(n_141), .B2(n_142), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_94), .B(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_95), .Y(n_479) );
INVxp67_ASAP7_75t_L g460 ( .A(n_96), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_97), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g501 ( .A(n_98), .Y(n_501) );
INVx1_ASAP7_75t_L g522 ( .A(n_99), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_100), .B(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_101), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_101), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_102), .Y(n_756) );
AND2x2_ASAP7_75t_L g450 ( .A(n_103), .B(n_158), .Y(n_450) );
AO221x2_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_737), .B1(n_744), .B2(n_751), .C(n_755), .Y(n_106) );
OAI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_109), .B(n_116), .Y(n_107) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g119 ( .A(n_111), .Y(n_119) );
INVx2_ASAP7_75t_L g427 ( .A(n_111), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g116 ( .A1(n_112), .A2(n_117), .B1(n_726), .B2(n_735), .C(n_736), .Y(n_116) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g735 ( .A(n_117), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_120), .B1(n_427), .B2(n_428), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g426 ( .A(n_121), .Y(n_426) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_121), .B(n_749), .Y(n_748) );
OR3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_353), .C(n_402), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_268), .C(n_296), .D(n_326), .E(n_340), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_186), .B1(n_218), .B2(n_223), .C(n_234), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_125), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g248 ( .A(n_126), .Y(n_248) );
AND2x2_ASAP7_75t_L g256 ( .A(n_126), .B(n_162), .Y(n_256) );
AND2x2_ASAP7_75t_L g279 ( .A(n_126), .B(n_161), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_126), .B(n_173), .Y(n_294) );
OR2x2_ASAP7_75t_L g303 ( .A(n_126), .B(n_241), .Y(n_303) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_126), .Y(n_306) );
AND2x2_ASAP7_75t_L g414 ( .A(n_126), .B(n_241), .Y(n_414) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_157), .Y(n_126) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_127), .A2(n_174), .B(n_185), .Y(n_173) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_128), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_130), .B(n_131), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_146), .B(n_154), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_143), .Y(n_135) );
INVx3_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_137), .Y(n_503) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
BUFx3_ASAP7_75t_L g230 ( .A(n_138), .Y(n_230) );
AND2x6_ASAP7_75t_L g440 ( .A(n_138), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g142 ( .A(n_139), .Y(n_142) );
INVx1_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx2_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_143), .A2(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
O2A1O1Ixp5_ASAP7_75t_SL g199 ( .A1(n_143), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_143), .B(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_144), .A2(n_153), .B1(n_229), .B2(n_231), .Y(n_228) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
INVx1_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
AND2x2_ASAP7_75t_L g436 ( .A(n_145), .B(n_150), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_145), .Y(n_441) );
O2A1O1Ixp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_152), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_148), .A2(n_171), .B(n_183), .C(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_148), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_152), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_153), .A2(n_171), .B1(n_191), .B2(n_193), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_153), .A2(n_171), .B1(n_244), .B2(n_245), .Y(n_243) );
INVx4_ASAP7_75t_L g514 ( .A(n_153), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_154), .B(n_242), .C(n_243), .Y(n_267) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_155), .A2(n_165), .B(n_168), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_175), .B(n_182), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_155), .A2(n_199), .B(n_203), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_155), .A2(n_209), .B(n_214), .Y(n_208) );
AND2x4_ASAP7_75t_L g435 ( .A(n_155), .B(n_436), .Y(n_435) );
INVx4_ASAP7_75t_SL g449 ( .A(n_155), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_155), .B(n_436), .Y(n_523) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_158), .A2(n_198), .B(n_206), .Y(n_197) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_208), .B(n_217), .Y(n_207) );
INVx2_ASAP7_75t_L g232 ( .A(n_158), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_158), .A2(n_434), .B(n_437), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_158), .A2(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g495 ( .A(n_158), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_159), .B(n_306), .Y(n_362) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
OAI311xp33_ASAP7_75t_L g304 ( .A1(n_160), .A2(n_305), .A3(n_306), .B1(n_307), .C1(n_322), .Y(n_304) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_173), .Y(n_160) );
AND2x2_ASAP7_75t_L g265 ( .A(n_161), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_161), .Y(n_272) );
AND2x2_ASAP7_75t_L g393 ( .A(n_161), .B(n_222), .Y(n_393) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_162), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g249 ( .A(n_162), .B(n_173), .Y(n_249) );
AND2x2_ASAP7_75t_L g301 ( .A(n_162), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g315 ( .A(n_162), .B(n_248), .Y(n_315) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_172), .Y(n_162) );
INVx4_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_163), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_163), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g222 ( .A(n_173), .Y(n_222) );
AND2x2_ASAP7_75t_L g264 ( .A(n_173), .B(n_248), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_179), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_177), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_177), .A2(n_526), .B(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_179), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_180), .A2(n_204), .B(n_205), .Y(n_203) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g445 ( .A(n_181), .Y(n_445) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_194), .Y(n_186) );
OR2x2_ASAP7_75t_L g359 ( .A(n_187), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_187), .B(n_365), .Y(n_376) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_188), .B(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g233 ( .A(n_189), .Y(n_233) );
AND2x2_ASAP7_75t_L g300 ( .A(n_189), .B(n_227), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_189), .B(n_207), .Y(n_311) );
AND2x2_ASAP7_75t_L g320 ( .A(n_189), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_194), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_194), .B(n_261), .Y(n_305) );
INVx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g292 ( .A(n_195), .B(n_251), .Y(n_292) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
INVx2_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
AND2x2_ASAP7_75t_L g319 ( .A(n_196), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
OR2x2_ASAP7_75t_L g336 ( .A(n_197), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_197), .Y(n_399) );
AND2x2_ASAP7_75t_L g238 ( .A(n_207), .B(n_233), .Y(n_238) );
INVx1_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
AND2x2_ASAP7_75t_L g280 ( .A(n_207), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g321 ( .A(n_207), .Y(n_321) );
INVx1_ASAP7_75t_L g337 ( .A(n_207), .Y(n_337) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_207), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_220), .B(n_325), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_220), .A2(n_310), .B1(n_359), .B2(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_221), .A2(n_403), .B(n_405), .C(n_423), .Y(n_402) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AND2x2_ASAP7_75t_L g313 ( .A(n_222), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g324 ( .A(n_222), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_223), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
AND2x2_ASAP7_75t_L g297 ( .A(n_224), .B(n_261), .Y(n_297) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g329 ( .A(n_225), .B(n_320), .Y(n_329) );
AND2x2_ASAP7_75t_L g348 ( .A(n_225), .B(n_262), .Y(n_348) );
AND2x4_ASAP7_75t_L g284 ( .A(n_226), .B(n_258), .Y(n_284) );
AND2x2_ASAP7_75t_L g422 ( .A(n_226), .B(n_398), .Y(n_422) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_227), .Y(n_251) );
INVx1_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
INVx1_ASAP7_75t_L g361 ( .A(n_227), .Y(n_361) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_230), .Y(n_447) );
INVx2_ASAP7_75t_L g515 ( .A(n_230), .Y(n_515) );
INVx1_ASAP7_75t_L g492 ( .A(n_232), .Y(n_492) );
OR2x2_ASAP7_75t_L g252 ( .A(n_233), .B(n_237), .Y(n_252) );
AND2x2_ASAP7_75t_L g261 ( .A(n_233), .B(n_262), .Y(n_261) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_233), .B(n_282), .Y(n_281) );
OAI221xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_239), .B1(n_250), .B2(n_253), .C(n_257), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_258), .B(n_260), .C(n_263), .Y(n_257) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g282 ( .A(n_237), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_237), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_237), .B(n_259), .Y(n_365) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_237), .Y(n_372) );
AND2x2_ASAP7_75t_L g290 ( .A(n_238), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g327 ( .A(n_238), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
INVx2_ASAP7_75t_L g318 ( .A(n_240), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_240), .A2(n_251), .B1(n_368), .B2(n_370), .C1(n_371), .C2(n_373), .Y(n_367) );
AND2x2_ASAP7_75t_L g424 ( .A(n_240), .B(n_393), .Y(n_424) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_248), .Y(n_240) );
INVx1_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
AO21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_246), .Y(n_241) );
INVx3_ASAP7_75t_L g462 ( .A(n_242), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_242), .B(n_482), .Y(n_481) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_242), .A2(n_498), .B(n_505), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_242), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_242), .A2(n_521), .B(n_528), .Y(n_520) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g266 ( .A(n_247), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g352 ( .A(n_249), .B(n_286), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_250), .A2(n_364), .B(n_366), .Y(n_363) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_251), .B(n_258), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_251), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx3_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
OR2x2_ASAP7_75t_L g369 ( .A(n_255), .B(n_291), .Y(n_369) );
AND2x2_ASAP7_75t_L g285 ( .A(n_256), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g323 ( .A(n_256), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_256), .B(n_317), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_256), .B(n_313), .Y(n_339) );
AND2x2_ASAP7_75t_L g343 ( .A(n_256), .B(n_325), .Y(n_343) );
INVxp67_ASAP7_75t_L g275 ( .A(n_258), .Y(n_275) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_260), .A2(n_333), .B1(n_338), .B2(n_339), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_260), .B(n_365), .Y(n_395) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g381 ( .A(n_261), .B(n_372), .Y(n_381) );
AND2x2_ASAP7_75t_L g410 ( .A(n_261), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g415 ( .A(n_261), .B(n_365), .Y(n_415) );
INVx1_ASAP7_75t_L g328 ( .A(n_262), .Y(n_328) );
BUFx2_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx1_ASAP7_75t_L g419 ( .A(n_263), .Y(n_419) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_266), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g278 ( .A(n_266), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
INVx3_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
OR2x2_ASAP7_75t_L g391 ( .A(n_266), .B(n_392), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B(n_276), .C(n_288), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_269), .A2(n_406), .B1(n_413), .B2(n_415), .C(n_416), .Y(n_405) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_283), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_279), .B(n_317), .Y(n_331) );
AND2x2_ASAP7_75t_L g373 ( .A(n_279), .B(n_313), .Y(n_373) );
INVx1_ASAP7_75t_SL g386 ( .A(n_280), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_280), .B(n_334), .Y(n_389) );
INVx1_ASAP7_75t_L g407 ( .A(n_281), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_285), .A2(n_375), .B1(n_377), .B2(n_381), .C(n_382), .Y(n_374) );
AND2x2_ASAP7_75t_L g401 ( .A(n_286), .B(n_393), .Y(n_401) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g385 ( .A(n_287), .Y(n_385) );
AOI21xp33_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_292), .B(n_293), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g356 ( .A(n_291), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
INVx1_ASAP7_75t_L g370 ( .A(n_293), .Y(n_370) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_301), .C(n_304), .Y(n_296) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_297), .A2(n_335), .A3(n_422), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g397 ( .A(n_300), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g418 ( .A(n_300), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_302), .B(n_317), .Y(n_345) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g420 ( .A(n_303), .B(n_317), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B1(n_316), .B2(n_319), .Y(n_307) );
NAND2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_311), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_311), .B(n_334), .Y(n_350) );
AND2x2_ASAP7_75t_L g404 ( .A(n_311), .B(n_399), .Y(n_404) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g379 ( .A(n_315), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OAI32xp33_ASAP7_75t_L g382 ( .A1(n_317), .A2(n_351), .A3(n_383), .B1(n_385), .B2(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g357 ( .A(n_320), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_320), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B(n_330), .C(n_332), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_328), .B(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_329), .A2(n_341), .B1(n_342), .B2(n_343), .C(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g341 ( .A(n_339), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_349), .B2(n_351), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND4xp25_ASAP7_75t_SL g406 ( .A(n_349), .B(n_407), .C(n_408), .D(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND4xp25_ASAP7_75t_SL g353 ( .A(n_354), .B(n_367), .C(n_374), .D(n_387), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_362), .C(n_363), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g384 ( .A(n_360), .Y(n_384) );
INVx2_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
OR2x2_ASAP7_75t_L g417 ( .A(n_372), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_394), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g413 ( .A(n_393), .B(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_396), .B(n_400), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR5x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_599), .C(n_677), .D(n_701), .E(n_718), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_471), .B(n_517), .C(n_576), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_451), .Y(n_431) );
AND2x2_ASAP7_75t_L g530 ( .A(n_432), .B(n_453), .Y(n_530) );
INVx5_ASAP7_75t_SL g558 ( .A(n_432), .Y(n_558) );
AND2x2_ASAP7_75t_L g594 ( .A(n_432), .B(n_579), .Y(n_594) );
OR2x2_ASAP7_75t_L g633 ( .A(n_432), .B(n_452), .Y(n_633) );
OR2x2_ASAP7_75t_L g664 ( .A(n_432), .B(n_555), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_432), .B(n_568), .Y(n_700) );
AND2x2_ASAP7_75t_L g712 ( .A(n_432), .B(n_555), .Y(n_712) );
OR2x6_ASAP7_75t_L g432 ( .A(n_433), .B(n_450), .Y(n_432) );
BUFx2_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_439), .A2(n_449), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_439), .A2(n_449), .B(n_510), .C(n_511), .Y(n_509) );
INVx5_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_446), .C(n_447), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_444), .A2(n_447), .B(n_479), .C(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g711 ( .A(n_451), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g574 ( .A(n_452), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_453), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_453), .Y(n_567) );
INVx3_ASAP7_75t_L g582 ( .A(n_453), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_453), .B(n_463), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_453), .B(n_558), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_453), .B(n_579), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_453), .B(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_L g662 ( .A(n_453), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_453), .B(n_520), .Y(n_676) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_461), .Y(n_453) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_462), .A2(n_508), .B(n_516), .Y(n_507) );
OR2x2_ASAP7_75t_L g568 ( .A(n_463), .B(n_520), .Y(n_568) );
AND2x2_ASAP7_75t_L g579 ( .A(n_463), .B(n_555), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_463), .B(n_582), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_463), .B(n_520), .Y(n_614) );
INVx1_ASAP7_75t_SL g626 ( .A(n_463), .Y(n_626) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g519 ( .A(n_464), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_464), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
AND2x2_ASAP7_75t_L g539 ( .A(n_473), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_473), .B(n_496), .Y(n_543) );
AND2x2_ASAP7_75t_L g546 ( .A(n_473), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_473), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g571 ( .A(n_473), .B(n_562), .Y(n_571) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_473), .Y(n_590) );
AND2x2_ASAP7_75t_L g611 ( .A(n_473), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g621 ( .A(n_473), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g667 ( .A(n_473), .B(n_550), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_473), .B(n_573), .Y(n_694) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g564 ( .A(n_474), .Y(n_564) );
AND2x2_ASAP7_75t_L g630 ( .A(n_474), .B(n_562), .Y(n_630) );
AND2x2_ASAP7_75t_L g714 ( .A(n_474), .B(n_582), .Y(n_714) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_481), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_483), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_483), .Y(n_703) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
AND2x2_ASAP7_75t_L g533 ( .A(n_484), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g542 ( .A(n_484), .B(n_540), .Y(n_542) );
INVx5_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
AND2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_507), .Y(n_573) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_484), .Y(n_610) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
AOI21xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_488), .B(n_492), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g651 ( .A(n_496), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_496), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g684 ( .A(n_496), .B(n_550), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_496), .A2(n_607), .B(n_714), .C(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
BUFx2_ASAP7_75t_L g534 ( .A(n_497), .Y(n_534) );
INVx2_ASAP7_75t_L g538 ( .A(n_497), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
INVx2_ASAP7_75t_L g540 ( .A(n_507), .Y(n_540) );
AND2x2_ASAP7_75t_L g547 ( .A(n_507), .B(n_538), .Y(n_547) );
AND2x2_ASAP7_75t_L g638 ( .A(n_507), .B(n_550), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AOI211x1_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_531), .B(n_544), .C(n_569), .Y(n_517) );
INVx1_ASAP7_75t_L g635 ( .A(n_518), .Y(n_635) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
INVx5_ASAP7_75t_SL g555 ( .A(n_520), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_520), .B(n_625), .Y(n_624) );
AOI311xp33_ASAP7_75t_L g643 ( .A1(n_520), .A2(n_644), .A3(n_646), .B(n_647), .C(n_653), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_520), .A2(n_591), .B(n_679), .C(n_682), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
INVxp67_ASAP7_75t_L g598 ( .A(n_530), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g531 ( .A(n_532), .B(n_535), .C(n_541), .D(n_543), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_532), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_536), .B(n_542), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_536), .B(n_549), .Y(n_669) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_537), .B(n_550), .Y(n_687) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
INVxp67_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
AND2x4_ASAP7_75t_L g549 ( .A(n_540), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g623 ( .A(n_540), .B(n_562), .Y(n_623) );
INVx1_ASAP7_75t_L g650 ( .A(n_540), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_540), .B(n_637), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_541), .B(n_611), .Y(n_631) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_542), .B(n_564), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_542), .B(n_611), .Y(n_710) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B(n_551), .C(n_559), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g563 ( .A(n_547), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g583 ( .A(n_548), .Y(n_583) );
AND2x2_ASAP7_75t_L g560 ( .A(n_549), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_549), .B(n_611), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_549), .B(n_630), .Y(n_654) );
OR2x2_ASAP7_75t_L g570 ( .A(n_550), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g602 ( .A(n_550), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_550), .B(n_562), .Y(n_617) );
AND2x2_ASAP7_75t_L g674 ( .A(n_550), .B(n_630), .Y(n_674) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_550), .Y(n_681) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_552), .A2(n_564), .B1(n_686), .B2(n_688), .C(n_691), .Y(n_685) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g575 ( .A(n_555), .B(n_558), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_555), .B(n_625), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_555), .B(n_582), .Y(n_690) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g675 ( .A(n_557), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g689 ( .A(n_557), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_558), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_558), .B(n_579), .Y(n_586) );
AND2x2_ASAP7_75t_L g656 ( .A(n_558), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_558), .B(n_605), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_558), .B(n_706), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_563), .B(n_565), .Y(n_559) );
INVx2_ASAP7_75t_L g592 ( .A(n_560), .Y(n_592) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
OR2x2_ASAP7_75t_L g616 ( .A(n_564), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_687), .Y(n_719) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AOI21xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_572), .B(n_574), .Y(n_569) );
INVx1_ASAP7_75t_L g723 ( .A(n_570), .Y(n_723) );
INVx2_ASAP7_75t_SL g637 ( .A(n_571), .Y(n_637) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_574), .A2(n_655), .B(n_719), .C(n_720), .Y(n_718) );
OAI322xp33_ASAP7_75t_SL g587 ( .A1(n_575), .A2(n_588), .A3(n_591), .B1(n_592), .B2(n_593), .C1(n_595), .C2(n_598), .Y(n_587) );
INVx2_ASAP7_75t_L g607 ( .A(n_575), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_583), .B1(n_584), .B2(n_586), .C(n_587), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp33_ASAP7_75t_SL g653 ( .A1(n_578), .A2(n_654), .B1(n_655), .B2(n_658), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_579), .B(n_582), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g652 ( .A(n_581), .B(n_614), .Y(n_652) );
INVx1_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_586), .A2(n_696), .B(n_698), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_621), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp67_ASAP7_75t_SL g649 ( .A(n_590), .B(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g706 ( .A(n_591), .Y(n_706) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_600), .B(n_627), .C(n_643), .D(n_659), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_608), .C(n_620), .Y(n_600) );
INVx1_ASAP7_75t_L g692 ( .A(n_601), .Y(n_692) );
AND2x2_ASAP7_75t_L g640 ( .A(n_602), .B(n_623), .Y(n_640) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_607), .B(n_642), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_613), .B1(n_616), .B2(n_618), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_610), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_611), .A2(n_650), .B(n_673), .C(n_675), .Y(n_672) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g657 ( .A(n_614), .Y(n_657) );
INVx1_ASAP7_75t_L g717 ( .A(n_615), .Y(n_717) );
NAND2xp33_ASAP7_75t_SL g707 ( .A(n_616), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g646 ( .A(n_625), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B(n_632), .C(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_639), .B2(n_641), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_637), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_642), .B(n_663), .Y(n_725) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_651), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_672), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_675), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_685), .C(n_695), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_704), .C(n_713), .Y(n_701) );
INVx1_ASAP7_75t_L g722 ( .A(n_702), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_709), .B2(n_711), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g736 ( .A(n_726), .Y(n_736) );
INVx1_ASAP7_75t_L g734 ( .A(n_727), .Y(n_734) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g752 ( .A(n_741), .Y(n_752) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_743), .Y(n_754) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_743), .Y(n_757) );
XOR2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_SL g769 ( .A(n_760), .Y(n_769) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule