module real_aes_7671_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g270 ( .A1(n_0), .A2(n_271), .B(n_272), .C(n_275), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_1), .B(n_212), .Y(n_276) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_3), .B(n_182), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_4), .A2(n_152), .B(n_155), .C(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_5), .A2(n_172), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_6), .A2(n_172), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_7), .B(n_212), .Y(n_525) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_8), .A2(n_139), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_9), .A2(n_459), .B1(n_462), .B2(n_463), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_9), .Y(n_463) );
AND2x6_ASAP7_75t_L g152 ( .A(n_10), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_11), .A2(n_152), .B(n_155), .C(n_158), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_12), .A2(n_47), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_12), .Y(n_460) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_13), .B(n_42), .Y(n_450) );
INVx1_ASAP7_75t_L g495 ( .A(n_14), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_15), .B(n_162), .Y(n_481) );
INVx1_ASAP7_75t_L g144 ( .A(n_16), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_17), .B(n_182), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_18), .A2(n_160), .B(n_503), .C(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_19), .B(n_212), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_20), .B(n_236), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_21), .A2(n_155), .B(n_199), .C(n_232), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_22), .A2(n_164), .B(n_274), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_23), .B(n_162), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_24), .B(n_162), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_25), .Y(n_553) );
INVx1_ASAP7_75t_L g545 ( .A(n_26), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_27), .A2(n_155), .B(n_195), .C(n_199), .Y(n_194) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_28), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_29), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_30), .B(n_454), .Y(n_455) );
INVx1_ASAP7_75t_L g536 ( .A(n_31), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_32), .A2(n_172), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g150 ( .A(n_33), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_34), .A2(n_174), .B(n_185), .C(n_220), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_35), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_36), .A2(n_274), .B(n_522), .C(n_524), .Y(n_521) );
INVxp67_ASAP7_75t_L g537 ( .A(n_37), .Y(n_537) );
OAI321xp33_ASAP7_75t_L g123 ( .A1(n_38), .A2(n_124), .A3(n_446), .B1(n_451), .B2(n_452), .C(n_455), .Y(n_123) );
INVx1_ASAP7_75t_L g451 ( .A(n_38), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_39), .B(n_197), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g520 ( .A(n_40), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_41), .A2(n_155), .B(n_199), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_42), .B(n_109), .Y(n_108) );
AOI222xp33_ASAP7_75t_SL g457 ( .A1(n_43), .A2(n_458), .B1(n_464), .B2(n_737), .C1(n_738), .C2(n_742), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_44), .A2(n_275), .B(n_493), .C(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_45), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_46), .Y(n_167) );
INVx1_ASAP7_75t_L g461 ( .A(n_47), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_48), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_49), .B(n_172), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_50), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_51), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_52), .A2(n_174), .B(n_176), .C(n_185), .Y(n_173) );
INVx1_ASAP7_75t_L g273 ( .A(n_53), .Y(n_273) );
INVx1_ASAP7_75t_L g177 ( .A(n_54), .Y(n_177) );
INVx1_ASAP7_75t_L g510 ( .A(n_55), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_56), .B(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_57), .A2(n_60), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_57), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_58), .Y(n_239) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_59), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_60), .Y(n_127) );
INVx1_ASAP7_75t_L g153 ( .A(n_61), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_62), .B(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_63), .B(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_64), .A2(n_206), .B(n_208), .C(n_210), .Y(n_205) );
INVx1_ASAP7_75t_L g143 ( .A(n_65), .Y(n_143) );
INVx1_ASAP7_75t_SL g523 ( .A(n_66), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_67), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_68), .B(n_182), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_69), .B(n_212), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_70), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g556 ( .A(n_71), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_72), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_73), .B(n_179), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_74), .A2(n_155), .B(n_185), .C(n_246), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_75), .Y(n_204) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_77), .A2(n_172), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_78), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_79), .A2(n_172), .B(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_80), .A2(n_104), .B1(n_117), .B2(n_746), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_81), .A2(n_230), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g501 ( .A(n_82), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_83), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_84), .B(n_178), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_85), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_86), .A2(n_172), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g504 ( .A(n_87), .Y(n_504) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g480 ( .A(n_89), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_90), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_91), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
OR2x2_ASAP7_75t_L g447 ( .A(n_92), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g467 ( .A(n_92), .B(n_449), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_93), .A2(n_155), .B(n_185), .C(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_94), .B(n_172), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_95), .Y(n_221) );
INVxp67_ASAP7_75t_L g209 ( .A(n_96), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_97), .B(n_139), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_98), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g247 ( .A(n_100), .Y(n_247) );
INVx2_ASAP7_75t_L g513 ( .A(n_101), .Y(n_513) );
AND2x2_ASAP7_75t_L g188 ( .A(n_102), .B(n_187), .Y(n_188) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_SL g746 ( .A(n_105), .Y(n_746) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g449 ( .A(n_112), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g736 ( .A(n_113), .B(n_449), .Y(n_736) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_113), .B(n_448), .Y(n_744) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_456), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g745 ( .A(n_122), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_124), .B(n_453), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22x1_ASAP7_75t_SL g738 ( .A1(n_129), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_738) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_130), .A2(n_465), .B1(n_468), .B2(n_734), .Y(n_464) );
OR3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_344), .C(n_409), .Y(n_130) );
NAND4xp25_ASAP7_75t_SL g131 ( .A(n_132), .B(n_285), .C(n_311), .D(n_334), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_213), .B1(n_254), .B2(n_261), .C(n_277), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_134), .A2(n_278), .B1(n_302), .B2(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_189), .Y(n_134) );
INVx1_ASAP7_75t_SL g338 ( .A(n_135), .Y(n_338) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
OR2x2_ASAP7_75t_L g259 ( .A(n_136), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g280 ( .A(n_136), .B(n_190), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_136), .B(n_200), .Y(n_293) );
AND2x2_ASAP7_75t_L g310 ( .A(n_136), .B(n_169), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_136), .B(n_257), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_136), .B(n_309), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_136), .B(n_189), .Y(n_431) );
AOI211xp5_ASAP7_75t_SL g442 ( .A1(n_136), .A2(n_348), .B(n_443), .C(n_444), .Y(n_442) );
INVx5_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_137), .B(n_190), .Y(n_314) );
AND2x2_ASAP7_75t_L g317 ( .A(n_137), .B(n_191), .Y(n_317) );
OR2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_190), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_137), .B(n_200), .Y(n_371) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_145), .B(n_166), .Y(n_137) );
INVx3_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_138), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_138), .A2(n_244), .B(n_252), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_138), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_138), .B(n_484), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_138), .B(n_548), .Y(n_547) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_138), .A2(n_552), .B(n_558), .Y(n_551) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_139), .A2(n_193), .B(n_194), .Y(n_192) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_141), .B(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_147), .A2(n_477), .B(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_147), .A2(n_187), .B(n_542), .C(n_543), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_147), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g172 ( .A(n_148), .B(n_152), .Y(n_172) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
INVx4_ASAP7_75t_SL g186 ( .A(n_152), .Y(n_186) );
BUFx3_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
INVx5_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_156), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_163), .Y(n_158) );
INVx5_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_160), .B(n_495), .Y(n_494) );
INVx4_ASAP7_75t_L g274 ( .A(n_162), .Y(n_274) );
INVx2_ASAP7_75t_L g493 ( .A(n_162), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_163), .A2(n_196), .B(n_198), .Y(n_195) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx2_ASAP7_75t_L g530 ( .A(n_168), .Y(n_530) );
INVx5_ASAP7_75t_SL g260 ( .A(n_169), .Y(n_260) );
AND2x2_ASAP7_75t_L g279 ( .A(n_169), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_169), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g365 ( .A(n_169), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g397 ( .A(n_169), .B(n_200), .Y(n_397) );
OR2x2_ASAP7_75t_L g403 ( .A(n_169), .B(n_293), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_169), .B(n_353), .Y(n_412) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_188), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_187), .Y(n_170) );
BUFx2_ASAP7_75t_L g230 ( .A(n_172), .Y(n_230) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_175), .A2(n_186), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_175), .A2(n_186), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_175), .A2(n_186), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_175), .A2(n_186), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_175), .A2(n_186), .B(n_510), .C(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_175), .A2(n_186), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_175), .A2(n_186), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_181), .C(n_183), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_178), .A2(n_183), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp5_ASAP7_75t_L g479 ( .A1(n_178), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_178), .A2(n_482), .B(n_556), .C(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_182), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g271 ( .A(n_182), .Y(n_271) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_182), .A2(n_207), .B1(n_536), .B2(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_182), .A2(n_235), .B(n_545), .C(n_546), .Y(n_544) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g275 ( .A(n_184), .Y(n_275) );
INVx1_ASAP7_75t_L g505 ( .A(n_184), .Y(n_505) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_187), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
INVx1_ASAP7_75t_L g240 ( .A(n_187), .Y(n_240) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_187), .A2(n_489), .B(n_496), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_200), .Y(n_189) );
AND2x2_ASAP7_75t_L g294 ( .A(n_190), .B(n_260), .Y(n_294) );
INVx1_ASAP7_75t_SL g307 ( .A(n_190), .Y(n_307) );
OR2x2_ASAP7_75t_L g342 ( .A(n_190), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g348 ( .A(n_190), .B(n_200), .Y(n_348) );
AND2x2_ASAP7_75t_L g406 ( .A(n_190), .B(n_257), .Y(n_406) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_191), .B(n_260), .Y(n_333) );
INVx3_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
OR2x2_ASAP7_75t_L g299 ( .A(n_200), .B(n_260), .Y(n_299) );
AND2x2_ASAP7_75t_L g309 ( .A(n_200), .B(n_307), .Y(n_309) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_200), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_200), .B(n_280), .Y(n_366) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_211), .Y(n_200) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_201), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_201), .A2(n_508), .B(n_514), .Y(n_507) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_201), .A2(n_518), .B(n_525), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_206), .A2(n_247), .B(n_248), .C(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_207), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_207), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_210), .B(n_535), .Y(n_534) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_212), .A2(n_267), .B(n_276), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_213), .A2(n_383), .B1(n_385), .B2(n_387), .C(n_390), .Y(n_382) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
AND2x2_ASAP7_75t_L g356 ( .A(n_215), .B(n_337), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_215), .B(n_415), .Y(n_419) );
OR2x2_ASAP7_75t_L g440 ( .A(n_215), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_215), .B(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx5_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
AND2x2_ASAP7_75t_L g364 ( .A(n_216), .B(n_227), .Y(n_364) );
AND2x2_ASAP7_75t_L g425 ( .A(n_216), .B(n_304), .Y(n_425) );
AND2x2_ASAP7_75t_L g438 ( .A(n_216), .B(n_257), .Y(n_438) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_241), .Y(n_225) );
AND2x4_ASAP7_75t_L g264 ( .A(n_226), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g283 ( .A(n_226), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
AND2x2_ASAP7_75t_L g359 ( .A(n_226), .B(n_337), .Y(n_359) );
AND2x2_ASAP7_75t_L g369 ( .A(n_226), .B(n_287), .Y(n_369) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_226), .Y(n_377) );
AND2x2_ASAP7_75t_L g389 ( .A(n_226), .B(n_266), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_226), .B(n_321), .Y(n_393) );
AND2x2_ASAP7_75t_L g430 ( .A(n_226), .B(n_425), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_226), .B(n_304), .Y(n_441) );
OR2x2_ASAP7_75t_L g443 ( .A(n_226), .B(n_379), .Y(n_443) );
INVx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g329 ( .A(n_227), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_227), .B(n_284), .Y(n_339) );
AND2x2_ASAP7_75t_L g351 ( .A(n_227), .B(n_266), .Y(n_351) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_227), .Y(n_381) );
AND2x4_ASAP7_75t_L g415 ( .A(n_227), .B(n_265), .Y(n_415) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_238), .Y(n_227) );
AOI21xp5_ASAP7_75t_SL g228 ( .A1(n_229), .A2(n_231), .B(n_236), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_237), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_240), .A2(n_476), .B(n_483), .Y(n_475) );
BUFx2_ASAP7_75t_L g263 ( .A(n_241), .Y(n_263) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g304 ( .A(n_242), .Y(n_304) );
AND2x2_ASAP7_75t_L g337 ( .A(n_242), .B(n_266), .Y(n_337) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g284 ( .A(n_243), .B(n_266), .Y(n_284) );
BUFx2_ASAP7_75t_L g330 ( .A(n_243), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g524 ( .A(n_250), .Y(n_524) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_256), .B(n_338), .Y(n_417) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_257), .B(n_280), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_257), .B(n_260), .Y(n_319) );
AND2x2_ASAP7_75t_L g374 ( .A(n_257), .B(n_310), .Y(n_374) );
AOI221xp5_ASAP7_75t_SL g311 ( .A1(n_258), .A2(n_312), .B1(n_320), .B2(n_322), .C(n_326), .Y(n_311) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g306 ( .A(n_259), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g347 ( .A(n_259), .B(n_348), .Y(n_347) );
OAI321xp33_ASAP7_75t_L g354 ( .A1(n_259), .A2(n_313), .A3(n_355), .B1(n_357), .B2(n_358), .C(n_360), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_260), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_263), .B(n_415), .Y(n_433) );
AND2x2_ASAP7_75t_L g320 ( .A(n_264), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_264), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
AND2x2_ASAP7_75t_L g303 ( .A(n_265), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_265), .B(n_378), .Y(n_408) );
INVx1_ASAP7_75t_L g445 ( .A(n_265), .Y(n_445) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_274), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g482 ( .A(n_275), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_282), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_279), .A2(n_389), .B(n_438), .C(n_439), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_280), .B(n_318), .Y(n_384) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_284), .B(n_287), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_284), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_284), .B(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_300), .B2(n_305), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g301 ( .A(n_287), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g324 ( .A(n_287), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g336 ( .A(n_287), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_287), .B(n_330), .Y(n_372) );
OR2x2_ASAP7_75t_L g379 ( .A(n_287), .B(n_304), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_287), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g429 ( .A(n_287), .B(n_415), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B1(n_295), .B2(n_297), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g335 ( .A(n_290), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_293), .A2(n_308), .B1(n_376), .B2(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g423 ( .A(n_294), .Y(n_423) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_298), .A2(n_335), .B1(n_338), .B2(n_339), .C(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g313 ( .A(n_299), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_303), .B(n_369), .Y(n_401) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_304), .Y(n_325) );
NAND2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
AND2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_353), .Y(n_352) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g396 ( .A(n_317), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_346), .B1(n_349), .B2(n_352), .C(n_354), .Y(n_345) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_324), .B(n_381), .Y(n_380) );
AOI21xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_328), .B(n_331), .Y(n_326) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_331), .Y(n_428) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g370 ( .A(n_333), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g391 ( .A(n_336), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_336), .B(n_396), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_339), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND4xp25_ASAP7_75t_L g344 ( .A(n_345), .B(n_363), .C(n_382), .D(n_395), .Y(n_344) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g353 ( .A(n_348), .Y(n_353) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_362), .Y(n_386) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_367), .C(n_375), .Y(n_363) );
AOI211xp5_ASAP7_75t_L g434 ( .A1(n_365), .A2(n_407), .B(n_435), .C(n_442), .Y(n_434) );
INVx1_ASAP7_75t_SL g394 ( .A(n_366), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_372), .B2(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_378), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_378), .B(n_389), .Y(n_422) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g399 ( .A(n_389), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_394), .Y(n_390) );
INVxp33_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI322xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_402), .C1(n_404), .C2(n_407), .Y(n_395) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND3xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_427), .C(n_434), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_416), .B2(n_418), .C(n_420), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g426 ( .A(n_415), .Y(n_426) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_430), .B2(n_431), .C(n_432), .Y(n_427) );
NAND2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g454 ( .A(n_447), .Y(n_454) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_455), .B(n_457), .C(n_745), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_458), .Y(n_737) );
INVx1_ASAP7_75t_L g462 ( .A(n_459), .Y(n_462) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g739 ( .A(n_466), .Y(n_739) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g740 ( .A(n_468), .Y(n_740) );
OR2x2_ASAP7_75t_SL g468 ( .A(n_469), .B(n_689), .Y(n_468) );
NAND5xp2_ASAP7_75t_L g469 ( .A(n_470), .B(n_601), .C(n_639), .D(n_660), .E(n_677), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_573), .C(n_594), .Y(n_470) );
OAI221xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_515), .B1(n_539), .B2(n_560), .C(n_564), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_485), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_474), .B(n_562), .Y(n_581) );
OR2x2_ASAP7_75t_L g608 ( .A(n_474), .B(n_498), .Y(n_608) );
AND2x2_ASAP7_75t_L g622 ( .A(n_474), .B(n_498), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_474), .B(n_488), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_474), .B(n_638), .Y(n_674) );
AND2x2_ASAP7_75t_L g703 ( .A(n_474), .B(n_613), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_474), .B(n_585), .Y(n_720) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g600 ( .A(n_475), .B(n_497), .Y(n_600) );
BUFx3_ASAP7_75t_L g625 ( .A(n_475), .Y(n_625) );
AND2x2_ASAP7_75t_L g654 ( .A(n_475), .B(n_498), .Y(n_654) );
AND3x2_ASAP7_75t_L g667 ( .A(n_475), .B(n_668), .C(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g590 ( .A(n_485), .Y(n_590) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
AOI32xp33_ASAP7_75t_L g645 ( .A1(n_486), .A2(n_597), .A3(n_646), .B1(n_649), .B2(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g572 ( .A(n_487), .B(n_497), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_487), .B(n_600), .Y(n_643) );
AND2x2_ASAP7_75t_L g650 ( .A(n_487), .B(n_622), .Y(n_650) );
OR2x2_ASAP7_75t_L g656 ( .A(n_487), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_487), .B(n_611), .Y(n_681) );
OR2x2_ASAP7_75t_L g699 ( .A(n_487), .B(n_527), .Y(n_699) );
BUFx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g563 ( .A(n_488), .B(n_507), .Y(n_563) );
INVx2_ASAP7_75t_L g585 ( .A(n_488), .Y(n_585) );
OR2x2_ASAP7_75t_L g607 ( .A(n_488), .B(n_507), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_488), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_488), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g668 ( .A(n_488), .B(n_562), .Y(n_668) );
INVx1_ASAP7_75t_SL g719 ( .A(n_497), .Y(n_719) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx1_ASAP7_75t_SL g562 ( .A(n_498), .Y(n_562) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_498), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_498), .B(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_498), .B(n_585), .C(n_703), .Y(n_714) );
INVx2_ASAP7_75t_L g613 ( .A(n_507), .Y(n_613) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_507), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
INVx1_ASAP7_75t_L g649 ( .A(n_516), .Y(n_649) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g567 ( .A(n_517), .B(n_550), .Y(n_567) );
INVx2_ASAP7_75t_L g584 ( .A(n_517), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_517), .B(n_551), .Y(n_589) );
AND2x2_ASAP7_75t_L g604 ( .A(n_517), .B(n_540), .Y(n_604) );
AND2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_588), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_526), .B(n_632), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_526), .B(n_589), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_526), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_526), .B(n_583), .Y(n_711) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g549 ( .A(n_527), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_527), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_540), .Y(n_593) );
AND2x2_ASAP7_75t_L g619 ( .A(n_527), .B(n_550), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_527), .B(n_659), .Y(n_658) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_531), .B(n_538), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_529), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g578 ( .A(n_531), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_540), .B(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g583 ( .A(n_540), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_SL g588 ( .A(n_540), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_540), .B(n_575), .Y(n_641) );
OR2x2_ASAP7_75t_L g651 ( .A(n_540), .B(n_577), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_540), .B(n_619), .Y(n_679) );
OR2x2_ASAP7_75t_L g709 ( .A(n_540), .B(n_550), .Y(n_709) );
AND2x2_ASAP7_75t_L g713 ( .A(n_540), .B(n_551), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_540), .B(n_589), .Y(n_726) );
AND2x2_ASAP7_75t_L g733 ( .A(n_540), .B(n_615), .Y(n_733) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_547), .Y(n_540) );
INVx1_ASAP7_75t_SL g676 ( .A(n_549), .Y(n_676) );
AND2x2_ASAP7_75t_L g615 ( .A(n_550), .B(n_577), .Y(n_615) );
AND2x2_ASAP7_75t_L g629 ( .A(n_550), .B(n_584), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_550), .B(n_588), .Y(n_632) );
INVx1_ASAP7_75t_L g659 ( .A(n_550), .Y(n_659) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g571 ( .A(n_551), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_561), .A2(n_607), .B(n_731), .C(n_732), .Y(n_730) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g637 ( .A(n_562), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_563), .B(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_622), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_568), .B(n_572), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_566), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g592 ( .A(n_567), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_567), .B(n_588), .Y(n_633) );
AND2x2_ASAP7_75t_L g724 ( .A(n_567), .B(n_575), .Y(n_724) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g597 ( .A(n_571), .B(n_584), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_582), .Y(n_598) );
OAI322xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_581), .A3(n_582), .B1(n_585), .B2(n_586), .C1(n_590), .C2(n_591), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
AND2x2_ASAP7_75t_L g685 ( .A(n_575), .B(n_597), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_575), .B(n_649), .Y(n_731) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g628 ( .A(n_577), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g694 ( .A(n_581), .B(n_607), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_582), .B(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_583), .B(n_615), .Y(n_672) );
AND2x2_ASAP7_75t_L g618 ( .A(n_584), .B(n_588), .Y(n_618) );
AND2x2_ASAP7_75t_L g626 ( .A(n_585), .B(n_627), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_585), .A2(n_664), .B(n_724), .C(n_725), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_586), .A2(n_599), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_588), .B(n_615), .Y(n_655) );
AND2x2_ASAP7_75t_L g661 ( .A(n_588), .B(n_629), .Y(n_661) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_597), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_589), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g705 ( .A(n_589), .Y(n_705) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_593), .A2(n_621), .B1(n_623), .B2(n_628), .Y(n_620) );
OAI22xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_595), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_630) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_600), .A2(n_702), .B1(n_704), .B2(n_706), .C(n_710), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B(n_609), .C(n_630), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g671 ( .A(n_607), .B(n_624), .Y(n_671) );
INVx1_ASAP7_75t_L g722 ( .A(n_607), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_608), .A2(n_610), .B1(n_614), .B2(n_617), .C(n_620), .Y(n_609) );
INVx2_ASAP7_75t_SL g664 ( .A(n_608), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g729 ( .A(n_611), .Y(n_729) );
AND2x2_ASAP7_75t_L g653 ( .A(n_612), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g638 ( .A(n_613), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g700 ( .A(n_616), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_624), .B(n_726), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g669 ( .A(n_627), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_628), .A2(n_640), .B(n_642), .C(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g717 ( .A(n_631), .Y(n_717) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_635), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_L g648 ( .A(n_638), .Y(n_648) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_651), .B1(n_652), .B2(n_655), .C1(n_656), .C2(n_658), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g684 ( .A(n_648), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_651), .B(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_652), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g657 ( .A(n_654), .Y(n_657) );
AND2x2_ASAP7_75t_L g721 ( .A(n_654), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g687 ( .A(n_657), .B(n_684), .Y(n_687) );
INVx1_ASAP7_75t_L g716 ( .A(n_658), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_665), .C(n_670), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_664), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_667), .A2(n_695), .A3(n_700), .B1(n_716), .B2(n_717), .C1(n_718), .C2(n_721), .Y(n_715) );
AND2x2_ASAP7_75t_L g702 ( .A(n_668), .B(n_703), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_673), .B2(n_675), .Y(n_670) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND5xp2_ASAP7_75t_L g689 ( .A(n_690), .B(n_701), .C(n_715), .D(n_723), .E(n_727), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_695), .B(n_696), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp33_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_703), .A2(n_728), .B(n_729), .C(n_730), .Y(n_727) );
AOI31xp33_ASAP7_75t_L g710 ( .A1(n_705), .A2(n_711), .A3(n_712), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g728 ( .A(n_726), .Y(n_728) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g741 ( .A(n_735), .Y(n_741) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
endmodule