module fake_jpeg_31151_n_73 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_6),
.B(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_14),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_1),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

OR2x4_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_2),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_3),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_29),
.C(n_26),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_20),
.C(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_21),
.B1(n_10),
.B2(n_11),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_53),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_9),
.B1(n_19),
.B2(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_7),
.B1(n_13),
.B2(n_15),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_48),
.C(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_45),
.Y(n_59)
);

OA21x2_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_61),
.B(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_58),
.C(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_68),
.B1(n_64),
.B2(n_67),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_69),
.Y(n_73)
);


endmodule