module fake_jpeg_2028_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_42),
.B1(n_37),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_42),
.B1(n_34),
.B2(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_46),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_57),
.B1(n_62),
.B2(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_48),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_44),
.B1(n_39),
.B2(n_40),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_18),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_36),
.C(n_17),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_36),
.B(n_2),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_11),
.B(n_12),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_108),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_24),
.B1(n_32),
.B2(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_109),
.B1(n_13),
.B2(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_8),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_15),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_94),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_92),
.C(n_25),
.Y(n_114)
);

OAI322xp33_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_121),
.A3(n_122),
.B1(n_109),
.B2(n_117),
.C1(n_26),
.C2(n_27),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_13),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_100),
.B1(n_107),
.B2(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_126),
.B1(n_106),
.B2(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_114),
.Y(n_130)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_128),
.A3(n_123),
.B1(n_119),
.B2(n_115),
.C(n_97),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_130),
.C(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_16),
.C(n_20),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_23),
.Y(n_139)
);


endmodule