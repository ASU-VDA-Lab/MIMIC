module real_jpeg_6824_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_44),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_1),
.A2(n_44),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_44),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_40),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_3),
.A2(n_40),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_40),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_4),
.Y(n_97)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_5),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_6),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_6),
.A2(n_88),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_77),
.B1(n_88),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_25),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_6),
.A2(n_330),
.B(n_332),
.C(n_340),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_6),
.B(n_356),
.C(n_358),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_6),
.B(n_147),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_6),
.B(n_268),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_6),
.B(n_74),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_7),
.Y(n_251)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_9),
.Y(n_424)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_43),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_12),
.A2(n_117),
.B1(n_120),
.B2(n_227),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_12),
.A2(n_86),
.B1(n_227),
.B2(n_336),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_12),
.A2(n_227),
.B1(n_366),
.B2(n_370),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_13),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_423),
.B(n_425),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_194),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_193),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_19),
.B(n_148),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_137),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_130),
.B2(n_131),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_57),
.B1(n_58),
.B2(n_129),
.Y(n_22)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_23),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B(n_41),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_24),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_25),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_25),
.B(n_134),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_25),
.B(n_226),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_31),
.Y(n_249)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_35),
.Y(n_229)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_41),
.B(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_46),
.B(n_88),
.Y(n_136)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_48),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_48),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_48),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_53),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_90),
.B1(n_91),
.B2(n_128),
.Y(n_58)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_59),
.B(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_59),
.A2(n_128),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_59),
.B(n_237),
.C(n_240),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_82),
.B(n_83),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_60),
.A2(n_181),
.B(n_188),
.Y(n_180)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_61),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_61),
.B(n_84),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_61),
.B(n_346),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_65),
.Y(n_339)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_80),
.Y(n_74)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_70),
.Y(n_357)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_74),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_74),
.B(n_346),
.Y(n_360)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_75),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_76),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_76),
.Y(n_265)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_79),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_79),
.Y(n_358)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_82),
.B(n_83),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_82),
.A2(n_157),
.B(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_88),
.A2(n_333),
.B(n_336),
.Y(n_332)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_122),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_140),
.B(n_147),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_92),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_115),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_96),
.Y(n_331)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_108),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_119),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_122),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_124),
.B(n_139),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_124),
.A2(n_139),
.B(n_147),
.Y(n_300)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_131),
.C(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_131),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_132),
.B(n_225),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_133),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_145),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_139),
.B(n_243),
.Y(n_271)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_146),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_147),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_165),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_154),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_155),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_157),
.B(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_162),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_189),
.B(n_190),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_167),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_180),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_189),
.B1(n_190),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_168),
.A2(n_180),
.B1(n_189),
.B2(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_168),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_168),
.A2(n_189),
.B1(n_329),
.B2(n_405),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_175),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_169),
.B(n_177),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_169),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_170),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_171),
.Y(n_369)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_180),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_188),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_188),
.B(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_230),
.B(n_422),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_196),
.B(n_199),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.C(n_206),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_200),
.Y(n_315)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_206),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_221),
.C(n_223),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_207),
.A2(n_208),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_209),
.B(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_210),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_213),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_214),
.A2(n_258),
.B(n_266),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_215),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_221),
.B(n_223),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_222),
.B(n_242),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_414),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_304),
.C(n_319),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_292),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_279),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_235),
.B(n_279),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.C(n_269),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_236),
.B(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_245),
.A2(n_246),
.B1(n_269),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_257),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_247),
.B(n_257),
.Y(n_287)
);

AOI32xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.A3(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_276),
.B(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_268),
.Y(n_383)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_274),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_274),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_275),
.B(n_382),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_276),
.B(n_364),
.Y(n_392)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_279),
.B(n_293),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.CI(n_286),
.CON(n_279),
.SN(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_289),
.C(n_290),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_292),
.A2(n_417),
.B(n_418),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_305),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_313),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_306),
.B(n_313),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_310),
.CI(n_312),
.CON(n_317),
.SN(n_317)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_317),
.B(n_318),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g428 ( 
.A(n_317),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_347),
.B(n_413),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_324),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.C(n_342),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_328),
.A2(n_342),
.B1(n_343),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_407),
.B(n_412),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_397),
.B(n_406),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_376),
.B(n_396),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_361),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_361),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_359),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_353),
.B1(n_359),
.B2(n_379),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_371),
.Y(n_361)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_374),
.C(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_384),
.B(n_395),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_380),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_391),
.B(n_394),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_400),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_403),
.C(n_404),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_411),
.Y(n_412)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_416),
.B(n_419),
.C(n_420),
.D(n_421),
.Y(n_414)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx8_ASAP7_75t_L g426 ( 
.A(n_424),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);


endmodule