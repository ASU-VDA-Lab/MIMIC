module fake_jpeg_9457_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_R g67 ( 
.A(n_36),
.B(n_16),
.Y(n_67)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_51),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_21),
.B2(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_19),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_24),
.B1(n_21),
.B2(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_72),
.B(n_84),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_81),
.B(n_61),
.Y(n_103)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_46),
.B1(n_35),
.B2(n_39),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_36),
.B1(n_35),
.B2(n_57),
.Y(n_102)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_36),
.B1(n_44),
.B2(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_42),
.B(n_46),
.C(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_51),
.A2(n_21),
.B1(n_38),
.B2(n_26),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_26),
.B1(n_38),
.B2(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_57),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_114),
.B1(n_97),
.B2(n_82),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_126),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_70),
.B1(n_55),
.B2(n_63),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_38),
.B1(n_22),
.B2(n_34),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_68),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_54),
.B(n_58),
.C(n_33),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_78),
.B(n_81),
.C(n_23),
.D(n_18),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_45),
.C(n_44),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_128),
.C(n_20),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_89),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_79),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_99),
.C(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_16),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_78),
.B1(n_60),
.B2(n_44),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_152),
.B1(n_157),
.B2(n_110),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_133),
.B(n_135),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_139),
.B1(n_150),
.B2(n_102),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_29),
.B(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_62),
.B1(n_83),
.B2(n_74),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_29),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_145),
.B(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_114),
.B1(n_108),
.B2(n_126),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_90),
.B1(n_97),
.B2(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_98),
.B1(n_80),
.B2(n_75),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_122),
.C(n_117),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_18),
.B1(n_23),
.B2(n_31),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_119),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_115),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_111),
.B1(n_121),
.B2(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_164),
.B1(n_179),
.B2(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_103),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_185),
.C(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_191),
.B1(n_31),
.B2(n_23),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_1),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_126),
.B(n_102),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_188),
.B1(n_162),
.B2(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_123),
.B1(n_128),
.B2(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_192),
.B1(n_146),
.B2(n_136),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_132),
.B1(n_138),
.B2(n_131),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_135),
.B(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_123),
.C(n_128),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_140),
.A2(n_118),
.B1(n_111),
.B2(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_125),
.B1(n_119),
.B2(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_94),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_194),
.B(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_195),
.B(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_202),
.B1(n_193),
.B2(n_183),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_130),
.B(n_136),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_200),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_127),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_215),
.C(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_163),
.A2(n_124),
.B1(n_53),
.B2(n_50),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_206),
.B(n_173),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_53),
.B(n_50),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_209),
.B1(n_166),
.B2(n_174),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_94),
.B1(n_34),
.B2(n_22),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_34),
.B1(n_22),
.B2(n_31),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_32),
.B(n_34),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_32),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_227),
.B1(n_248),
.B2(n_209),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_191),
.B1(n_178),
.B2(n_171),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_175),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_235),
.C(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_196),
.A2(n_192),
.B1(n_175),
.B2(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_182),
.C(n_186),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_199),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_161),
.B(n_174),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_203),
.B(n_202),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_196),
.A2(n_161),
.B1(n_189),
.B2(n_4),
.Y(n_242)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_2),
.C(n_3),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_217),
.C(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_15),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_222),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_210),
.B1(n_208),
.B2(n_220),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_194),
.B(n_198),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_223),
.B(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_248),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_231),
.C(n_240),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_263),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_230),
.B(n_224),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_236),
.B(n_226),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_207),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_199),
.B1(n_211),
.B2(n_213),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_267),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_216),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_213),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_269),
.C(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_12),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_211),
.B1(n_212),
.B2(n_217),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_207),
.C(n_3),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_269),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_276),
.B(n_261),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_263),
.C(n_235),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_277),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_287),
.B(n_270),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_234),
.C(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_243),
.C(n_225),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_13),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_13),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_12),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_252),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_253),
.B1(n_251),
.B2(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_2),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_298),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_9),
.B(n_11),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_250),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_301),
.C(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_260),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_281),
.B(n_256),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_262),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_257),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_284),
.C(n_271),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_308),
.B(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_272),
.B(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_283),
.C(n_255),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_301),
.C(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_11),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_290),
.C(n_291),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_308),
.B(n_313),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_288),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_5),
.B(n_6),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_320),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_302),
.B(n_304),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_328),
.C(n_318),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_321),
.C(n_6),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_325),
.Y(n_334)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.C(n_282),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_7),
.Y(n_336)
);


endmodule