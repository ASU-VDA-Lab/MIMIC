module fake_jpeg_3216_n_180 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_25),
.Y(n_33)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_10),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_26),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_16),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_4),
.B(n_6),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_71),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_82),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_63),
.B1(n_59),
.B2(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_23),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_38),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_62),
.C(n_93),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_34),
.B(n_38),
.C(n_35),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_69),
.B(n_80),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_52),
.B1(n_24),
.B2(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_101),
.B1(n_77),
.B2(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_107),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_99),
.Y(n_114)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_44),
.B1(n_10),
.B2(n_11),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_108),
.B1(n_110),
.B2(n_98),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_83),
.B1(n_68),
.B2(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_72),
.B1(n_60),
.B2(n_69),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_90),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_116),
.B(n_123),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_72),
.B1(n_60),
.B2(n_57),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_127),
.B1(n_110),
.B2(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_62),
.Y(n_122)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_57),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_130),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_94),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_95),
.C(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_108),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_97),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_114),
.A3(n_129),
.B1(n_126),
.B2(n_99),
.C1(n_107),
.C2(n_124),
.Y(n_150)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_98),
.B(n_112),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_107),
.B(n_102),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_122),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_130),
.B1(n_116),
.B2(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_151),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_135),
.B1(n_145),
.B2(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_141),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_138),
.C(n_132),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.C(n_163),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_154),
.B1(n_152),
.B2(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_132),
.C(n_134),
.Y(n_159)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_162),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_140),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_162),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_154),
.C(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.C(n_163),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_158),
.B1(n_160),
.B2(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_171),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_144),
.B1(n_161),
.B2(n_165),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_165),
.B(n_171),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_170),
.C(n_173),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_169),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);


endmodule