module real_jpeg_16848_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_2),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_4),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_6),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

AND2x4_ASAP7_75t_SL g71 ( 
.A(n_6),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_6),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_6),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_6),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_7),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_7),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_7),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_7),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_7),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_55),
.Y(n_54)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_10),
.B(n_64),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_10),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_10),
.B(n_36),
.Y(n_112)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_12),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_12),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_12),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_12),
.B(n_254),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_13),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_300),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_268),
.B(n_298),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_225),
.B(n_262),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_188),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_152),
.B(n_187),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_121),
.B(n_151),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_93),
.B(n_120),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_58),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_26),
.B(n_58),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_43),
.C(n_51),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_28),
.A2(n_41),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_103),
.B(n_112),
.C(n_141),
.Y(n_159)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_32),
.A2(n_33),
.B1(n_127),
.B2(n_136),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_32),
.B(n_136),
.C(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_32),
.B(n_141),
.C(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_37),
.C(n_41),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_33),
.B(n_292),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_34),
.B(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_37),
.A2(n_38),
.B1(n_164),
.B2(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_38),
.B(n_200),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_38),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_38),
.B(n_80),
.C(n_164),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_43),
.A2(n_51),
.B1(n_52),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_43),
.A2(n_44),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_47),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_47),
.A2(n_48),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_48),
.B(n_212),
.C(n_216),
.Y(n_234)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_53),
.A2(n_54),
.B1(n_99),
.B2(n_101),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_63),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_54),
.B(n_99),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_54),
.A2(n_99),
.B(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_54),
.B(n_62),
.C(n_132),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_55),
.Y(n_180)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_77),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_78),
.C(n_92),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_70),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_109),
.B(n_113),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_71),
.B(n_76),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_62),
.A2(n_63),
.B1(n_111),
.B2(n_112),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_96),
.B(n_98),
.C(n_103),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_75),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_73),
.A2(n_76),
.B1(n_131),
.B2(n_132),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_127),
.C(n_132),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_91),
.B2(n_92),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_90),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_84),
.C(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_80),
.A2(n_90),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_84),
.A2(n_236),
.B1(n_237),
.B2(n_241),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_84),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_84),
.B(n_234),
.C(n_237),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_84),
.B(n_211),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_84),
.A2(n_174),
.B1(n_175),
.B2(n_236),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_148),
.B1(n_163),
.B2(n_169),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_90),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_107),
.B(n_119),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_96),
.B(n_111),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_96),
.B(n_112),
.C(n_175),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_96),
.A2(n_117),
.B1(n_199),
.B2(n_205),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_96),
.B(n_201),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_99),
.A2(n_101),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_99),
.B(n_148),
.C(n_164),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_115),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_114),
.B(n_118),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_112),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_117),
.B(n_200),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_137),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_137),
.C(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

OR2x6_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_131),
.A2(n_132),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_146),
.C(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g292 ( 
.A1(n_141),
.A2(n_143),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_170),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_157),
.C(n_170),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_162),
.C(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_161),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_186),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_178),
.C(n_186),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_181),
.B(n_185),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_181),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_181),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_190),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_208),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_209),
.C(n_224),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_206),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_197),
.C(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_224),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_222),
.C(n_223),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_211),
.B(n_236),
.C(n_279),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_261),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_261),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_227),
.B(n_229),
.C(n_246),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_245),
.B2(n_246),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_272),
.C(n_273),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_251),
.C(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_258),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_297),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_297),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_286),
.C(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_286),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_284),
.C(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_332),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_305),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_325),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_324),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule