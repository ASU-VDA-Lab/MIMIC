module real_jpeg_25899_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVxp67_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_0),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_0),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_0),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_33),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_0),
.B(n_52),
.Y(n_260)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_17),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_52),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_2),
.B(n_49),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_2),
.B(n_47),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_66),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_2),
.B(n_27),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_4),
.B(n_33),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_4),
.B(n_52),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_6),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_6),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_17),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_6),
.B(n_52),
.Y(n_315)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_49),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_8),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_33),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_47),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_66),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_27),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_9),
.B(n_52),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_9),
.B(n_33),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_49),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_47),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_66),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_27),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_9),
.B(n_70),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_11),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_33),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_52),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_49),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_11),
.B(n_47),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_11),
.B(n_66),
.Y(n_316)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_13),
.B(n_66),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_14),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_14),
.B(n_33),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_14),
.B(n_52),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_14),
.B(n_49),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_14),
.B(n_47),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_14),
.B(n_66),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_16),
.B(n_47),
.Y(n_128)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_17),
.Y(n_149)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_17),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_21),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_71),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_22),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_23),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_60),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_30),
.B(n_84),
.C(n_94),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_30),
.A2(n_38),
.B1(n_83),
.B2(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_32),
.B(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_36),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_36),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_39),
.B(n_45),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_40),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_41),
.A2(n_42),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_44),
.B(n_165),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_45),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_52),
.Y(n_166)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_54),
.B(n_71),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_55),
.A2(n_56),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_57),
.B(n_62),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_59),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_61),
.B(n_63),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_74),
.C(n_76),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_65),
.A2(n_69),
.B1(n_75),
.B2(n_332),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_69),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_77),
.A2(n_78),
.B1(n_95),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_89),
.C(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_84),
.C(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_86),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_91),
.CI(n_92),
.CON(n_100),
.SN(n_100)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_95),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_102),
.C(n_105),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_97),
.B(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_99),
.B(n_100),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_100),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.C(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_118),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.CI(n_121),
.CON(n_118),
.SN(n_118)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_343),
.C(n_344),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_335),
.C(n_336),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_319),
.C(n_320),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_296),
.C(n_297),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_263),
.C(n_264),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_233),
.C(n_234),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_211),
.C(n_212),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_193),
.C(n_194),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_171),
.C(n_172),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_157),
.C(n_162),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_155),
.C(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_147),
.Y(n_152)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_152),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.C(n_167),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_184),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_177),
.C(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_183),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_192),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_197),
.C(n_202),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_205),
.C(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_210),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_228),
.C(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_222),
.C(n_223),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_216),
.Y(n_221)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_221),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_223),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.CI(n_226),
.CON(n_223),
.SN(n_223)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_225),
.C(n_226),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.CI(n_231),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_238),
.C(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_240),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.CI(n_243),
.CON(n_240),
.SN(n_240)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_256),
.C(n_261),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_256),
.B1(n_261),
.B2(n_262),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_252),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_287),
.C(n_288),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_259),
.C(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_283),
.B2(n_295),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_284),
.C(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_269),
.C(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_315),
.C(n_316),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.CI(n_294),
.CON(n_289),
.SN(n_289)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_317),
.B2(n_318),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_309),
.C(n_317),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_323),
.C(n_334),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_334),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_329),
.C(n_330),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_340),
.C(n_342),
.Y(n_343)
);


endmodule