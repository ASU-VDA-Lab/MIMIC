module real_jpeg_12225_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_30),
.B1(n_37),
.B2(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_3),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_119),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_4),
.A2(n_55),
.B1(n_58),
.B2(n_119),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_30),
.B1(n_37),
.B2(n_119),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_5),
.A2(n_41),
.B1(n_55),
.B2(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_55),
.B1(n_58),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_168),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_7),
.A2(n_30),
.B1(n_37),
.B2(n_168),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_10),
.A2(n_55),
.B1(n_58),
.B2(n_65),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_30),
.B1(n_37),
.B2(n_65),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_55),
.B1(n_58),
.B2(n_63),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_12),
.A2(n_30),
.B1(n_37),
.B2(n_63),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_13),
.B(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_13),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_60),
.B(n_195),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_186),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_13),
.A2(n_43),
.B(n_46),
.C(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_13),
.B(n_78),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_13),
.B(n_34),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_13),
.B(n_51),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_13),
.A2(n_58),
.B(n_72),
.C(n_257),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_14),
.A2(n_55),
.B1(n_58),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_71),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_14),
.A2(n_30),
.B1(n_37),
.B2(n_71),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_15),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_55),
.B1(n_58),
.B2(n_155),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_155),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_15),
.A2(n_30),
.B1(n_37),
.B2(n_155),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_16),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_16),
.A2(n_36),
.B1(n_55),
.B2(n_58),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_16),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_325)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_321),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_308),
.B(n_320),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_133),
.B(n_305),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_120),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_95),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_23),
.B(n_95),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_81),
.C(n_93),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_52),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_26),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_28),
.B1(n_52),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_27),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_34),
.B(n_35),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_29),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_29),
.A2(n_34),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_29),
.A2(n_34),
.B1(n_175),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_29),
.A2(n_34),
.B1(n_146),
.B2(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_29),
.A2(n_34),
.B1(n_189),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_29),
.A2(n_34),
.B1(n_186),
.B2(n_242),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_29),
.A2(n_34),
.B1(n_235),
.B2(n_242),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_30),
.B(n_244),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_109),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_33),
.A2(n_144),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_37),
.A2(n_47),
.B(n_186),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_40),
.A2(n_44),
.B1(n_51),
.B2(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_43),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_42),
.A2(n_58),
.A3(n_74),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_43),
.B(n_75),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_49),
.B1(n_51),
.B2(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_51),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_44),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_44),
.A2(n_51),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_44),
.A2(n_51),
.B1(n_149),
.B2(n_180),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_44),
.A2(n_51),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_44),
.A2(n_51),
.B1(n_221),
.B2(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_48),
.A2(n_113),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_48),
.A2(n_150),
.B1(n_179),
.B2(n_259),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_53),
.A2(n_54),
.B1(n_84),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_53),
.A2(n_54),
.B1(n_118),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_53),
.A2(n_54),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_53),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_54),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_55),
.B(n_186),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_55),
.A2(n_57),
.A3(n_60),
.B1(n_196),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_56),
.B(n_58),
.Y(n_210)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_61),
.B(n_186),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_81),
.B1(n_93),
.B2(n_94),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_68),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_70),
.A2(n_76),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_72),
.A2(n_78),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_72),
.A2(n_78),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_72),
.A2(n_78),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_76),
.A2(n_91),
.B1(n_115),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_76),
.A2(n_115),
.B1(n_116),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_76),
.A2(n_115),
.B1(n_170),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_76),
.A2(n_167),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_83),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_87),
.C(n_89),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_83),
.B(n_123),
.C(n_126),
.Y(n_309)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_92),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_87),
.B(n_129),
.C(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.C(n_103),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.C(n_117),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_105),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_290)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_120),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_121),
.B(n_122),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_132),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_158),
.B(n_304),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_135),
.B(n_156),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_136),
.B(n_139),
.Y(n_302)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_140),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.C(n_153),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_141),
.A2(n_142),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_143),
.B(n_147),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_151),
.B(n_153),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_152),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_299),
.B(n_303),
.Y(n_158)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_286),
.B1(n_297),
.B2(n_298),
.C(n_330),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_270),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_213),
.B(n_269),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_190),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_163),
.B(n_190),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.C(n_181),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_164),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_172),
.C(n_174),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_173),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_173),
.A2(n_283),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_173),
.A2(n_283),
.B1(n_316),
.B2(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_177),
.A2(n_181),
.B1(n_182),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_177),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_204),
.B2(n_212),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_191),
.B(n_205),
.C(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_193),
.B(n_199),
.C(n_203),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_206),
.B(n_209),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_263),
.B(n_268),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_251),
.B(n_262),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_231),
.B(n_250),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_217),
.B(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.C(n_229),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_239),
.B(n_249),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_237),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_245),
.B(n_248),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_258),
.C(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_272),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_281),
.C(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);


endmodule