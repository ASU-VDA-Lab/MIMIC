module fake_aes_2665_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_25;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
AND2x2_ASAP7_75t_SL g23 ( .A(n_19), .B(n_13), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_15), .B1(n_11), .B2(n_16), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
AOI33xp33_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_22), .A3(n_20), .B1(n_18), .B2(n_21), .B3(n_0), .Y(n_27) );
OAI22xp5_ASAP7_75t_SL g28 ( .A1(n_23), .A2(n_21), .B1(n_2), .B2(n_1), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_24), .Y(n_29) );
INVx3_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
CKINVDCx16_ASAP7_75t_R g32 ( .A(n_31), .Y(n_32) );
NAND2xp5_ASAP7_75t_SL g33 ( .A(n_32), .B(n_30), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_30), .Y(n_34) );
OAI222xp33_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_30), .B1(n_28), .B2(n_25), .C1(n_2), .C2(n_26), .Y(n_35) );
NAND2x1p5_ASAP7_75t_L g36 ( .A(n_34), .B(n_30), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_30), .Y(n_37) );
AOI222xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_35), .B1(n_28), .B2(n_25), .C1(n_10), .C2(n_9), .Y(n_38) );
endmodule