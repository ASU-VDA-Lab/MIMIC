module fake_jpeg_20282_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_42),
.B(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_35),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_21),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_48),
.B1(n_20),
.B2(n_24),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_60),
.B1(n_21),
.B2(n_1),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_17),
.B1(n_29),
.B2(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_29),
.B1(n_17),
.B2(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_78),
.Y(n_112)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_92),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_77),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_30),
.B1(n_24),
.B2(n_34),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_84),
.A2(n_91),
.B1(n_98),
.B2(n_2),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_45),
.C(n_19),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_96),
.C(n_0),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_99),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_28),
.B1(n_41),
.B2(n_26),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_97),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_19),
.C(n_26),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_26),
.B1(n_28),
.B2(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_33),
.B1(n_11),
.B2(n_15),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_33),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_104),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_21),
.A3(n_36),
.B1(n_15),
.B2(n_14),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_15),
.B(n_14),
.C(n_13),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_0),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_116),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_135),
.B(n_81),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_131),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_14),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_122),
.B(n_12),
.C(n_7),
.D(n_8),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_13),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_132),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_12),
.B(n_11),
.C(n_4),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_76),
.B(n_92),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_97),
.B1(n_96),
.B2(n_66),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_11),
.C(n_12),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_72),
.B(n_3),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_4),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_136),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_143),
.B(n_149),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_156),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_78),
.B1(n_76),
.B2(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_148),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_159),
.B(n_164),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_151),
.B1(n_158),
.B2(n_111),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_137),
.B1(n_127),
.B2(n_111),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_99),
.B(n_95),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_153),
.B(n_121),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_95),
.B(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_90),
.B1(n_105),
.B2(n_106),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_68),
.B(n_7),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_69),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_85),
.B(n_82),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_69),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_110),
.C(n_135),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_168),
.C(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_135),
.C(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_111),
.B1(n_107),
.B2(n_131),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_189),
.B1(n_142),
.B2(n_145),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_129),
.C(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_146),
.B(n_145),
.Y(n_176)
);

INVx2_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_139),
.C(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_142),
.C(n_146),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_130),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_183),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_124),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_186),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_123),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_132),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_108),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_108),
.B1(n_66),
.B2(n_106),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_119),
.A3(n_136),
.B1(n_71),
.B2(n_126),
.C1(n_82),
.C2(n_8),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_119),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_147),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_82),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_82),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_158),
.B(n_152),
.C(n_153),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_179),
.B(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_181),
.B1(n_171),
.B2(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_183),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_215),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_143),
.C(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_167),
.C(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_162),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_157),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_166),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_177),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_239),
.B(n_218),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_204),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_204),
.C(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_189),
.B1(n_191),
.B2(n_175),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_201),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_186),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_224),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_191),
.B1(n_182),
.B2(n_170),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_240),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_149),
.B1(n_185),
.B2(n_172),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_205),
.B1(n_200),
.B2(n_198),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_192),
.B(n_149),
.C(n_147),
.D(n_162),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_161),
.B1(n_163),
.B2(n_136),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_202),
.B1(n_136),
.B2(n_8),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_210),
.B1(n_202),
.B2(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_252),
.B1(n_257),
.B2(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_253),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_220),
.Y(n_247)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_223),
.B(n_208),
.C(n_202),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_255),
.C(n_256),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_198),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_214),
.C(n_199),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_209),
.C(n_214),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_219),
.C(n_199),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_240),
.C(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_266),
.C(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_230),
.B1(n_200),
.B2(n_205),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_229),
.C(n_234),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_221),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_269),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_239),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_202),
.B1(n_234),
.B2(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_260),
.C(n_269),
.Y(n_281)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_246),
.C(n_244),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_278),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_245),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_261),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_258),
.B(n_265),
.C(n_268),
.D(n_263),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_271),
.C(n_265),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_247),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_257),
.B(n_274),
.Y(n_287)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.C(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_273),
.C(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_248),
.A3(n_272),
.B1(n_284),
.B2(n_280),
.C1(n_251),
.C2(n_259),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_260),
.C(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_296),
.B(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_279),
.Y(n_299)
);


endmodule