module fake_netlist_1_2372_n_50 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_50);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_50;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_46;
wire n_48;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_9), .Y(n_18) );
INVx6_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_14), .B(n_0), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_10), .B(n_13), .Y(n_22) );
INVx5_ASAP7_75t_L g23 ( .A(n_11), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_3), .B(n_0), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_1), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_18), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_19), .B(n_1), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_16), .B(n_2), .Y(n_28) );
NOR2x2_ASAP7_75t_L g29 ( .A(n_17), .B(n_2), .Y(n_29) );
AND2x4_ASAP7_75t_L g30 ( .A(n_26), .B(n_24), .Y(n_30) );
AND2x4_ASAP7_75t_L g31 ( .A(n_25), .B(n_24), .Y(n_31) );
NAND3xp33_ASAP7_75t_L g32 ( .A(n_28), .B(n_22), .C(n_20), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_27), .Y(n_33) );
O2A1O1Ixp33_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_22), .B(n_29), .C(n_21), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVxp67_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_32), .Y(n_39) );
OAI22xp5_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_36), .B1(n_29), .B2(n_19), .Y(n_40) );
OAI22xp5_ASAP7_75t_L g41 ( .A1(n_38), .A2(n_23), .B1(n_4), .B2(n_5), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_42), .Y(n_43) );
AND2x4_ASAP7_75t_L g44 ( .A(n_41), .B(n_23), .Y(n_44) );
NOR3xp33_ASAP7_75t_SL g45 ( .A(n_40), .B(n_3), .C(n_4), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_43), .Y(n_46) );
INVx1_ASAP7_75t_L g47 ( .A(n_44), .Y(n_47) );
NAND3xp33_ASAP7_75t_L g48 ( .A(n_45), .B(n_23), .C(n_5), .Y(n_48) );
OR2x2_ASAP7_75t_L g49 ( .A(n_46), .B(n_44), .Y(n_49) );
OA22x2_ASAP7_75t_L g50 ( .A1(n_49), .A2(n_47), .B1(n_48), .B2(n_6), .Y(n_50) );
endmodule