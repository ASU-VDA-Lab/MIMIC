module fake_jpeg_24105_n_260 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_13),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_30),
.A2(n_28),
.B(n_20),
.C(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_23),
.Y(n_51)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_16),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_27),
.B1(n_16),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_52),
.B1(n_58),
.B2(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_50),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_17),
.C(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_54),
.B1(n_44),
.B2(n_20),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_35),
.B1(n_25),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_79),
.B1(n_40),
.B2(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_26),
.B1(n_24),
.B2(n_17),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_47),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_26),
.B1(n_21),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_40),
.A2(n_28),
.B1(n_20),
.B2(n_22),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_29),
.B1(n_19),
.B2(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_54),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_86),
.B(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_63),
.B1(n_60),
.B2(n_70),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_45),
.B(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_52),
.C(n_53),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_93),
.B(n_100),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_18),
.B(n_22),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_74),
.A3(n_65),
.B1(n_61),
.B2(n_66),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_60),
.B1(n_70),
.B2(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_99),
.Y(n_107)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_47),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_73),
.B1(n_28),
.B2(n_18),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_118),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_81),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_123),
.B(n_126),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_70),
.B1(n_78),
.B2(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_80),
.B1(n_71),
.B2(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_46),
.B1(n_32),
.B2(n_31),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_46),
.C(n_29),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_46),
.B1(n_29),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_101),
.B1(n_85),
.B2(n_99),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_29),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_11),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_90),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_141),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_133),
.Y(n_156)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_120),
.B1(n_109),
.B2(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_143),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_81),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_92),
.B(n_100),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_106),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_87),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_93),
.B(n_125),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_110),
.B1(n_121),
.B2(n_124),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_157),
.B1(n_165),
.B2(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_138),
.B(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_161),
.B(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_120),
.B1(n_123),
.B2(n_101),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_155),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_126),
.B1(n_100),
.B2(n_92),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_89),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_126),
.B1(n_115),
.B2(n_103),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_111),
.C(n_118),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_129),
.C(n_136),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_97),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_93),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_129),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_180),
.C(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_184),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_84),
.B1(n_97),
.B2(n_139),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_141),
.C(n_131),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_141),
.C(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_132),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_155),
.B1(n_159),
.B2(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_82),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_154),
.C(n_160),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_189),
.C(n_158),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_81),
.C(n_144),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_83),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_198),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_186),
.C(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_204),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_165),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_202),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_203),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_161),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_164),
.C(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_175),
.C(n_166),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_206),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_213),
.C(n_217),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_186),
.C(n_185),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_139),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_178),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_205),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_219),
.C(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_175),
.C(n_173),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_199),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_173),
.B(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_230),
.B1(n_10),
.B2(n_9),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_173),
.C(n_152),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_229),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_11),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_211),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_140),
.B(n_133),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_133),
.B1(n_91),
.B2(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_207),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_91),
.B1(n_10),
.B2(n_9),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_231),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_91),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_240),
.B1(n_1),
.B2(n_4),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_234),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_244),
.B1(n_238),
.B2(n_240),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_224),
.B(n_5),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_247),
.B(n_5),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_4),
.B(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_249),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_246),
.B(n_6),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_5),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_252),
.A2(n_7),
.B(n_240),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_7),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_256),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_254),
.B(n_257),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_259),
.Y(n_260)
);


endmodule