module fake_jpeg_1245_n_651 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_651);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_651;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_19),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_59),
.B(n_110),
.C(n_55),
.Y(n_156)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_61),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_62),
.B(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_129),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_70),
.Y(n_160)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx8_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_72),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_100),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_1),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_93),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_1),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_33),
.B(n_2),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_43),
.C(n_41),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_2),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_33),
.B(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_106),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_2),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_39),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_24),
.B(n_3),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_114),
.Y(n_169)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_3),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_27),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_118),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_24),
.B(n_4),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_27),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_5),
.Y(n_204)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_39),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_134),
.B(n_140),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_136),
.B(n_156),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_62),
.B(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_39),
.B1(n_58),
.B2(n_36),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_141),
.A2(n_58),
.B1(n_29),
.B2(n_30),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_145),
.B(n_146),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_28),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_151),
.B(n_153),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_28),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_57),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_155),
.B(n_159),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_39),
.C(n_57),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_34),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_57),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_63),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_165),
.B(n_168),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_24),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_41),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_172),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_26),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_86),
.B(n_36),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_55),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_186),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_58),
.B1(n_34),
.B2(n_29),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_181),
.A2(n_148),
.B(n_160),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_77),
.B(n_43),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_42),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_74),
.B(n_42),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_76),
.B(n_45),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_49),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_205),
.Y(n_289)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_83),
.B(n_45),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_91),
.B(n_26),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_95),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_217),
.Y(n_293)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_124),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_224),
.Y(n_333)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

CKINVDCx12_ASAP7_75t_R g227 ( 
.A(n_180),
.Y(n_227)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_185),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_231),
.Y(n_326)
);

INVx6_ASAP7_75t_SL g232 ( 
.A(n_180),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_232),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_233),
.A2(n_245),
.B1(n_249),
.B2(n_261),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_234),
.B(n_248),
.C(n_272),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_56),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_277),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_149),
.A2(n_122),
.B1(n_119),
.B2(n_116),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_237),
.A2(n_143),
.B1(n_198),
.B2(n_210),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_238),
.B(n_150),
.C(n_212),
.Y(n_335)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_184),
.B(n_50),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_243),
.B(n_250),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_185),
.A2(n_34),
.B1(n_38),
.B2(n_30),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_142),
.A2(n_115),
.B1(n_111),
.B2(n_105),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_246),
.A2(n_270),
.B1(n_273),
.B2(n_287),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_131),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_130),
.A2(n_29),
.B1(n_38),
.B2(n_30),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_169),
.B(n_38),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_252),
.Y(n_355)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_258),
.Y(n_347)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_259),
.Y(n_343)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_260),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_130),
.A2(n_103),
.B1(n_53),
.B2(n_35),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_161),
.B(n_6),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_264),
.Y(n_307)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_137),
.B(n_6),
.Y(n_264)
);

BUFx16f_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_265),
.Y(n_303)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_195),
.Y(n_267)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_138),
.B(n_7),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_274),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_191),
.A2(n_35),
.B1(n_53),
.B2(n_9),
.Y(n_270)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_219),
.A2(n_35),
.B1(n_53),
.B2(n_10),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_139),
.B(n_7),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_174),
.B(n_8),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_278),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_183),
.B(n_8),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_133),
.B(n_10),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_164),
.Y(n_279)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_132),
.B(n_10),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_283),
.Y(n_344)
);

BUFx12_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_133),
.B(n_13),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_141),
.A2(n_156),
.B1(n_219),
.B2(n_143),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_192),
.B1(n_213),
.B2(n_210),
.Y(n_320)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_164),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_294),
.Y(n_332)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_191),
.A2(n_35),
.B1(n_53),
.B2(n_13),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_173),
.B(n_53),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_297),
.Y(n_325)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_158),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_295),
.B(n_171),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_181),
.B(n_53),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_299),
.Y(n_357)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

OA22x2_ASAP7_75t_SL g301 ( 
.A1(n_224),
.A2(n_189),
.B1(n_188),
.B2(n_167),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_301),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_148),
.B(n_192),
.C(n_175),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_304),
.A2(n_285),
.B(n_267),
.C(n_229),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_152),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_306),
.A2(n_314),
.B1(n_315),
.B2(n_342),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_177),
.B1(n_154),
.B2(n_201),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_276),
.A2(n_177),
.B1(n_154),
.B2(n_201),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_160),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_319),
.B(n_300),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_320),
.A2(n_330),
.B1(n_265),
.B2(n_232),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_235),
.A2(n_150),
.B(n_212),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_293),
.A2(n_147),
.B1(n_199),
.B2(n_200),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_335),
.B(n_300),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_237),
.A2(n_199),
.B1(n_200),
.B2(n_198),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_240),
.B1(n_226),
.B2(n_222),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_221),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_345),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_254),
.A2(n_171),
.B1(n_176),
.B2(n_213),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_224),
.B(n_221),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_224),
.B(n_194),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_348),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_242),
.B(n_194),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_353),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_230),
.B(n_176),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_291),
.Y(n_370)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_255),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_L g433 ( 
.A1(n_366),
.A2(n_371),
.B(n_373),
.Y(n_433)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_370),
.B(n_386),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_244),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_236),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_375),
.B1(n_385),
.B2(n_266),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_378),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_239),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_383),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_300),
.B1(n_294),
.B2(n_299),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_314),
.B1(n_315),
.B2(n_357),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_247),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_265),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_399),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_333),
.A2(n_225),
.B1(n_252),
.B2(n_293),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_313),
.B(n_259),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_260),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_391),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_388),
.A2(n_285),
.B(n_312),
.Y(n_442)
);

INVx2_ASAP7_75t_R g389 ( 
.A(n_304),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_389),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_296),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_345),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_394),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_308),
.B(n_253),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_397),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_308),
.B(n_289),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_307),
.B(n_251),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_401),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_359),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_279),
.B1(n_257),
.B2(n_258),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_402),
.A2(n_309),
.B(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_403),
.A2(n_355),
.B1(n_332),
.B2(n_256),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_303),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_405),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_332),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_325),
.B(n_292),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_302),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_305),
.B(n_288),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_340),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_335),
.C(n_305),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_425),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_306),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_413),
.A2(n_423),
.B1(n_428),
.B2(n_444),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_424),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_328),
.B1(n_323),
.B2(n_326),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_402),
.B1(n_382),
.B2(n_394),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_326),
.B1(n_301),
.B2(n_302),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_352),
.C(n_331),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_321),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_426),
.B(n_322),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_427),
.A2(n_429),
.B(n_405),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_367),
.A2(n_301),
.B1(n_331),
.B2(n_355),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_398),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_368),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_343),
.C(n_358),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_403),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_389),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_379),
.A2(n_390),
.B1(n_382),
.B2(n_396),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_378),
.B(n_317),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_446),
.B(n_407),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_371),
.Y(n_447)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_377),
.Y(n_450)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_476),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_452),
.A2(n_465),
.B1(n_468),
.B2(n_437),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_373),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_455),
.B(n_461),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_416),
.B(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_383),
.Y(n_458)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_408),
.Y(n_460)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_460),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_372),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_439),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_464),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_397),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_422),
.A2(n_379),
.B1(n_394),
.B2(n_389),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_388),
.B(n_384),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_467),
.A2(n_472),
.B(n_478),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_444),
.A2(n_381),
.B1(n_374),
.B2(n_361),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_439),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_471),
.Y(n_498)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_429),
.A2(n_361),
.B(n_388),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_482),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_416),
.B(n_434),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_477),
.Y(n_503)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_415),
.A2(n_362),
.B(n_312),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_414),
.B(n_401),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_481),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_363),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_411),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_437),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_L g546 ( 
.A1(n_485),
.A2(n_470),
.B(n_477),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_453),
.B1(n_468),
.B2(n_454),
.Y(n_523)
);

AOI32xp33_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_432),
.A3(n_446),
.B1(n_421),
.B2(n_391),
.Y(n_488)
);

AOI21xp33_ASAP7_75t_L g525 ( 
.A1(n_488),
.A2(n_464),
.B(n_456),
.Y(n_525)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_454),
.A2(n_419),
.B1(n_413),
.B2(n_441),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_492),
.A2(n_494),
.B1(n_453),
.B2(n_452),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_421),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_496),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_457),
.A2(n_436),
.B1(n_441),
.B2(n_420),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_409),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_387),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_497),
.B(n_499),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_445),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_425),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_500),
.B(n_509),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_420),
.C(n_436),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_501),
.B(n_504),
.C(n_516),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_443),
.C(n_365),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_447),
.B(n_443),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_369),
.Y(n_512)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_448),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_513),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_451),
.B(n_393),
.C(n_329),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_486),
.A2(n_457),
.B1(n_462),
.B2(n_469),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_519),
.A2(n_523),
.B1(n_494),
.B2(n_506),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_520),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_474),
.Y(n_522)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_528),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_495),
.B(n_465),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_526),
.B(n_485),
.Y(n_562)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_527),
.Y(n_572)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_484),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_529),
.B(n_530),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_504),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_532),
.Y(n_555)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_483),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_537),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_534),
.A2(n_535),
.B1(n_506),
.B2(n_470),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_492),
.A2(n_459),
.B1(n_467),
.B2(n_478),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_511),
.A2(n_489),
.B1(n_515),
.B2(n_507),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_496),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_499),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_SL g539 ( 
.A(n_491),
.B(n_490),
.C(n_508),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_542),
.C(n_545),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_490),
.B(n_472),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_502),
.Y(n_560)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_495),
.B(n_463),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_473),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_508),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_546),
.A2(n_438),
.B(n_431),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_516),
.C(n_510),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_549),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_510),
.C(n_491),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_502),
.C(n_485),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_550),
.B(n_563),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_556),
.B(n_560),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_561),
.A2(n_567),
.B1(n_534),
.B2(n_535),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_565),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_536),
.B(n_530),
.C(n_526),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_564),
.A2(n_546),
.B1(n_522),
.B2(n_539),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_543),
.B(n_514),
.C(n_362),
.Y(n_566)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_566),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_519),
.A2(n_482),
.B1(n_471),
.B2(n_460),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_536),
.B(n_438),
.C(n_431),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_571),
.C(n_541),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_540),
.Y(n_569)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_569),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_570),
.A2(n_412),
.B(n_364),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_317),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_551),
.A2(n_547),
.B(n_518),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_580),
.B1(n_584),
.B2(n_570),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_552),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_576),
.B(n_579),
.Y(n_608)
);

BUFx12_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_577),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_578),
.A2(n_582),
.B1(n_449),
.B2(n_339),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_568),
.B(n_520),
.C(n_531),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_561),
.A2(n_517),
.B1(n_449),
.B2(n_466),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_557),
.B(n_400),
.C(n_412),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_591),
.C(n_548),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_558),
.A2(n_554),
.B1(n_572),
.B2(n_567),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_586),
.A2(n_334),
.B(n_340),
.Y(n_609)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_559),
.Y(n_588)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_588),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_563),
.B(n_392),
.C(n_350),
.Y(n_591)
);

BUFx24_ASAP7_75t_SL g592 ( 
.A(n_555),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_592),
.B(n_585),
.Y(n_600)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_593),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_591),
.B(n_549),
.C(n_550),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_596),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_598),
.B1(n_599),
.B2(n_607),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_571),
.C(n_564),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_556),
.C(n_565),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_597),
.B(n_590),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_575),
.B(n_562),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_589),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_580),
.A2(n_310),
.B1(n_360),
.B2(n_329),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_603),
.A2(n_295),
.B1(n_175),
.B2(n_268),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_350),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_286),
.Y(n_620)
);

FAx1_ASAP7_75t_SL g606 ( 
.A(n_590),
.B(n_349),
.CI(n_347),
.CON(n_606),
.SN(n_606)
);

XNOR2x2_ASAP7_75t_SL g621 ( 
.A(n_606),
.B(n_282),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_586),
.A2(n_334),
.B(n_322),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_609),
.A2(n_573),
.B1(n_316),
.B2(n_310),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_612),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_582),
.C(n_583),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_617),
.Y(n_630)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_616),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_593),
.B(n_573),
.C(n_577),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_601),
.B(n_577),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_618),
.B(n_619),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_608),
.B(n_316),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_605),
.C(n_607),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g631 ( 
.A(n_621),
.B(n_623),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_SL g622 ( 
.A(n_598),
.B(n_223),
.C(n_282),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_609),
.Y(n_632)
);

AOI31xp67_ASAP7_75t_L g624 ( 
.A1(n_617),
.A2(n_597),
.A3(n_596),
.B(n_594),
.Y(n_624)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_624),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_614),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_625),
.A2(n_627),
.B1(n_612),
.B2(n_620),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_610),
.A2(n_599),
.B1(n_603),
.B2(n_604),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_632),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_630),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_635),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_615),
.C(n_622),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_SL g641 ( 
.A(n_636),
.B(n_631),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_629),
.A2(n_633),
.B1(n_631),
.B2(n_624),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_637),
.B(n_640),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_606),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_641),
.B(n_643),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_638),
.Y(n_643)
);

AOI322xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_634),
.A3(n_639),
.B1(n_640),
.B2(n_631),
.C1(n_621),
.C2(n_606),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_SL g647 ( 
.A1(n_645),
.A2(n_642),
.B(n_223),
.C(n_280),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_646),
.C(n_223),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_228),
.B1(n_271),
.B2(n_206),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_223),
.B1(n_263),
.B2(n_218),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_218),
.Y(n_651)
);


endmodule