module fake_jpeg_16710_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_9),
.B(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_68),
.B(n_87),
.Y(n_171)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_29),
.B1(n_23),
.B2(n_37),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_110),
.Y(n_131)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_14),
.B1(n_21),
.B2(n_20),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_15),
.C(n_25),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_88),
.C(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_38),
.B(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_15),
.C(n_25),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_10),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_16),
.B1(n_28),
.B2(n_21),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_93),
.A2(n_97),
.B1(n_108),
.B2(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_41),
.A2(n_16),
.B1(n_30),
.B2(n_19),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_96),
.A2(n_93),
.B1(n_112),
.B2(n_108),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_66),
.B1(n_63),
.B2(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_45),
.B(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_2),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_40),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_52),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_40),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_12),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_11),
.Y(n_122)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_61),
.A2(n_36),
.B1(n_34),
.B2(n_15),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_160),
.Y(n_172)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_137),
.Y(n_174)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_73),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_133),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_135),
.B(n_141),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_34),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_143),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_155),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_78),
.A2(n_11),
.B(n_27),
.C(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_64),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_78),
.B(n_2),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_71),
.B(n_2),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_167),
.B1(n_163),
.B2(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_79),
.B(n_111),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_69),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_80),
.B1(n_75),
.B2(n_91),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_3),
.C(n_7),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_8),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_88),
.B(n_3),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_10),
.Y(n_196)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_184),
.A2(n_188),
.B(n_192),
.Y(n_236)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_210),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_9),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_72),
.B(n_116),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_72),
.B(n_102),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_198),
.B1(n_205),
.B2(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_190),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_75),
.B1(n_91),
.B2(n_99),
.Y(n_198)
);

BUFx24_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_113),
.B(n_77),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_203),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_124),
.A2(n_117),
.B1(n_100),
.B2(n_92),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_100),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_203),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_130),
.A2(n_113),
.B1(n_152),
.B2(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_214),
.B1(n_217),
.B2(n_144),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_134),
.B1(n_168),
.B2(n_125),
.Y(n_222)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_182),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_147),
.A2(n_149),
.B1(n_166),
.B2(n_150),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_140),
.B1(n_131),
.B2(n_134),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_164),
.B(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_139),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_140),
.A2(n_123),
.B1(n_161),
.B2(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_219),
.B(n_221),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_224),
.B1(n_232),
.B2(n_253),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_222),
.B(n_237),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_225),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_129),
.B1(n_138),
.B2(n_127),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_175),
.B(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_136),
.C(n_207),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_172),
.B(n_136),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_240),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_238),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_213),
.B1(n_175),
.B2(n_209),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_244),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_180),
.B(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_188),
.B(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_258),
.C(n_200),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_176),
.B(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_187),
.A2(n_201),
.B1(n_204),
.B2(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_239),
.B1(n_218),
.B2(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_184),
.B(n_176),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_200),
.B(n_181),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_204),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_202),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_202),
.B(n_195),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_195),
.B(n_185),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_262),
.B(n_280),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_260),
.B(n_276),
.Y(n_311)
);

AO22x2_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_181),
.B1(n_197),
.B2(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_281),
.B1(n_289),
.B2(n_262),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_235),
.B(n_226),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_265),
.B(n_277),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_220),
.B1(n_222),
.B2(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_271),
.B(n_284),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_281),
.B1(n_282),
.B2(n_289),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_236),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_283),
.C(n_290),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_232),
.B(n_246),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_219),
.A3(n_224),
.B1(n_243),
.B2(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_253),
.B(n_258),
.Y(n_280)
);

AO21x2_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_223),
.B(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_233),
.A2(n_244),
.B1(n_239),
.B2(n_242),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_231),
.A2(n_218),
.B1(n_229),
.B2(n_241),
.Y(n_284)
);

AOI22x1_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_229),
.B1(n_234),
.B2(n_238),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_247),
.C(n_234),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_251),
.A2(n_235),
.B(n_232),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_273),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_263),
.B1(n_280),
.B2(n_318),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_272),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_303),
.B(n_304),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_283),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_279),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_306),
.A2(n_310),
.B1(n_313),
.B2(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_279),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_268),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_263),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_274),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_276),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_263),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_287),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_322),
.C(n_330),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_275),
.C(n_265),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_317),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_338),
.C(n_340),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_300),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_331),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_293),
.B1(n_302),
.B2(n_316),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_337),
.A2(n_307),
.B1(n_309),
.B2(n_314),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_317),
.C(n_316),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_293),
.C(n_298),
.Y(n_340)
);

XOR2x2_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_311),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_297),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_315),
.C(n_301),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_330),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_346),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_347),
.A2(n_351),
.B1(n_358),
.B2(n_343),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_350),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_339),
.B(n_340),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_294),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_360),
.C(n_322),
.Y(n_365)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_336),
.Y(n_359)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_338),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_368),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_372),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_347),
.A2(n_335),
.B(n_342),
.Y(n_364)
);

AOI21xp33_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_349),
.B(n_357),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_369),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_328),
.C(n_337),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_328),
.C(n_341),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_296),
.B1(n_303),
.B2(n_348),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_357),
.B1(n_368),
.B2(n_363),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_360),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_374),
.A2(n_370),
.B1(n_367),
.B2(n_369),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_380),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_378),
.B(n_379),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_364),
.A2(n_371),
.B1(n_362),
.B2(n_361),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_379),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_367),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_373),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_385),
.B(n_387),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_366),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_373),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_385),
.C(n_382),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_388),
.B(n_380),
.Y(n_391)
);

AO21x1_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_375),
.B(n_382),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_378),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_375),
.C(n_365),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_376),
.Y(n_395)
);


endmodule