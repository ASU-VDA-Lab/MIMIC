module fake_jpeg_29240_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_36),
.B1(n_29),
.B2(n_16),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_67),
.B1(n_60),
.B2(n_57),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_39),
.C(n_19),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_61),
.C(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_47),
.B1(n_52),
.B2(n_42),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_62),
.B(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_6),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_4),
.B(n_5),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_6),
.B(n_7),
.Y(n_68)
);

NAND5xp2_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_10),
.C(n_12),
.D(n_13),
.E(n_14),
.Y(n_78)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_8),
.B(n_9),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_78),
.B1(n_69),
.B2(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_73),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_76),
.B(n_71),
.C(n_69),
.D(n_70),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_15),
.B(n_17),
.C(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_22),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_27),
.B(n_24),
.C(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_23),
.Y(n_86)
);


endmodule