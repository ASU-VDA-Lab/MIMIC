module fake_netlist_1_12404_n_49 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_49);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_49;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_48;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
AND2x4_ASAP7_75t_L g17 ( .A(n_15), .B(n_13), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_10), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_1), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_1), .B(n_2), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_8), .B(n_2), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_4), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_20), .Y(n_27) );
AND2x6_ASAP7_75t_SL g28 ( .A(n_22), .B(n_0), .Y(n_28) );
OAI21xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_17), .B(n_23), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_25), .B(n_17), .Y(n_30) );
INVxp67_ASAP7_75t_SL g31 ( .A(n_30), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_25), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_26), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI31xp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_32), .A3(n_23), .B(n_28), .Y(n_36) );
OAI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_32), .B1(n_18), .B2(n_26), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_37), .B(n_24), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g40 ( .A(n_36), .B(n_24), .Y(n_40) );
BUFx2_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
NOR2x1_ASAP7_75t_L g42 ( .A(n_40), .B(n_24), .Y(n_42) );
OAI22xp5_ASAP7_75t_L g43 ( .A1(n_39), .A2(n_21), .B1(n_4), .B2(n_3), .Y(n_43) );
OAI22xp5_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_21), .B1(n_3), .B2(n_6), .Y(n_44) );
HB1xp67_ASAP7_75t_L g45 ( .A(n_41), .Y(n_45) );
NOR3xp33_ASAP7_75t_L g46 ( .A(n_43), .B(n_21), .C(n_7), .Y(n_46) );
XNOR2xp5_ASAP7_75t_L g47 ( .A(n_45), .B(n_5), .Y(n_47) );
OAI22xp5_ASAP7_75t_L g48 ( .A1(n_44), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_48) );
AOI22xp33_ASAP7_75t_L g49 ( .A1(n_48), .A2(n_16), .B1(n_46), .B2(n_47), .Y(n_49) );
endmodule