module fake_netlist_5_1050_n_1593 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1593);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1593;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_72),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_41),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_87),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_52),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_57),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_53),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_28),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_115),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_65),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_30),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_38),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_35),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_30),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_20),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_25),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_7),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_83),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_49),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_39),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_37),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_41),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_135),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_22),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_21),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_81),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_21),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_47),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_74),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_26),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_11),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_59),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_78),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_43),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_46),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_36),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_2),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_3),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_40),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_34),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_103),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_45),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_138),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_50),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_45),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_71),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_35),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_102),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_54),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_123),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_114),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_10),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_15),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_29),
.Y(n_277)
);

BUFx8_ASAP7_75t_SL g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_38),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_12),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_18),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_104),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_122),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_16),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_8),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_56),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_60),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_131),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_145),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_113),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_97),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_120),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_95),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_93),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_86),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_43),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_174),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_187),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_191),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_187),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_187),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_187),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_187),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_234),
.B(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_158),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_161),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_177),
.B(n_4),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_171),
.B(n_5),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_165),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_173),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_276),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_191),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_179),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_181),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_198),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_184),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_188),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_189),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_234),
.B(n_5),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_168),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_192),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_294),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_294),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_168),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_299),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_194),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_204),
.B(n_234),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_174),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_155),
.B(n_10),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_170),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_170),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_160),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_258),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_258),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_172),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_199),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_200),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_202),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_176),
.B(n_11),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_207),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_182),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_304),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_315),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_316),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_320),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_152),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_321),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_152),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_303),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_305),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_326),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_311),
.B(n_243),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_331),
.B(n_293),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_306),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_166),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_172),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_166),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_231),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_307),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_359),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_329),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_334),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_335),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_323),
.B(n_178),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_340),
.B(n_231),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_307),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_308),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_309),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_309),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_344),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_351),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_325),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_367),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_331),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_332),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_R g434 ( 
.A(n_312),
.B(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_369),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_374),
.B(n_371),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_433),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_431),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_375),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_374),
.B(n_337),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_405),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_395),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_403),
.B(n_155),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_185),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_394),
.A2(n_319),
.B1(n_354),
.B2(n_370),
.Y(n_453)
);

BUFx8_ASAP7_75t_SL g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_405),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_417),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_417),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_386),
.B(n_348),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_401),
.B(n_417),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_337),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_403),
.B(n_197),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_411),
.A2(n_245),
.B1(n_255),
.B2(n_153),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_302),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_408),
.B(n_414),
.Y(n_468)
);

NOR2x1p5_ASAP7_75t_L g469 ( 
.A(n_372),
.B(n_156),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_348),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_339),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_185),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_411),
.A2(n_228),
.B1(n_284),
.B2(n_197),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_206),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_386),
.B(n_366),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_383),
.B(n_339),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_408),
.B(n_206),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_389),
.B(n_228),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_387),
.B(n_398),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_431),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_406),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_408),
.B(n_284),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_434),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_408),
.B(n_175),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_411),
.A2(n_283),
.B1(n_251),
.B2(n_236),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_377),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_342),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_411),
.B(n_343),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_380),
.B(n_175),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_413),
.A2(n_167),
.B1(n_205),
.B2(n_208),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_381),
.B(n_353),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_384),
.B(n_355),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_393),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_407),
.B(n_355),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_391),
.B(n_175),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_164),
.C(n_157),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_409),
.B(n_341),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_410),
.B(n_221),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_392),
.B(n_226),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_413),
.B(n_186),
.C(n_183),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_404),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_420),
.B(n_361),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_415),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_396),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_424),
.B(n_361),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_428),
.B(n_201),
.C(n_190),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_362),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_373),
.B(n_169),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_415),
.B(n_175),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_373),
.B(n_362),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_376),
.B(n_196),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_423),
.B(n_226),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_379),
.B(n_363),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_379),
.B(n_364),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_382),
.B(n_175),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_382),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_435),
.A2(n_287),
.B1(n_219),
.B2(n_218),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_388),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_432),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_388),
.B(n_364),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_399),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_399),
.B(n_209),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_402),
.B(n_365),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_402),
.B(n_217),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_416),
.B(n_221),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_418),
.B(n_286),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_419),
.B(n_233),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_422),
.B(n_233),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_422),
.B(n_223),
.Y(n_562)
);

INVx6_ASAP7_75t_L g563 ( 
.A(n_432),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

AND2x6_ASAP7_75t_L g565 ( 
.A(n_427),
.B(n_223),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_300),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_432),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_425),
.A2(n_280),
.B1(n_268),
.B2(n_203),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_432),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_425),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_432),
.B(n_300),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_458),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_483),
.B(n_214),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_438),
.B(n_215),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_459),
.B(n_154),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_463),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

BUFx5_ASAP7_75t_L g582 ( 
.A(n_474),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_534),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_491),
.B(n_216),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_159),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_460),
.B(n_477),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_345),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_443),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_495),
.B(n_163),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_550),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_436),
.B(n_223),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_496),
.B(n_223),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_470),
.B(n_346),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_472),
.B(n_180),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_523),
.Y(n_597)
);

O2A1O1Ixp5_ASAP7_75t_L g598 ( 
.A1(n_451),
.A2(n_224),
.B(n_195),
.C(n_271),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_470),
.B(n_496),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_472),
.B(n_193),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_453),
.A2(n_213),
.B(n_235),
.C(n_222),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_472),
.B(n_210),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_457),
.B(n_473),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_473),
.B(n_220),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_451),
.A2(n_279),
.B1(n_257),
.B2(n_247),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_464),
.B(n_269),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_530),
.A2(n_270),
.B(n_298),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_500),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_464),
.A2(n_247),
.B1(n_257),
.B2(n_279),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_545),
.B(n_547),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_500),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_550),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_468),
.A2(n_347),
.B1(n_350),
.B2(n_349),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_559),
.B(n_211),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_445),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_570),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_453),
.A2(n_223),
.B1(n_261),
.B2(n_290),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_448),
.B(n_212),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_466),
.B(n_365),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_468),
.B(n_227),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_555),
.B(n_238),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_501),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_531),
.B(n_261),
.Y(n_625)
);

CKINVDCx11_ASAP7_75t_R g626 ( 
.A(n_484),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_449),
.B(n_225),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_493),
.A2(n_263),
.B(n_289),
.C(n_288),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_523),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_523),
.Y(n_630)
);

AOI22x1_ASAP7_75t_SL g631 ( 
.A1(n_484),
.A2(n_301),
.B1(n_241),
.B2(n_242),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_452),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_551),
.B(n_261),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_455),
.B(n_229),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_456),
.B(n_232),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_549),
.B(n_230),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_246),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_538),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_474),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_493),
.A2(n_261),
.B1(n_290),
.B2(n_230),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_445),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_488),
.A2(n_295),
.B1(n_293),
.B2(n_230),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_461),
.B(n_237),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_480),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_248),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_570),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_462),
.B(n_239),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_542),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_474),
.A2(n_290),
.B1(n_261),
.B2(n_262),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_465),
.B(n_252),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_479),
.A2(n_297),
.B1(n_296),
.B2(n_244),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_475),
.B(n_240),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_488),
.B(n_266),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_506),
.B(n_267),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_474),
.A2(n_290),
.B1(n_259),
.B2(n_264),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_479),
.A2(n_272),
.B1(n_292),
.B2(n_250),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_506),
.B(n_249),
.Y(n_659)
);

NOR2x1p5_ASAP7_75t_L g660 ( 
.A(n_494),
.B(n_273),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_492),
.B(n_290),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_532),
.B(n_265),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_488),
.B(n_274),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_474),
.A2(n_295),
.B1(n_282),
.B2(n_275),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_492),
.B(n_256),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_442),
.Y(n_667)
);

AO221x1_ASAP7_75t_L g668 ( 
.A1(n_499),
.A2(n_295),
.B1(n_14),
.B2(n_16),
.C(n_18),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_254),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_452),
.B(n_253),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_452),
.B(n_573),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_553),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_573),
.B(n_61),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_535),
.B(n_55),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_515),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_571),
.B(n_69),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_498),
.B(n_533),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_490),
.B(n_147),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_535),
.B(n_144),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_557),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_466),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_505),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_539),
.B(n_132),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_129),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_558),
.B(n_118),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_557),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_558),
.B(n_112),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_454),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_490),
.B(n_110),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_560),
.B(n_107),
.Y(n_690)
);

AND2x6_ASAP7_75t_SL g691 ( 
.A(n_466),
.B(n_13),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_560),
.B(n_101),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_520),
.B(n_14),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_481),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_19),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_561),
.B(n_96),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_498),
.B(n_19),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_561),
.B(n_92),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_520),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_471),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_482),
.B(n_89),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_482),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_481),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_82),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_566),
.B(n_77),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_552),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_566),
.B(n_75),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_503),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_554),
.B(n_70),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_525),
.B(n_23),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_503),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_509),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_509),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_450),
.B(n_46),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_440),
.B(n_24),
.C(n_26),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_450),
.B(n_29),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_514),
.B(n_521),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_514),
.B(n_31),
.Y(n_719)
);

O2A1O1Ixp5_ASAP7_75t_L g720 ( 
.A1(n_562),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_510),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_469),
.B(n_33),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_516),
.B(n_34),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_516),
.B(n_37),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_SL g725 ( 
.A(n_546),
.B(n_40),
.C(n_42),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_485),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_517),
.B(n_526),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_517),
.B(n_527),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_482),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_513),
.B(n_489),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_487),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_487),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_546),
.B(n_568),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_521),
.B(n_522),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_522),
.B(n_536),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_523),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_478),
.B(n_508),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_574),
.B(n_568),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_624),
.B(n_609),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_671),
.A2(n_603),
.B(n_587),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_667),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_727),
.A2(n_528),
.B(n_446),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_728),
.A2(n_441),
.B(n_446),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_585),
.B(n_562),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_612),
.B(n_556),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_630),
.A2(n_441),
.B(n_467),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_667),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_575),
.B(n_556),
.Y(n_748)
);

AO32x1_ASAP7_75t_L g749 ( 
.A1(n_686),
.A2(n_536),
.A3(n_510),
.B1(n_529),
.B2(n_486),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_630),
.A2(n_692),
.B(n_619),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_599),
.B(n_583),
.Y(n_751)
);

NOR2x1_ASAP7_75t_L g752 ( 
.A(n_730),
.B(n_519),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_618),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_623),
.B(n_504),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_588),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_619),
.A2(n_502),
.B(n_489),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_636),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_576),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_601),
.A2(n_537),
.B(n_544),
.C(n_572),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_467),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_608),
.A2(n_629),
.B(n_597),
.Y(n_762)
);

OR2x6_ASAP7_75t_SL g763 ( 
.A(n_688),
.B(n_454),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_548),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_577),
.B(n_548),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_597),
.A2(n_497),
.B(n_524),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_621),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_578),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_646),
.B(n_572),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_677),
.B(n_543),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_646),
.B(n_537),
.C(n_564),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_621),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_629),
.A2(n_497),
.B(n_524),
.Y(n_774)
);

AOI21x1_ASAP7_75t_L g775 ( 
.A1(n_718),
.A2(n_512),
.B(n_563),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_669),
.B(n_564),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_733),
.B(n_543),
.Y(n_777)
);

INVx3_ASAP7_75t_SL g778 ( 
.A(n_726),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_622),
.A2(n_512),
.B1(n_543),
.B2(n_563),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_673),
.A2(n_567),
.B(n_569),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_512),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_614),
.B(n_655),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_701),
.B(n_563),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_569),
.B(n_482),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_622),
.B(n_482),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_656),
.B(n_565),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_647),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_659),
.B(n_565),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_734),
.A2(n_569),
.B(n_507),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_735),
.A2(n_507),
.B(n_565),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_601),
.A2(n_507),
.B(n_565),
.C(n_628),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_623),
.B(n_565),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_628),
.A2(n_507),
.B(n_698),
.C(n_719),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_607),
.A2(n_677),
.B1(n_708),
.B2(n_706),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_637),
.B(n_664),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_637),
.B(n_663),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_607),
.B(n_580),
.Y(n_798)
);

CKINVDCx6p67_ASAP7_75t_R g799 ( 
.A(n_626),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_674),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_735),
.A2(n_579),
.B(n_594),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_632),
.B(n_638),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_611),
.A2(n_737),
.B(n_602),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_581),
.B(n_592),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_651),
.B(n_633),
.Y(n_805)
);

AOI21xp33_ASAP7_75t_L g806 ( 
.A1(n_698),
.A2(n_679),
.B(n_683),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_613),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_681),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_682),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_736),
.Y(n_810)
);

NOR2x1_ASAP7_75t_L g811 ( 
.A(n_660),
.B(n_684),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_594),
.A2(n_697),
.B(n_699),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_711),
.B(n_643),
.C(n_700),
.Y(n_813)
);

O2A1O1Ixp5_ASAP7_75t_L g814 ( 
.A1(n_593),
.A2(n_666),
.B(n_662),
.C(n_690),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_647),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_596),
.A2(n_600),
.B(n_593),
.Y(n_816)
);

AO22x1_ASAP7_75t_L g817 ( 
.A1(n_711),
.A2(n_705),
.B1(n_694),
.B2(n_696),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_642),
.B(n_649),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_586),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_670),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_584),
.B(n_589),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_661),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_591),
.B(n_590),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_685),
.B(n_687),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_620),
.A2(n_644),
.B(n_654),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_719),
.A2(n_633),
.B(n_725),
.C(n_604),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_693),
.A2(n_657),
.B1(n_668),
.B2(n_665),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_689),
.A2(n_662),
.B(n_724),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_666),
.A2(n_606),
.B1(n_648),
.B2(n_635),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_653),
.Y(n_830)
);

OAI321xp33_ASAP7_75t_L g831 ( 
.A1(n_605),
.A2(n_610),
.A3(n_640),
.B1(n_707),
.B2(n_665),
.C(n_722),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_661),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_653),
.B(n_625),
.Y(n_833)
);

NAND3x1_ASAP7_75t_L g834 ( 
.A(n_716),
.B(n_720),
.C(n_631),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_625),
.B(n_709),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_650),
.A2(n_657),
.B1(n_640),
.B2(n_605),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_682),
.B(n_710),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_617),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_610),
.B(n_670),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_721),
.B(n_714),
.Y(n_840)
);

NAND2x1_ASAP7_75t_L g841 ( 
.A(n_736),
.B(n_675),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_639),
.A2(n_736),
.B(n_634),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_639),
.A2(n_627),
.B(n_650),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_661),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_616),
.B(n_652),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_689),
.A2(n_678),
.B(n_675),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_675),
.A2(n_702),
.B(n_703),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_658),
.B(n_675),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_713),
.A2(n_695),
.B1(n_731),
.B2(n_641),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_645),
.A2(n_732),
.B(n_704),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_703),
.B(n_729),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_715),
.B(n_723),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_703),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_717),
.A2(n_676),
.B(n_598),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_582),
.B(n_676),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_691),
.B(n_582),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_703),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_729),
.A2(n_671),
.B(n_630),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_729),
.A2(n_671),
.B(n_630),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_582),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_582),
.B(n_624),
.Y(n_861)
);

AOI33xp33_ASAP7_75t_L g862 ( 
.A1(n_582),
.A2(n_610),
.A3(n_605),
.B1(n_499),
.B2(n_458),
.B3(n_476),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_632),
.B(n_576),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_599),
.B(n_587),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_599),
.B(n_587),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_599),
.B(n_587),
.Y(n_868)
);

CKINVDCx10_ASAP7_75t_R g869 ( 
.A(n_626),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_599),
.A2(n_622),
.B(n_575),
.C(n_619),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_624),
.B(n_609),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_726),
.B(n_491),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_619),
.A2(n_599),
.B1(n_603),
.B2(n_622),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_599),
.B(n_583),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_599),
.B(n_587),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_599),
.B(n_583),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_L g878 ( 
.A1(n_646),
.A2(n_403),
.B(n_394),
.Y(n_878)
);

OAI22xp33_ASAP7_75t_L g879 ( 
.A1(n_624),
.A2(n_518),
.B1(n_612),
.B2(n_609),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_680),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_599),
.A2(n_622),
.B(n_575),
.C(n_619),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_SL g883 ( 
.A(n_688),
.B(n_494),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_661),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_599),
.B(n_583),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_621),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_680),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_599),
.B(n_587),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_619),
.A2(n_599),
.B1(n_603),
.B2(n_622),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_599),
.B(n_587),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_619),
.A2(n_599),
.B1(n_603),
.B2(n_622),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_599),
.B(n_583),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_671),
.A2(n_603),
.B(n_483),
.Y(n_896)
);

AO32x1_ASAP7_75t_L g897 ( 
.A1(n_686),
.A2(n_680),
.A3(n_591),
.B1(n_589),
.B2(n_584),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_599),
.B(n_587),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_599),
.B(n_587),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_599),
.B(n_583),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_865),
.B(n_866),
.Y(n_901)
);

BUFx12f_ASAP7_75t_L g902 ( 
.A(n_755),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_868),
.B(n_876),
.Y(n_903)
);

O2A1O1Ixp5_ASAP7_75t_L g904 ( 
.A1(n_806),
.A2(n_870),
.B(n_881),
.C(n_824),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_797),
.A2(n_878),
.B(n_899),
.C(n_898),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_775),
.A2(n_785),
.B(n_850),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_808),
.Y(n_907)
);

BUFx4f_ASAP7_75t_L g908 ( 
.A(n_778),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_L g909 ( 
.A1(n_874),
.A2(n_890),
.B(n_893),
.C(n_795),
.Y(n_909)
);

AOI21x1_ASAP7_75t_SL g910 ( 
.A1(n_786),
.A2(n_793),
.B(n_748),
.Y(n_910)
);

AO31x2_ASAP7_75t_L g911 ( 
.A1(n_828),
.A2(n_873),
.A3(n_896),
.B(n_895),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_889),
.B(n_891),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_805),
.A2(n_836),
.B(n_845),
.C(n_826),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_844),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_800),
.A2(n_862),
.B(n_867),
.C(n_863),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_741),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_746),
.A2(n_846),
.B(n_743),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_796),
.B(n_819),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_758),
.B(n_782),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_742),
.A2(n_847),
.B(n_842),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_817),
.B(n_747),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_809),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_767),
.Y(n_923)
);

OAI21x1_ASAP7_75t_L g924 ( 
.A1(n_780),
.A2(n_774),
.B(n_766),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_770),
.A2(n_882),
.B(n_885),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_888),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_745),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_739),
.B(n_871),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_892),
.A2(n_750),
.B(n_777),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_810),
.A2(n_860),
.B(n_776),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_750),
.A2(n_803),
.B(n_814),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_SL g933 ( 
.A1(n_848),
.A2(n_851),
.B(n_761),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_754),
.B(n_823),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_879),
.B(n_751),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_773),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_794),
.A2(n_827),
.B(n_831),
.C(n_861),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_844),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_875),
.B(n_877),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_810),
.A2(n_843),
.B(n_855),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_886),
.B(n_894),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_900),
.B(n_818),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_820),
.B(n_772),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_738),
.A2(n_839),
.B1(n_807),
.B2(n_856),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_816),
.A2(n_756),
.B(n_801),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_781),
.B(n_821),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_858),
.A2(n_859),
.B(n_854),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_887),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_825),
.A2(n_840),
.B(n_841),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_804),
.B(n_864),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_759),
.B(n_768),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_825),
.A2(n_812),
.B(n_779),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_769),
.A2(n_792),
.B(n_760),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_883),
.B(n_802),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_798),
.A2(n_784),
.B(n_764),
.Y(n_955)
);

AO31x2_ASAP7_75t_L g956 ( 
.A1(n_765),
.A2(n_787),
.A3(n_789),
.B(n_791),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_834),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_804),
.B(n_852),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_838),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_830),
.Y(n_960)
);

AO31x2_ASAP7_75t_L g961 ( 
.A1(n_791),
.A2(n_835),
.A3(n_833),
.B(n_897),
.Y(n_961)
);

OAI22x1_ASAP7_75t_L g962 ( 
.A1(n_864),
.A2(n_811),
.B1(n_752),
.B2(n_744),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_844),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_897),
.A2(n_749),
.A3(n_790),
.B(n_815),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_810),
.A2(n_761),
.B(n_851),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_829),
.B(n_771),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_832),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_790),
.A2(n_853),
.B(n_857),
.Y(n_968)
);

AOI21xp33_ASAP7_75t_L g969 ( 
.A1(n_753),
.A2(n_788),
.B(n_783),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_853),
.A2(n_857),
.B(n_757),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_872),
.B(n_799),
.Y(n_971)
);

AOI21xp33_ASAP7_75t_L g972 ( 
.A1(n_849),
.A2(n_757),
.B(n_884),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_832),
.A2(n_897),
.B(n_749),
.Y(n_973)
);

AO31x2_ASAP7_75t_L g974 ( 
.A1(n_749),
.A2(n_837),
.A3(n_822),
.B(n_884),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_822),
.A2(n_763),
.B(n_869),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_740),
.A2(n_762),
.B(n_671),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_755),
.B(n_574),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_865),
.B(n_866),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_796),
.B(n_898),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_755),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_775),
.A2(n_785),
.B(n_850),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_808),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_755),
.B(n_574),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_775),
.A2(n_785),
.B(n_850),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_870),
.A2(n_881),
.B(n_740),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_739),
.B(n_609),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_809),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_869),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_740),
.A2(n_762),
.B(n_671),
.Y(n_989)
);

CKINVDCx6p67_ASAP7_75t_R g990 ( 
.A(n_869),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_740),
.A2(n_762),
.B(n_671),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_865),
.B(n_866),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_820),
.B(n_772),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_755),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_L g995 ( 
.A1(n_878),
.A2(n_836),
.B(n_797),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_775),
.A2(n_785),
.B(n_850),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_808),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_796),
.B(n_898),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_870),
.A2(n_881),
.B(n_797),
.C(n_878),
.Y(n_999)
);

NOR4xp25_ASAP7_75t_L g1000 ( 
.A(n_870),
.B(n_881),
.C(n_831),
.D(n_878),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_739),
.B(n_609),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_806),
.A2(n_881),
.B(n_870),
.C(n_824),
.Y(n_1002)
);

AO31x2_ASAP7_75t_L g1003 ( 
.A1(n_870),
.A2(n_881),
.A3(n_828),
.B(n_874),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_869),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_796),
.B(n_898),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_865),
.B(n_868),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_755),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_865),
.B(n_868),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_809),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_865),
.B(n_868),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_865),
.B(n_868),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_872),
.B(n_505),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_844),
.Y(n_1014)
);

AO221x1_ASAP7_75t_L g1015 ( 
.A1(n_836),
.A2(n_893),
.B1(n_890),
.B2(n_874),
.C(n_879),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_755),
.B(n_574),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_951),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_988),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_901),
.B(n_903),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_L g1020 ( 
.A(n_987),
.B(n_1010),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_986),
.B(n_1001),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_918),
.B(n_977),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_950),
.B(n_921),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_912),
.A2(n_978),
.B1(n_992),
.B2(n_1009),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_913),
.A2(n_995),
.B(n_905),
.C(n_999),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_980),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_SL g1027 ( 
.A1(n_973),
.A2(n_944),
.B(n_941),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_929),
.B(n_1006),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1015),
.A2(n_935),
.B1(n_979),
.B2(n_998),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_928),
.B(n_1005),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_953),
.A2(n_945),
.B(n_930),
.Y(n_1031)
);

BUFx4_ASAP7_75t_SL g1032 ( 
.A(n_1004),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1011),
.B(n_1012),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_990),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_967),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_954),
.A2(n_919),
.B1(n_944),
.B2(n_992),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_916),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_908),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_934),
.B(n_946),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_914),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_957),
.A2(n_958),
.B1(n_921),
.B2(n_928),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_909),
.B(n_985),
.C(n_904),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_926),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_908),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1000),
.B(n_942),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_914),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_902),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_983),
.B(n_1016),
.Y(n_1048)
);

BUFx12f_ASAP7_75t_L g1049 ( 
.A(n_922),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1000),
.B(n_939),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_980),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_994),
.B(n_921),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_994),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_1008),
.Y(n_1054)
);

INVx8_ASAP7_75t_L g1055 ( 
.A(n_938),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_927),
.Y(n_1056)
);

OR2x2_ASAP7_75t_SL g1057 ( 
.A(n_971),
.B(n_907),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_963),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_937),
.B(n_915),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_982),
.B(n_997),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_938),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_933),
.B(n_975),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_936),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_938),
.B(n_1014),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_1007),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_959),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_923),
.B(n_948),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_960),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_943),
.B(n_993),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1013),
.B(n_993),
.Y(n_1070)
);

AND3x1_ASAP7_75t_SL g1071 ( 
.A(n_962),
.B(n_943),
.C(n_1002),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1007),
.B(n_1014),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_SL g1073 ( 
.A1(n_932),
.A2(n_955),
.B(n_969),
.C(n_972),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_970),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_940),
.A2(n_949),
.B(n_917),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_974),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_974),
.Y(n_1077)
);

CKINVDCx11_ASAP7_75t_R g1078 ( 
.A(n_910),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_968),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_965),
.B(n_920),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_961),
.Y(n_1081)
);

OAI321xp33_ASAP7_75t_L g1082 ( 
.A1(n_925),
.A2(n_1003),
.A3(n_931),
.B1(n_911),
.B2(n_961),
.C(n_952),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_L g1083 ( 
.A(n_972),
.B(n_969),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_911),
.B(n_956),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_911),
.B(n_956),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_956),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_964),
.Y(n_1087)
);

AO22x2_ASAP7_75t_L g1088 ( 
.A1(n_964),
.A2(n_947),
.B1(n_906),
.B2(n_981),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_984),
.B(n_996),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_SL g1090 ( 
.A(n_924),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_967),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_901),
.Y(n_1092)
);

OR2x2_ASAP7_75t_SL g1093 ( 
.A(n_971),
.B(n_485),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_L g1094 ( 
.A(n_901),
.B(n_870),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_951),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_916),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_951),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_901),
.A2(n_878),
.B(n_403),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_914),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_901),
.B(n_865),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_901),
.B(n_865),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_986),
.B(n_609),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_980),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_967),
.B(n_966),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_951),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_914),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_912),
.A2(n_619),
.B1(n_866),
.B2(n_865),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_908),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_976),
.A2(n_991),
.B(n_989),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_901),
.B(n_865),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_912),
.A2(n_619),
.B1(n_866),
.B2(n_865),
.Y(n_1111)
);

OR2x2_ASAP7_75t_SL g1112 ( 
.A(n_971),
.B(n_485),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_951),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_951),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_951),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_901),
.B(n_865),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_907),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_901),
.B(n_865),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_901),
.B(n_865),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1015),
.A2(n_878),
.B1(n_797),
.B2(n_836),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_913),
.A2(n_878),
.B(n_881),
.C(n_870),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_914),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_950),
.B(n_921),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_950),
.B(n_921),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_929),
.B(n_595),
.Y(n_1125)
);

NAND2x1_ASAP7_75t_L g1126 ( 
.A(n_967),
.B(n_832),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_909),
.A2(n_806),
.B(n_881),
.C(n_870),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_901),
.B(n_865),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_986),
.B(n_609),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_914),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_951),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_986),
.B(n_609),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1021),
.A2(n_1125),
.B1(n_1098),
.B2(n_1120),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_1055),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1056),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_1055),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1028),
.B(n_1092),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_SL g1138 ( 
.A1(n_1102),
.A2(n_1132),
.B1(n_1129),
.B2(n_1042),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1026),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1055),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1036),
.A2(n_1039),
.B1(n_1119),
.B2(n_1118),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1039),
.A2(n_1128),
.B1(n_1119),
.B2(n_1118),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1068),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1098),
.A2(n_1041),
.B1(n_1042),
.B2(n_1094),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1121),
.A2(n_1025),
.B(n_1070),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1051),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1043),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1023),
.A2(n_1123),
.B1(n_1124),
.B2(n_1031),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_1127),
.A2(n_1109),
.B(n_1082),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_SL g1151 ( 
.A(n_1018),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1052),
.A2(n_1124),
.B1(n_1023),
.B2(n_1123),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1048),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1046),
.Y(n_1154)
);

BUFx2_ASAP7_75t_SL g1155 ( 
.A(n_1040),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1053),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1066),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1027),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1024),
.B(n_1019),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1019),
.B(n_1033),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_1059),
.A2(n_1033),
.B1(n_1116),
.B2(n_1101),
.Y(n_1161)
);

OAI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1100),
.A2(n_1128),
.B1(n_1116),
.B2(n_1110),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1017),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1037),
.Y(n_1164)
);

OAI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1100),
.A2(n_1101),
.B1(n_1110),
.B2(n_1022),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1095),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1059),
.A2(n_1107),
.B1(n_1111),
.B2(n_1030),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1065),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1053),
.A2(n_1103),
.B1(n_1107),
.B2(n_1111),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1045),
.B(n_1050),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1097),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1113),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1131),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1088),
.A2(n_1080),
.B(n_1085),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1032),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1046),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1045),
.B(n_1050),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1105),
.Y(n_1178)
);

CKINVDCx11_ASAP7_75t_R g1179 ( 
.A(n_1049),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1096),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1103),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1084),
.B(n_1081),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1062),
.A2(n_1069),
.B1(n_1071),
.B2(n_1020),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1114),
.B(n_1115),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1072),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1083),
.A2(n_1089),
.B(n_1073),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1099),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1064),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1088),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1086),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1057),
.A2(n_1117),
.B1(n_1063),
.B2(n_1112),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1067),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1093),
.A2(n_1058),
.B1(n_1074),
.B2(n_1062),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1062),
.A2(n_1078),
.B1(n_1104),
.B2(n_1047),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1060),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1126),
.A2(n_1090),
.B(n_1104),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1108),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1034),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1099),
.Y(n_1200)
);

AND2x2_ASAP7_75t_SL g1201 ( 
.A(n_1104),
.B(n_1090),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1086),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1099),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1104),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1076),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1044),
.A2(n_1086),
.B1(n_1035),
.B2(n_1091),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_SL g1207 ( 
.A(n_1054),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1065),
.B(n_1061),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1065),
.Y(n_1209)
);

INVx6_ASAP7_75t_L g1210 ( 
.A(n_1040),
.Y(n_1210)
);

BUFx2_ASAP7_75t_R g1211 ( 
.A(n_1061),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1079),
.A2(n_1077),
.B(n_1087),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1106),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1106),
.Y(n_1214)
);

INVx8_ASAP7_75t_L g1215 ( 
.A(n_1106),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1122),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1122),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1130),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1130),
.A2(n_865),
.B1(n_868),
.B2(n_866),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1056),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1056),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1080),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1026),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1056),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1056),
.Y(n_1225)
);

BUFx8_ASAP7_75t_L g1226 ( 
.A(n_1018),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1056),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1021),
.A2(n_878),
.B1(n_797),
.B2(n_813),
.Y(n_1228)
);

CKINVDCx6p67_ASAP7_75t_R g1229 ( 
.A(n_1018),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1029),
.B(n_1092),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1075),
.A2(n_924),
.B(n_917),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1170),
.B(n_1177),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1205),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1201),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1159),
.B(n_1143),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1170),
.B(n_1177),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1189),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1212),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1212),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1174),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1162),
.A2(n_1142),
.B(n_1231),
.Y(n_1241)
);

CKINVDCx6p67_ASAP7_75t_R g1242 ( 
.A(n_1179),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1182),
.B(n_1159),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1158),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1158),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1182),
.B(n_1139),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1204),
.B(n_1197),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1175),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1139),
.B(n_1167),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1186),
.A2(n_1169),
.B(n_1190),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1186),
.A2(n_1202),
.B(n_1190),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1150),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1153),
.B(n_1137),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1138),
.B(n_1160),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1186),
.A2(n_1202),
.B(n_1146),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1145),
.A2(n_1204),
.B(n_1230),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1175),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1222),
.B(n_1183),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1161),
.B(n_1230),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1165),
.B(n_1133),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1148),
.A2(n_1157),
.B(n_1228),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1201),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1206),
.A2(n_1219),
.B(n_1194),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1150),
.A2(n_1195),
.B(n_1149),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1150),
.B(n_1144),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1220),
.B(n_1225),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1191),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1135),
.A2(n_1224),
.B(n_1221),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1210),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1156),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1193),
.B(n_1198),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1181),
.B(n_1185),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1178),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1163),
.A2(n_1172),
.B(n_1173),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1184),
.B(n_1171),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1188),
.A2(n_1192),
.B(n_1166),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1191),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1196),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1152),
.B(n_1218),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1208),
.B(n_1216),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1266),
.B(n_1232),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1266),
.B(n_1214),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1254),
.A2(n_1179),
.B1(n_1229),
.B2(n_1191),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1251),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1240),
.B(n_1217),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1240),
.B(n_1214),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1232),
.B(n_1176),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1236),
.B(n_1176),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1236),
.B(n_1176),
.Y(n_1292)
);

OAI31xp33_ASAP7_75t_L g1293 ( 
.A1(n_1260),
.A2(n_1164),
.A3(n_1180),
.B(n_1209),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1247),
.B(n_1155),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1260),
.B(n_1180),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1245),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1243),
.B(n_1154),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1243),
.B(n_1154),
.Y(n_1298)
);

NOR2x1_ASAP7_75t_SL g1299 ( 
.A(n_1247),
.B(n_1155),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1256),
.B(n_1252),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1247),
.B(n_1168),
.Y(n_1301)
);

NAND2x1_ASAP7_75t_L g1302 ( 
.A(n_1247),
.B(n_1210),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1247),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1247),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1256),
.B(n_1200),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1248),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1256),
.B(n_1200),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1256),
.B(n_1154),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1241),
.A2(n_1215),
.B(n_1168),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_1267),
.B(n_1262),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1250),
.B(n_1187),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1293),
.B(n_1253),
.C(n_1241),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1284),
.B(n_1237),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1284),
.B(n_1237),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1293),
.B(n_1235),
.C(n_1261),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1295),
.B(n_1273),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1284),
.B(n_1255),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1305),
.B(n_1246),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1305),
.B(n_1246),
.Y(n_1319)
);

NOR3xp33_ASAP7_75t_L g1320 ( 
.A(n_1309),
.B(n_1276),
.C(n_1281),
.Y(n_1320)
);

AND4x1_ASAP7_75t_L g1321 ( 
.A(n_1286),
.B(n_1249),
.C(n_1259),
.D(n_1242),
.Y(n_1321)
);

NAND4xp25_ASAP7_75t_L g1322 ( 
.A(n_1286),
.B(n_1265),
.C(n_1274),
.D(n_1276),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1301),
.A2(n_1258),
.B1(n_1259),
.B2(n_1262),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1309),
.A2(n_1249),
.B(n_1264),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1300),
.A2(n_1281),
.B(n_1274),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1311),
.B(n_1261),
.C(n_1282),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1302),
.B(n_1283),
.C(n_1271),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1304),
.A2(n_1262),
.B1(n_1234),
.B2(n_1258),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1290),
.B(n_1265),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1290),
.B(n_1275),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1303),
.A2(n_1277),
.B1(n_1280),
.B2(n_1282),
.C(n_1244),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1294),
.A2(n_1234),
.B1(n_1262),
.B2(n_1211),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1311),
.B(n_1261),
.C(n_1270),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1294),
.A2(n_1234),
.B1(n_1262),
.B2(n_1242),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1291),
.B(n_1270),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1291),
.B(n_1233),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1311),
.B(n_1261),
.C(n_1244),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1304),
.B(n_1271),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1291),
.B(n_1292),
.Y(n_1340)
);

AOI221xp5_ASAP7_75t_L g1341 ( 
.A1(n_1303),
.A2(n_1277),
.B1(n_1280),
.B2(n_1283),
.C(n_1278),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1307),
.B(n_1250),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1307),
.B(n_1250),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1292),
.B(n_1233),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1294),
.B(n_1238),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1301),
.A2(n_1258),
.B1(n_1263),
.B2(n_1242),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1292),
.B(n_1269),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1308),
.B(n_1238),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1288),
.A2(n_1264),
.B(n_1261),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1294),
.A2(n_1207),
.B1(n_1268),
.B2(n_1279),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1297),
.B(n_1269),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1297),
.B(n_1268),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1308),
.B(n_1239),
.Y(n_1353)
);

OA211x2_ASAP7_75t_L g1354 ( 
.A1(n_1302),
.A2(n_1310),
.B(n_1299),
.C(n_1304),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1342),
.B(n_1343),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1348),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1347),
.B(n_1300),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_SL g1358 ( 
.A(n_1312),
.B(n_1304),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1353),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1316),
.B(n_1312),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1353),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1345),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1351),
.B(n_1287),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1345),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1317),
.B(n_1318),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1314),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1338),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1327),
.B(n_1287),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_1325),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1322),
.B(n_1278),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1319),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1324),
.B(n_1304),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1349),
.B(n_1304),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1340),
.B(n_1304),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1334),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1331),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1336),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1354),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1320),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1339),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1335),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1330),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1359),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1357),
.B(n_1337),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1366),
.B(n_1294),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1366),
.B(n_1294),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1381),
.B(n_1326),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1366),
.B(n_1294),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1380),
.B(n_1299),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1381),
.B(n_1341),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1359),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1370),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1356),
.B(n_1329),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1356),
.B(n_1352),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1362),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1357),
.B(n_1344),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1356),
.B(n_1328),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1326),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1360),
.B(n_1332),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1384),
.B(n_1379),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1372),
.A2(n_1315),
.B(n_1321),
.Y(n_1403)
);

INVx3_ASAP7_75t_R g1404 ( 
.A(n_1383),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1384),
.B(n_1298),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1362),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1359),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1380),
.B(n_1362),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1361),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1364),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1361),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1365),
.B(n_1302),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1373),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1357),
.B(n_1289),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1365),
.B(n_1285),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1298),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1368),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1365),
.B(n_1285),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1377),
.B(n_1296),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1379),
.B(n_1298),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1376),
.B(n_1285),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1404),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1396),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1403),
.A2(n_1383),
.B1(n_1372),
.B2(n_1358),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1369),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1400),
.B(n_1369),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1396),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1383),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1409),
.B(n_1391),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1385),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1392),
.B(n_1378),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1395),
.B(n_1355),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1392),
.B(n_1378),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1393),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1393),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1408),
.B(n_1370),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1395),
.B(n_1423),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1407),
.Y(n_1441)
);

NOR3xp33_ASAP7_75t_L g1442 ( 
.A(n_1389),
.B(n_1350),
.C(n_1374),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1394),
.B(n_1370),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1409),
.B(n_1380),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1394),
.B(n_1420),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1399),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1420),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1407),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1414),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1423),
.B(n_1355),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1404),
.A2(n_1358),
.B1(n_1371),
.B2(n_1333),
.Y(n_1452)
);

INVxp33_ASAP7_75t_L g1453 ( 
.A(n_1409),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_L g1454 ( 
.A(n_1397),
.B(n_1371),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1414),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1410),
.B(n_1363),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1410),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1405),
.B(n_1378),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1414),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1413),
.B(n_1355),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1412),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1412),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1415),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1417),
.B(n_1378),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1461),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1461),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1425),
.B(n_1386),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1432),
.B(n_1409),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1440),
.B(n_1387),
.Y(n_1470)
);

INVx3_ASAP7_75t_SL g1471 ( 
.A(n_1444),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1431),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1432),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1430),
.B(n_1386),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1457),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1432),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1398),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1463),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1424),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1437),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1454),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1427),
.B(n_1380),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1428),
.B(n_1402),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1429),
.B(n_1447),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1444),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1454),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1438),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1444),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1443),
.B(n_1268),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1426),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1433),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1451),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1452),
.B(n_1229),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1445),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1434),
.B(n_1398),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1436),
.B(n_1415),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1440),
.B(n_1422),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1445),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1481),
.B(n_1487),
.Y(n_1501)
);

NOR2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1472),
.B(n_1279),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1491),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1491),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1471),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1495),
.A2(n_1321),
.B(n_1442),
.Y(n_1506)
);

AOI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1472),
.A2(n_1439),
.B1(n_1443),
.B2(n_1453),
.C(n_1464),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1479),
.B(n_1500),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1494),
.B(n_1435),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1473),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1471),
.A2(n_1453),
.B1(n_1439),
.B2(n_1406),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1484),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1466),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1482),
.A2(n_1464),
.B1(n_1435),
.B2(n_1374),
.C(n_1375),
.Y(n_1516)
);

CKINVDCx16_ASAP7_75t_R g1517 ( 
.A(n_1495),
.Y(n_1517)
);

AOI222xp33_ASAP7_75t_L g1518 ( 
.A1(n_1479),
.A2(n_1374),
.B1(n_1375),
.B2(n_1451),
.C1(n_1450),
.C2(n_1460),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1473),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1500),
.A2(n_1375),
.B1(n_1397),
.B2(n_1406),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1496),
.B(n_1476),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1490),
.A2(n_1391),
.B1(n_1354),
.B2(n_1382),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1496),
.B(n_1450),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1485),
.A2(n_1279),
.B(n_1411),
.C(n_1164),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1469),
.B(n_1391),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1505),
.B(n_1469),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1517),
.B(n_1489),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1503),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1504),
.Y(n_1529)
);

NOR2xp67_ASAP7_75t_SL g1530 ( 
.A(n_1508),
.B(n_1257),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1509),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1501),
.B(n_1485),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1502),
.Y(n_1533)
);

CKINVDCx16_ASAP7_75t_R g1534 ( 
.A(n_1521),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1510),
.B(n_1519),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1506),
.B(n_1490),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1507),
.B(n_1486),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1483),
.Y(n_1538)
);

NOR3xp33_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1489),
.C(n_1483),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1523),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1525),
.B(n_1490),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1512),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1513),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1524),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1534),
.B(n_1514),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1531),
.Y(n_1546)
);

NOR3xp33_ASAP7_75t_L g1547 ( 
.A(n_1527),
.B(n_1516),
.C(n_1515),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1530),
.B(n_1477),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1538),
.A2(n_1516),
.B1(n_1524),
.B2(n_1520),
.C(n_1475),
.Y(n_1549)
);

NAND4xp25_ASAP7_75t_L g1550 ( 
.A(n_1532),
.B(n_1518),
.C(n_1522),
.D(n_1478),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1527),
.A2(n_1467),
.B(n_1493),
.C(n_1492),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1470),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1537),
.A2(n_1474),
.B1(n_1468),
.B2(n_1497),
.C(n_1498),
.Y(n_1553)
);

OAI211xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1536),
.A2(n_1499),
.B(n_1456),
.C(n_1465),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1546),
.B(n_1528),
.Y(n_1557)
);

NOR3xp33_ASAP7_75t_L g1558 ( 
.A(n_1545),
.B(n_1535),
.C(n_1540),
.Y(n_1558)
);

NOR3xp33_ASAP7_75t_SL g1559 ( 
.A(n_1550),
.B(n_1544),
.C(n_1529),
.Y(n_1559)
);

NOR2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1555),
.B(n_1542),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1551),
.Y(n_1561)
);

XNOR2x1_ASAP7_75t_SL g1562 ( 
.A(n_1552),
.B(n_1533),
.Y(n_1562)
);

AOI211x1_ASAP7_75t_L g1563 ( 
.A1(n_1554),
.A2(n_1541),
.B(n_1543),
.C(n_1441),
.Y(n_1563)
);

NOR3x1_ASAP7_75t_L g1564 ( 
.A(n_1547),
.B(n_1533),
.C(n_1411),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1559),
.B(n_1549),
.C(n_1539),
.Y(n_1565)
);

OAI21xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1562),
.A2(n_1541),
.B(n_1553),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1561),
.A2(n_1391),
.B(n_1456),
.C(n_1226),
.Y(n_1567)
);

AOI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1563),
.A2(n_1449),
.B1(n_1459),
.B2(n_1455),
.C(n_1448),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1557),
.B(n_1387),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1569),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1565),
.A2(n_1566),
.B1(n_1556),
.B2(n_1558),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1567),
.B(n_1560),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1568),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1565),
.A2(n_1564),
.B1(n_1449),
.B2(n_1459),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1565),
.A2(n_1455),
.B1(n_1364),
.B2(n_1382),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1571),
.A2(n_1570),
.B1(n_1572),
.B2(n_1573),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1574),
.B(n_1226),
.C(n_1151),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1575),
.B(n_1199),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1570),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1570),
.B(n_1458),
.Y(n_1580)
);

NAND5xp2_ASAP7_75t_L g1581 ( 
.A(n_1576),
.B(n_1226),
.C(n_1199),
.D(n_1346),
.E(n_1323),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1579),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1578),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1582),
.Y(n_1584)
);

AOI211xp5_ASAP7_75t_L g1585 ( 
.A1(n_1584),
.A2(n_1577),
.B(n_1583),
.C(n_1581),
.Y(n_1585)
);

AO21x2_ASAP7_75t_L g1586 ( 
.A1(n_1585),
.A2(n_1580),
.B(n_1462),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1586),
.A2(n_1199),
.B1(n_1203),
.B2(n_1462),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1587),
.A2(n_1586),
.B(n_1382),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1588),
.A2(n_1364),
.B(n_1388),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_R g1590 ( 
.A1(n_1589),
.A2(n_1421),
.B1(n_1418),
.B2(n_1367),
.Y(n_1590)
);

AOI322xp5_ASAP7_75t_L g1591 ( 
.A1(n_1589),
.A2(n_1419),
.A3(n_1416),
.B1(n_1388),
.B2(n_1390),
.C1(n_1421),
.C2(n_1376),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1590),
.A2(n_1141),
.B1(n_1215),
.B2(n_1134),
.C(n_1136),
.Y(n_1592)
);

AOI211xp5_ASAP7_75t_L g1593 ( 
.A1(n_1592),
.A2(n_1591),
.B(n_1141),
.C(n_1213),
.Y(n_1593)
);


endmodule