module fake_netlist_6_4773_n_843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_843;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_57),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_160),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_43),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_25),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_79),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_121),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_40),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_120),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_139),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_122),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_28),
.B(n_126),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_31),
.B(n_157),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_131),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_76),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_53),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_64),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_98),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_112),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_104),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_136),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_41),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_82),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_167),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_190),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

CKINVDCx6p67_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

OAI22x1_ASAP7_75t_SL g244 ( 
.A1(n_223),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_178),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_217),
.Y(n_246)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_18),
.Y(n_247)
);

CKINVDCx11_ASAP7_75t_R g248 ( 
.A(n_186),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_19),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_1),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_189),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

CKINVDCx9p33_ASAP7_75t_R g261 ( 
.A(n_179),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_20),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_21),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_4),
.B(n_5),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_22),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_198),
.A2(n_5),
.B(n_6),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_174),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_23),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_224),
.A2(n_6),
.B(n_7),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_175),
.B(n_7),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_176),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_182),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_200),
.B(n_8),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_9),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_181),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_185),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

AND3x2_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_9),
.C(n_10),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_245),
.B(n_183),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_193),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_288),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_248),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_248),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_253),
.Y(n_306)
);

BUFx6f_ASAP7_75t_SL g307 ( 
.A(n_253),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_242),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_243),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_R g312 ( 
.A(n_282),
.B(n_188),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_270),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_288),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_284),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_257),
.B(n_196),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_290),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_261),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_252),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_266),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_258),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_R g336 ( 
.A(n_281),
.B(n_191),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_286),
.B(n_279),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_279),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_277),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_336),
.B(n_250),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_271),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_271),
.Y(n_347)
);

NAND2x1p5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_250),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_321),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_283),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_250),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_336),
.B(n_271),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_295),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_251),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_251),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_278),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_247),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_247),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_278),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_278),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_315),
.B(n_240),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_268),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_295),
.B(n_268),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_277),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_294),
.B(n_299),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_254),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_292),
.B(n_206),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_281),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_277),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_314),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_312),
.B(n_203),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_293),
.B(n_240),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_302),
.B(n_244),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_333),
.B(n_254),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_340),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_309),
.B(n_204),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_298),
.B(n_281),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_265),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_262),
.C(n_249),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_326),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_292),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_277),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_291),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_303),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_304),
.B(n_209),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_295),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_300),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_306),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_272),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_310),
.B(n_254),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_269),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_246),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_369),
.Y(n_415)
);

O2A1O1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_362),
.A2(n_246),
.B(n_265),
.C(n_280),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_350),
.B(n_280),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_269),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_SL g422 ( 
.A(n_395),
.B(n_213),
.C(n_211),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_280),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_214),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_272),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_361),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_351),
.B(n_219),
.Y(n_432)
);

OR2x2_ASAP7_75t_SL g433 ( 
.A(n_401),
.B(n_11),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

O2A1O1Ixp5_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_345),
.B(n_347),
.C(n_367),
.Y(n_435)
);

O2A1O1Ixp5_ASAP7_75t_L g436 ( 
.A1(n_370),
.A2(n_267),
.B(n_266),
.C(n_264),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_344),
.B(n_267),
.Y(n_438)
);

NOR2x2_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_11),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_376),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_355),
.A2(n_234),
.B1(n_221),
.B2(n_222),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_398),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_374),
.B(n_375),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_379),
.A2(n_409),
.B1(n_347),
.B2(n_345),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_363),
.A2(n_264),
.B1(n_247),
.B2(n_267),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_380),
.B(n_220),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_378),
.B(n_24),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_356),
.B(n_227),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_360),
.B(n_228),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_387),
.A2(n_403),
.B1(n_406),
.B2(n_364),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_383),
.B(n_229),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_404),
.B(n_12),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_379),
.A2(n_238),
.B1(n_237),
.B2(n_235),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_SL g460 ( 
.A(n_405),
.B(n_233),
.C(n_14),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_348),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_348),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_372),
.B(n_13),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_399),
.B(n_254),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_385),
.B(n_254),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_14),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_368),
.B(n_371),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_247),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_390),
.B(n_247),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_400),
.B(n_264),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_365),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_SL g479 ( 
.A(n_440),
.B(n_392),
.C(n_389),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_15),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_424),
.A2(n_264),
.B(n_247),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_432),
.A2(n_264),
.B1(n_99),
.B2(n_100),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_418),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_15),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_SL g490 ( 
.A(n_454),
.B(n_16),
.C(n_17),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_461),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

O2A1O1Ixp5_ASAP7_75t_L g493 ( 
.A1(n_426),
.A2(n_264),
.B(n_26),
.C(n_27),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_101),
.C(n_29),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

O2A1O1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_417),
.A2(n_17),
.B(n_30),
.C(n_34),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_470),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_437),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_477),
.B(n_42),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_44),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_461),
.B(n_46),
.Y(n_501)
);

NOR3xp33_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_50),
.C(n_51),
.Y(n_502)
);

NAND2x1p5_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_54),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_172),
.B(n_58),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_426),
.A2(n_412),
.B(n_435),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_429),
.B(n_56),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_467),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_446),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_458),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_425),
.A2(n_67),
.B(n_68),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_446),
.B(n_70),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_436),
.A2(n_170),
.B(n_72),
.Y(n_513)
);

OAI22x1_ASAP7_75t_L g514 ( 
.A1(n_459),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_429),
.B(n_75),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

BUFx2_ASAP7_75t_SL g517 ( 
.A(n_428),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_462),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_472),
.A2(n_81),
.B(n_84),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_443),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_473),
.A2(n_86),
.B(n_87),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_88),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_449),
.A2(n_89),
.B(n_90),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_93),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_SL g530 ( 
.A1(n_438),
.A2(n_169),
.B(n_95),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_422),
.B(n_94),
.C(n_96),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_416),
.A2(n_102),
.B(n_103),
.C(n_105),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_471),
.A2(n_106),
.B(n_107),
.Y(n_533)
);

OR2x6_ASAP7_75t_SL g534 ( 
.A(n_439),
.B(n_108),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_109),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_505),
.A2(n_420),
.B(n_431),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_500),
.A2(n_448),
.B(n_421),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_513),
.A2(n_420),
.B(n_431),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_504),
.A2(n_475),
.B(n_444),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_491),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_484),
.B(n_469),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_485),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_454),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_482),
.A2(n_444),
.B(n_450),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_524),
.A2(n_450),
.B(n_468),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_486),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_500),
.A2(n_421),
.B(n_455),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_534),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_495),
.B(n_466),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_516),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_527),
.A2(n_453),
.B(n_441),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_527),
.A2(n_441),
.B(n_460),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_519),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_492),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

AOI22x1_ASAP7_75t_L g559 ( 
.A1(n_514),
.A2(n_433),
.B1(n_456),
.B2(n_114),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

BUFx4_ASAP7_75t_SL g561 ( 
.A(n_531),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_517),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_508),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

OAI21x1_ASAP7_75t_SL g565 ( 
.A1(n_512),
.A2(n_456),
.B(n_113),
.Y(n_565)
);

AOI21xp33_ASAP7_75t_L g566 ( 
.A1(n_481),
.A2(n_111),
.B(n_115),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_489),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_523),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_535),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

AO21x2_ASAP7_75t_L g573 ( 
.A1(n_512),
.A2(n_116),
.B(n_117),
.Y(n_573)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_494),
.A2(n_118),
.B(n_119),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_503),
.Y(n_576)
);

AOI22x1_ASAP7_75t_L g577 ( 
.A1(n_520),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

BUFx24_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

AOI21x1_ASAP7_75t_L g580 ( 
.A1(n_501),
.A2(n_128),
.B(n_130),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_528),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_525),
.B(n_521),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_493),
.A2(n_133),
.B(n_137),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_548),
.Y(n_584)
);

CKINVDCx6p67_ASAP7_75t_R g585 ( 
.A(n_538),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_570),
.A2(n_506),
.B1(n_502),
.B2(n_531),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_564),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_563),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_539),
.A2(n_511),
.B(n_494),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_570),
.A2(n_498),
.B1(n_483),
.B2(n_515),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_563),
.Y(n_593)
);

BUFx5_ASAP7_75t_L g594 ( 
.A(n_579),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

BUFx8_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_567),
.B(n_582),
.Y(n_598)
);

AOI222xp33_ASAP7_75t_L g599 ( 
.A1(n_545),
.A2(n_568),
.B1(n_550),
.B2(n_572),
.C1(n_542),
.C2(n_575),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_579),
.A2(n_490),
.B1(n_479),
.B2(n_509),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_571),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_564),
.B(n_518),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_581),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_559),
.A2(n_526),
.B1(n_533),
.B2(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_544),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_569),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_542),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_551),
.A2(n_530),
.B1(n_496),
.B2(n_532),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_542),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_541),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_557),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_552),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_558),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_562),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_540),
.A2(n_507),
.B(n_140),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_554),
.A2(n_138),
.B(n_142),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_552),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_556),
.B(n_148),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_555),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_560),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_576),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_596),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_555),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_605),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_588),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_585),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_584),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_595),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_591),
.B(n_564),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_599),
.B(n_578),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_603),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_599),
.B(n_578),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_598),
.B(n_578),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_597),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_605),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_588),
.B(n_576),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_601),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_586),
.A2(n_609),
.B(n_592),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_591),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_607),
.B(n_578),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_611),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_576),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_589),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_611),
.B(n_576),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_612),
.B(n_565),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_611),
.B(n_580),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_613),
.B(n_573),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_593),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_615),
.Y(n_655)
);

AO31x2_ASAP7_75t_L g656 ( 
.A1(n_600),
.A2(n_540),
.A3(n_554),
.B(n_583),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_611),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_600),
.A2(n_566),
.B1(n_549),
.B2(n_574),
.Y(n_658)
);

BUFx10_ASAP7_75t_L g659 ( 
.A(n_619),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_594),
.B(n_537),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_592),
.A2(n_577),
.B1(n_574),
.B2(n_573),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_616),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_622),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_583),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_616),
.Y(n_665)
);

CKINVDCx16_ASAP7_75t_R g666 ( 
.A(n_606),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_586),
.A2(n_561),
.B1(n_547),
.B2(n_162),
.Y(n_667)
);

INVx4_ASAP7_75t_R g668 ( 
.A(n_594),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_SL g669 ( 
.A(n_604),
.B(n_561),
.C(n_547),
.Y(n_669)
);

BUFx4f_ASAP7_75t_SL g670 ( 
.A(n_614),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_625),
.B(n_546),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_608),
.B(n_546),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_SL g673 ( 
.A1(n_594),
.A2(n_536),
.B1(n_161),
.B2(n_164),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_620),
.B(n_156),
.Y(n_674)
);

NOR2x1_ASAP7_75t_L g675 ( 
.A(n_587),
.B(n_536),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_623),
.B(n_165),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_650),
.B(n_646),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_637),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_650),
.B(n_587),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_629),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_635),
.B(n_618),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_638),
.B(n_618),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_671),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_649),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_653),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_644),
.B(n_594),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_664),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_648),
.B(n_623),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_645),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_632),
.B(n_624),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_633),
.B(n_624),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_643),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_639),
.B(n_609),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_654),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_667),
.A2(n_604),
.B1(n_602),
.B2(n_617),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_675),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_656),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_675),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_672),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_672),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_634),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_660),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_655),
.B(n_617),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_663),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_669),
.B(n_602),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_668),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_662),
.B(n_626),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_665),
.B(n_626),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_641),
.B(n_590),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_677),
.B(n_658),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_679),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_677),
.B(n_661),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_686),
.B(n_630),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_701),
.B(n_651),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_712),
.B(n_630),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_697),
.B(n_651),
.C(n_676),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_678),
.B(n_657),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_686),
.B(n_666),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_678),
.B(n_657),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_712),
.B(n_634),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_679),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_688),
.B(n_666),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_704),
.B(n_652),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_696),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_681),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_685),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_701),
.B(n_657),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_678),
.B(n_659),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_709),
.B(n_659),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_693),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_701),
.B(n_652),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_694),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_694),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_704),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_684),
.B(n_673),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_739),
.B(n_682),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_718),
.B(n_683),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_729),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_714),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_737),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_718),
.B(n_683),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_727),
.B(n_682),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_717),
.B(n_707),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_724),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_721),
.B(n_698),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_738),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_730),
.Y(n_753)
);

NOR2x1_ASAP7_75t_L g754 ( 
.A(n_719),
.B(n_700),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_720),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_728),
.B(n_702),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_735),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_741),
.B(n_698),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_732),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_719),
.A2(n_695),
.B1(n_687),
.B2(n_692),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_731),
.Y(n_761)
);

OA222x2_ASAP7_75t_L g762 ( 
.A1(n_754),
.A2(n_713),
.B1(n_715),
.B2(n_726),
.C1(n_708),
.C2(n_710),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_756),
.B(n_690),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_755),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_744),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_743),
.B(n_716),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_758),
.Y(n_767)
);

NAND4xp75_ASAP7_75t_L g768 ( 
.A(n_749),
.B(n_707),
.C(n_695),
.D(n_692),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

NOR2x1p5_ASAP7_75t_L g770 ( 
.A(n_747),
.B(n_690),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_750),
.Y(n_771)
);

AND4x1_ASAP7_75t_L g772 ( 
.A(n_760),
.B(n_740),
.C(n_734),
.D(n_710),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_748),
.B(n_726),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_742),
.B(n_725),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_772),
.A2(n_760),
.B(n_748),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_749),
.B1(n_717),
.B2(n_691),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_769),
.B(n_742),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_765),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_770),
.B(n_750),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_L g781 ( 
.A1(n_775),
.A2(n_774),
.B(n_767),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_779),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

OAI21xp33_ASAP7_75t_SL g784 ( 
.A1(n_777),
.A2(n_769),
.B(n_762),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_780),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_784),
.B(n_776),
.C(n_777),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_785),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_781),
.B(n_763),
.C(n_767),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_782),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_787),
.B(n_783),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_786),
.B(n_636),
.Y(n_791)
);

OAI222xp33_ASAP7_75t_L g792 ( 
.A1(n_791),
.A2(n_789),
.B1(n_764),
.B2(n_788),
.C1(n_766),
.C2(n_751),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_790),
.A2(n_627),
.B(n_631),
.Y(n_793)
);

OAI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_791),
.A2(n_740),
.B(n_713),
.C(n_771),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_792),
.A2(n_670),
.B1(n_608),
.B2(n_642),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_794),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_793),
.B(n_711),
.Y(n_797)
);

NOR2x1_ASAP7_75t_L g798 ( 
.A(n_793),
.B(n_711),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_794),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_792),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_795),
.B(n_731),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_796),
.Y(n_802)
);

AOI221xp5_ASAP7_75t_L g803 ( 
.A1(n_800),
.A2(n_799),
.B1(n_798),
.B2(n_797),
.C(n_709),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_800),
.A2(n_758),
.B(n_706),
.Y(n_804)
);

NOR2x1_ASAP7_75t_L g805 ( 
.A(n_800),
.B(n_674),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_797),
.B(n_722),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_797),
.B(n_733),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_R g808 ( 
.A(n_802),
.B(n_166),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_801),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_805),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_804),
.Y(n_811)
);

BUFx12f_ASAP7_75t_L g812 ( 
.A(n_806),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_807),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_803),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_813),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_SL g816 ( 
.A1(n_809),
.A2(n_810),
.B1(n_814),
.B2(n_812),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_811),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_808),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_SL g819 ( 
.A1(n_809),
.A2(n_708),
.B1(n_723),
.B2(n_703),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_813),
.Y(n_820)
);

XNOR2x1_ASAP7_75t_L g821 ( 
.A(n_814),
.B(n_168),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_813),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_809),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_816),
.A2(n_689),
.B1(n_746),
.B2(n_752),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_815),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_820),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_823),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_822),
.Y(n_828)
);

AOI31xp33_ASAP7_75t_L g829 ( 
.A1(n_821),
.A2(n_723),
.A3(n_691),
.B(n_687),
.Y(n_829)
);

AO22x2_ASAP7_75t_L g830 ( 
.A1(n_817),
.A2(n_745),
.B1(n_757),
.B2(n_753),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_818),
.B(n_759),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_819),
.A2(n_703),
.B1(n_680),
.B2(n_689),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_827),
.B(n_689),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_825),
.A2(n_828),
.B1(n_826),
.B2(n_831),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_SL g835 ( 
.A1(n_824),
.A2(n_703),
.B1(n_680),
.B2(n_647),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_829),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_SL g837 ( 
.A1(n_832),
.A2(n_703),
.B1(n_680),
.B2(n_647),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_836),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_833),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_SL g840 ( 
.A1(n_838),
.A2(n_834),
.B1(n_835),
.B2(n_837),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_840),
.A2(n_839),
.B1(n_830),
.B2(n_703),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_700),
.B1(n_715),
.B2(n_705),
.C(n_699),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_842),
.A2(n_705),
.B1(n_736),
.B2(n_699),
.Y(n_843)
);


endmodule