module real_jpeg_25150_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_35),
.B1(n_68),
.B2(n_70),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_35),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_21),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_3),
.A2(n_25),
.B(n_94),
.C(n_241),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_22),
.B1(n_25),
.B2(n_181),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_3),
.B(n_57),
.C(n_73),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_3),
.A2(n_68),
.B1(n_70),
.B2(n_181),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_3),
.A2(n_54),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_136),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_37),
.B1(n_43),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_22),
.B1(n_25),
.B2(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_68),
.B1(n_70),
.B2(n_84),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_84),
.Y(n_201)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_7),
.A2(n_29),
.B1(n_43),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_7),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_7),
.A2(n_68),
.B1(n_70),
.B2(n_121),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_121),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_8),
.Y(n_94)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_10),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_68),
.B1(n_70),
.B2(n_88),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_22),
.B1(n_25),
.B2(n_88),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_88),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_42),
.B1(n_68),
.B2(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_11),
.A2(n_22),
.B1(n_25),
.B2(n_42),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_22),
.B1(n_25),
.B2(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_12),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_12),
.A2(n_68),
.B1(n_70),
.B2(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_43),
.B1(n_98),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_98),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_22),
.B1(n_25),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_13),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_13),
.A2(n_31),
.B1(n_43),
.B2(n_172),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_13),
.A2(n_68),
.B1(n_70),
.B2(n_172),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_172),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_15),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_22),
.B1(n_25),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_189)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_16),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_16),
.A2(n_55),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_16),
.Y(n_204)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_16),
.A2(n_55),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_34),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_27),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_21),
.A2(n_27),
.B1(n_120),
.B2(n_213),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_21),
.A2(n_27),
.B1(n_41),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_22),
.A2(n_25),
.B1(n_94),
.B2(n_95),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_22),
.A2(n_26),
.B(n_182),
.C(n_192),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_24),
.B(n_25),
.C(n_38),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_27),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_27),
.A2(n_124),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_30),
.B(n_181),
.Y(n_182)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_33),
.A2(n_83),
.B(n_85),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_33),
.B(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_83),
.B1(n_122),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_33),
.A2(n_122),
.B1(n_144),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_33),
.A2(n_85),
.B(n_212),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_36),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_40),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_40),
.B(n_357),
.Y(n_358)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_43),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_356),
.B(n_358),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_344),
.B(n_355),
.Y(n_47)
);

OAI31xp33_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_147),
.A3(n_161),
.B(n_341),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_125),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_50),
.B(n_125),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_89),
.C(n_105),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_51),
.A2(n_89),
.B1(n_90),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_51),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_79),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_53),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_53),
.A2(n_64),
.B1(n_65),
.B2(n_80),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_61),
.B(n_63),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_63),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_54),
.A2(n_188),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_54),
.A2(n_60),
.B1(n_110),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_54),
.A2(n_270),
.B(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_55),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_73),
.B2(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_56),
.B(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_61),
.B(n_181),
.Y(n_274)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_71),
.B1(n_78),
.B2(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_70),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_68),
.B(n_262),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_70),
.A2(n_95),
.B(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_78),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_71),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_71),
.A2(n_78),
.B1(n_236),
.B2(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_76),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_76),
.A2(n_101),
.B1(n_115),
.B2(n_176),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_76),
.B(n_181),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_76),
.A2(n_177),
.B(n_251),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_78),
.B(n_178),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_104),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_99),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_92),
.A2(n_93),
.B1(n_138),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_92),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_92),
.A2(n_210),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_93),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_93),
.A2(n_117),
.B(n_196),
.Y(n_320)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_101),
.A2(n_235),
.B(n_237),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_101),
.A2(n_237),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_105),
.A2(n_106),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.C(n_118),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_107),
.A2(n_108),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_109),
.Y(n_313)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_111),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_111),
.A2(n_244),
.B(n_268),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_116),
.B(n_118),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_143),
.B2(n_146),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_140),
.C(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_136),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_135),
.A2(n_136),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_136),
.B(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_140),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_140),
.B(n_154),
.C(n_158),
.Y(n_354)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_146),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_143),
.B(n_150),
.C(n_153),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_148),
.A2(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_160),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_149),
.B(n_160),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_155),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_159),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_334),
.B(n_340),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_324),
.B(n_333),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_222),
.B(n_307),
.C(n_323),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_205),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_165),
.B(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_183),
.C(n_193),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_166),
.A2(n_167),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_179),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_174),
.C(n_179),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_183),
.A2(n_184),
.B1(n_193),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_190),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_193),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_200),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_214),
.B1(n_215),
.B2(n_221),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g360 ( 
.A(n_206),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.CI(n_211),
.CON(n_206),
.SN(n_206)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_216),
.B(n_220),
.C(n_221),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_217),
.B(n_219),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_300),
.B(n_306),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_255),
.B(n_299),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_247),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_227),
.B(n_247),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_246),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_234),
.C(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.C(n_252),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_252),
.B1(n_253),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_293),
.B(n_298),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_283),
.B(n_292),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_271),
.B(n_282),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_278),
.B(n_281),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_291),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.C(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_322),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_322),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_312),
.C(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_319),
.C(n_321),
.Y(n_332)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_326),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.C(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_346),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_350),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_357)
);


endmodule