module fake_jpeg_26841_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_265;
wire n_115;
wire n_123;
wire n_192;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_20),
.B1(n_32),
.B2(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_50),
.B1(n_53),
.B2(n_42),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_34),
.B2(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_33),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_37),
.B1(n_41),
.B2(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g115 ( 
.A(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_65),
.B(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_72),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_40),
.C(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_26),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_76),
.B1(n_16),
.B2(n_40),
.Y(n_110)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_37),
.B(n_41),
.C(n_39),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_31),
.B(n_17),
.C(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_16),
.B1(n_30),
.B2(n_22),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_93),
.B1(n_40),
.B2(n_39),
.Y(n_104)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_97),
.B1(n_62),
.B2(n_40),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_90),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_31),
.B1(n_23),
.B2(n_18),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_33),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_35),
.B(n_25),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_117),
.B1(n_81),
.B2(n_75),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_0),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_86),
.B(n_67),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_63),
.Y(n_116)
);

AOI22x1_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_35),
.B1(n_30),
.B2(n_22),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_35),
.B1(n_22),
.B2(n_2),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_77),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_35),
.B1(n_1),
.B2(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_131),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_129),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_139),
.B1(n_151),
.B2(n_11),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_88),
.B1(n_74),
.B2(n_63),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_146),
.B1(n_152),
.B2(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_113),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_147),
.B(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_79),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_98),
.C(n_97),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_150),
.C(n_157),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_111),
.B(n_102),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_115),
.B(n_82),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_66),
.B1(n_90),
.B2(n_96),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_92),
.C(n_67),
.Y(n_150)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_110),
.B1(n_111),
.B2(n_106),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_95),
.B1(n_87),
.B2(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_64),
.C(n_85),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_126),
.B(n_107),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_158),
.A2(n_163),
.B(n_174),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_11),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_161),
.C(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_133),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_115),
.B1(n_105),
.B2(n_118),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_169),
.B1(n_174),
.B2(n_185),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_0),
.B(n_5),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_11),
.C(n_6),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_0),
.B(n_6),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_148),
.B(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_131),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_6),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_134),
.C(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

OA21x2_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_201),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_147),
.C(n_152),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_161),
.C(n_184),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_140),
.B(n_8),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_7),
.B(n_10),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_168),
.B1(n_185),
.B2(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_15),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_171),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_15),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_178),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

AOI31xp33_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_162),
.A3(n_188),
.B(n_160),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_232),
.C(n_196),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_170),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_191),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_163),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_166),
.C(n_176),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_172),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_210),
.B(n_231),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_209),
.B(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_205),
.B(n_190),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_240),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_207),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_243),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_209),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_230),
.C(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_193),
.C(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_249),
.C(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_211),
.C(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_190),
.B(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_256),
.C(n_263),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_203),
.B1(n_219),
.B2(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_222),
.B1(n_206),
.B2(n_181),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_226),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_228),
.C(n_207),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_237),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_248),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_192),
.B1(n_251),
.B2(n_240),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_192),
.B1(n_176),
.B2(n_183),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_247),
.B1(n_215),
.B2(n_235),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_208),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_7),
.Y(n_285)
);

XNOR2x2_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_199),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_213),
.B(n_182),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_259),
.B(n_238),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_248),
.C(n_192),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_285),
.C(n_277),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_276),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_13),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_267),
.B(n_273),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_291),
.C(n_281),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_12),
.C(n_13),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_280),
.A3(n_282),
.B1(n_278),
.B2(n_15),
.C1(n_14),
.C2(n_12),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_295),
.CI(n_289),
.CON(n_297),
.SN(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_293),
.C(n_288),
.Y(n_298)
);

OAI31xp33_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_297),
.A3(n_296),
.B(n_13),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);


endmodule