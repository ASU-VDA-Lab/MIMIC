module fake_jpeg_17330_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_32),
.B1(n_13),
.B2(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_33),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_1),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_21),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_22),
.B(n_24),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_58),
.B(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_62),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_60),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_25),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.C(n_77),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_50),
.B1(n_56),
.B2(n_49),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_53),
.C(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_53),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_52),
.B(n_51),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_75),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_90),
.CI(n_71),
.CON(n_98),
.SN(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_90),
.C(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_71),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_76),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_70),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_94),
.B1(n_83),
.B2(n_95),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_69),
.B1(n_82),
.B2(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_93),
.C(n_92),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_92),
.C(n_96),
.Y(n_103)
);

XOR2x2_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_94),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_104),
.B(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.C(n_105),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_104),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_109),
.Y(n_112)
);


endmodule