module fake_jpeg_11351_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_46),
.B1(n_25),
.B2(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_17),
.B1(n_29),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_68),
.B1(n_39),
.B2(n_38),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_69),
.B1(n_23),
.B2(n_20),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_73),
.Y(n_80)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_17),
.B1(n_29),
.B2(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_28),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_39),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_42),
.B(n_40),
.C(n_43),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_77),
.A2(n_21),
.B(n_19),
.C(n_35),
.D(n_27),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_128)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_107),
.B1(n_61),
.B2(n_48),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_104),
.Y(n_130)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_99),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_18),
.B1(n_32),
.B2(n_26),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_18),
.B1(n_32),
.B2(n_26),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_24),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_37),
.C(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_26),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_19),
.B(n_35),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_108),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_21),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_82),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_84),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_121),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_53),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_102),
.C(n_33),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_102),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_76),
.A3(n_100),
.B1(n_98),
.B2(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_132),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_93),
.B1(n_86),
.B2(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_13),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_105),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_30),
.B(n_21),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_142),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_72),
.B1(n_71),
.B2(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_158),
.B1(n_162),
.B2(n_172),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_154),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_147),
.A2(n_159),
.B(n_163),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_92),
.B1(n_91),
.B2(n_83),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_155),
.B1(n_4),
.B2(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_92),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_157),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_81),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_83),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_134),
.B1(n_111),
.B2(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_116),
.B1(n_125),
.B2(n_139),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_135),
.B1(n_133),
.B2(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_95),
.B1(n_30),
.B2(n_35),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_19),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_166),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_0),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_15),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_0),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_3),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_14),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_3),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_13),
.C(n_12),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_11),
.C(n_10),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_119),
.B1(n_115),
.B2(n_112),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_185),
.B1(n_190),
.B2(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_150),
.B1(n_149),
.B2(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_184),
.B1(n_187),
.B2(n_199),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_114),
.B1(n_119),
.B2(n_11),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_186),
.B(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

AOI22x1_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_206),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_4),
.C(n_6),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_174),
.C(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_142),
.A2(n_171),
.B1(n_144),
.B2(n_155),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_216),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_154),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_225),
.Y(n_239)
);

AOI221xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.C(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_177),
.A2(n_172),
.B1(n_173),
.B2(n_168),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_184),
.B1(n_192),
.B2(n_178),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_168),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_230),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_170),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_143),
.C(n_163),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_197),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_6),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_234),
.C(n_186),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_7),
.C(n_8),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_242),
.C(n_259),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_218),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_177),
.B1(n_193),
.B2(n_175),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_243),
.B1(n_249),
.B2(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_175),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_217),
.B1(n_233),
.B2(n_228),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_250),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_252),
.B1(n_222),
.B2(n_224),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_220),
.B1(n_179),
.B2(n_213),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_200),
.B1(n_187),
.B2(n_192),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_214),
.A2(n_185),
.B1(n_200),
.B2(n_176),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_203),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_256),
.B1(n_243),
.B2(n_257),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_232),
.C(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_235),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_219),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_218),
.B1(n_226),
.B2(n_236),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_251),
.B1(n_260),
.B2(n_253),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_188),
.C(n_190),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_7),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_8),
.C(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_250),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_252),
.B1(n_248),
.B2(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_280),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_272),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_268),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_291),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_278),
.B1(n_296),
.B2(n_290),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_273),
.B1(n_279),
.B2(n_265),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_257),
.B(n_9),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_9),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_267),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_300),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_264),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_266),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_264),
.B(n_276),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_308),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_281),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_310),
.B(n_314),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_301),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_291),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_298),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_323),
.B(n_326),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_293),
.C(n_302),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_316),
.C(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_329),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_283),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_302),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_328),
.B(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.B(n_312),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_326),
.B1(n_325),
.B2(n_295),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_312),
.B(n_297),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_297),
.Y(n_337)
);


endmodule