module fake_netlist_5_2111_n_2267 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_239, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2267);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_239;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2267;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_99),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_42),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_83),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_108),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_35),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_161),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_242),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_182),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_81),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_117),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_65),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_121),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_212),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_112),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_109),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_58),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_227),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_167),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_61),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_32),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_87),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_135),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_92),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_170),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_210),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_177),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_183),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_14),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_190),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_78),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_111),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_133),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_77),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_153),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_175),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_96),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_71),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_36),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_188),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_42),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_39),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_28),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_164),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_75),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_16),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_69),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_181),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_132),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_69),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_192),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_186),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_180),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_94),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_30),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_101),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_138),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_88),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_62),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_146),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_220),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_34),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_15),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_152),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_201),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_115),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_233),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_124),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_122),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_6),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_19),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_20),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_230),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_171),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_79),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_149),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_140),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_57),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_98),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_113),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_34),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_72),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_5),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_67),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_13),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_159),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_200),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_3),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_125),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_75),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_63),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_216),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_14),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_179),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_102),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_126),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_119),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_151),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_107),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_39),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_222),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_53),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_2),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_62),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_97),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_231),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_218),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_43),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_23),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_27),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_44),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_189),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_178),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_4),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_50),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_187),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_221),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_73),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_54),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_185),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_11),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_6),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_241),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_214),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_147),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_46),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_49),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_81),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_40),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_137),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_128),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_106),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_33),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_217),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_142),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_56),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_15),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_25),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_228),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_168),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_19),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_203),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_83),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_105),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_55),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_26),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_65),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_51),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_93),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_155),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_160),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_224),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_197),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_165),
.Y(n_437)
);

BUFx2_ASAP7_75t_SL g438 ( 
.A(n_130),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_154),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_174),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_194),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_176),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_55),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_29),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_2),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_7),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_129),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_193),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_116),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_157),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_232),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_148),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_90),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_45),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_48),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_236),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_50),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_91),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_11),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_61),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_52),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_66),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_240),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_25),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_208),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_225),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_38),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_40),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_60),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_80),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_32),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_0),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_79),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_27),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_243),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_258),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_258),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_340),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_262),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_248),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_252),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_295),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_384),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_310),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_328),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_254),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_295),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_295),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_295),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_295),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_340),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_295),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_360),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_358),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_445),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_437),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_445),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_256),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_257),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_244),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_263),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_468),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_266),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_249),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_273),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_303),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_468),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_249),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_265),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_278),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_365),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_278),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_311),
.Y(n_532)
);

INVxp33_ASAP7_75t_SL g533 ( 
.A(n_245),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_389),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_311),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_378),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_339),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_267),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_365),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_268),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_303),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_411),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_463),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_270),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_266),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_339),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_367),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_367),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_365),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_378),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_454),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_272),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_412),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_273),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_279),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_389),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_387),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_282),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_389),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_285),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_387),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_299),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_329),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_299),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_315),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_315),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_320),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_320),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_324),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_276),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_286),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_324),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_352),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_352),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_287),
.Y(n_579)
);

INVxp33_ASAP7_75t_SL g580 ( 
.A(n_251),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_355),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_288),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_276),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_290),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_355),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_361),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_294),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_361),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_365),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_365),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_363),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_305),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_275),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_365),
.Y(n_595)
);

BUFx2_ASAP7_75t_SL g596 ( 
.A(n_259),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_363),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_381),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_381),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_308),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_318),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_325),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_473),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_395),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_284),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_247),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_323),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_323),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_484),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_482),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_584),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_497),
.Y(n_615)
);

OA21x2_ASAP7_75t_L g616 ( 
.A1(n_498),
.A2(n_250),
.B(n_247),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_500),
.Y(n_617)
);

INVx6_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_483),
.B(n_323),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_493),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_511),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_559),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_498),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_560),
.B(n_412),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_496),
.A2(n_274),
.B(n_246),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_480),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_559),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_514),
.B(n_259),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_513),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_496),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_499),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_502),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_505),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_505),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_506),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_506),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_606),
.B(n_322),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_508),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_508),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_509),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_509),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_533),
.B(n_322),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_479),
.B(n_436),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_485),
.B(n_255),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_510),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_519),
.A2(n_321),
.B1(n_460),
.B2(n_331),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_512),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_479),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_567),
.B(n_403),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_512),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_526),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_481),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_523),
.A2(n_261),
.B1(n_269),
.B2(n_260),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_538),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_515),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_517),
.B(n_246),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_517),
.B(n_274),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_541),
.A2(n_556),
.B1(n_477),
.B2(n_495),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_520),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_521),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_540),
.B(n_544),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_555),
.B(n_313),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_558),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_521),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_524),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_524),
.Y(n_676)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_527),
.B(n_438),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_545),
.B(n_436),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_527),
.Y(n_679)
);

AND3x2_ASAP7_75t_L g680 ( 
.A(n_495),
.B(n_332),
.C(n_313),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_562),
.B(n_332),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_566),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_594),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_481),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_564),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_486),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_486),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_487),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_487),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_489),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_566),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_575),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_489),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_534),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_560),
.B(n_280),
.Y(n_695)
);

CKINVDCx6p67_ASAP7_75t_R g696 ( 
.A(n_603),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_563),
.B(n_280),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_568),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_490),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_490),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_492),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_568),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_570),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_570),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_371),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_684),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_672),
.B(n_583),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_678),
.B(n_585),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_619),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_607),
.B(n_580),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_620),
.B(n_588),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_678),
.B(n_593),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_619),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_612),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_684),
.Y(n_716)
);

INVxp33_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_678),
.B(n_600),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_632),
.B(n_601),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_625),
.A2(n_596),
.B1(n_476),
.B2(n_289),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_635),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_R g722 ( 
.A(n_621),
.B(n_602),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_695),
.B(n_478),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_684),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_649),
.B(n_574),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_662),
.B(n_605),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_686),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_686),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_695),
.B(n_501),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_689),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_635),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_657),
.A2(n_370),
.B1(n_391),
.B2(n_317),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_622),
.B(n_634),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_681),
.B(n_525),
.Y(n_734)
);

INVxp33_ASAP7_75t_SL g735 ( 
.A(n_660),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_677),
.B(n_436),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_668),
.A2(n_536),
.B1(n_561),
.B2(n_551),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_SL g738 ( 
.A(n_638),
.B(n_565),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_629),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_SL g740 ( 
.A1(n_705),
.A2(n_503),
.B1(n_253),
.B2(n_264),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_689),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_689),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_696),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_610),
.B(n_656),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_625),
.A2(n_289),
.B1(n_359),
.B2(n_271),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_671),
.B(n_596),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_658),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_627),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_658),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_617),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_624),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_690),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_492),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_624),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_690),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_610),
.B(n_494),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_650),
.B(n_436),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_690),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_627),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_614),
.B(n_534),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_501),
.Y(n_764)
);

OAI21xp33_ASAP7_75t_SL g765 ( 
.A1(n_626),
.A2(n_359),
.B(n_271),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_687),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_663),
.B(n_403),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_645),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_616),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_645),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_673),
.B(n_403),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_627),
.B(n_531),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_685),
.B(n_531),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_645),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_638),
.B(n_438),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_647),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_610),
.B(n_494),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_696),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_658),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_692),
.Y(n_783)
);

BUFx6f_ASAP7_75t_SL g784 ( 
.A(n_644),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_694),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_693),
.Y(n_786)
);

INVx6_ASAP7_75t_L g787 ( 
.A(n_686),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_697),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_647),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_686),
.Y(n_790)
);

BUFx8_ASAP7_75t_SL g791 ( 
.A(n_683),
.Y(n_791)
);

AND3x1_ASAP7_75t_L g792 ( 
.A(n_654),
.B(n_399),
.C(n_395),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_656),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_656),
.B(n_661),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_694),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_647),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_656),
.B(n_542),
.Y(n_797)
);

INVxp33_ASAP7_75t_L g798 ( 
.A(n_654),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_658),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_694),
.B(n_403),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_699),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_658),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_644),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_694),
.B(n_440),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_652),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_644),
.B(n_440),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_686),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_651),
.B(n_542),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_650),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_699),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_644),
.B(n_543),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_658),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_688),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_677),
.A2(n_488),
.B1(n_504),
.B2(n_491),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_659),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_680),
.Y(n_816)
);

INVxp33_ASAP7_75t_L g817 ( 
.A(n_683),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_616),
.A2(n_399),
.B1(n_427),
.B2(n_408),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_682),
.B(n_440),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_700),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_682),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_691),
.A2(n_443),
.B1(n_423),
.B2(n_557),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_700),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_616),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_650),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_665),
.A2(n_507),
.B1(n_333),
.B2(n_330),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_661),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_688),
.B(n_581),
.Y(n_831)
);

BUFx4f_ASAP7_75t_L g832 ( 
.A(n_616),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_652),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_650),
.B(n_436),
.Y(n_834)
);

BUFx4f_ASAP7_75t_L g835 ( 
.A(n_688),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_698),
.B(n_563),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_698),
.B(n_522),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_613),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_688),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_659),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_569),
.C(n_283),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_613),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_702),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_615),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_688),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

XOR2xp5_ASAP7_75t_L g847 ( 
.A(n_703),
.B(n_281),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_615),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_628),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_626),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_659),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_250),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_703),
.B(n_440),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_628),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_688),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_701),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_636),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_704),
.B(n_292),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_636),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_701),
.B(n_326),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_637),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_665),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_659),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_637),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_704),
.B(n_336),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_665),
.B(n_337),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_666),
.B(n_341),
.Y(n_867)
);

BUFx8_ASAP7_75t_SL g868 ( 
.A(n_666),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_664),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_609),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_821),
.B(n_342),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_843),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_862),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_701),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_719),
.B(n_701),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_772),
.A2(n_666),
.B(n_410),
.C(n_417),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_818),
.A2(n_427),
.B1(n_429),
.B2(n_408),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_723),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_772),
.B(n_701),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_SL g881 ( 
.A(n_828),
.B(n_725),
.C(n_726),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_748),
.B(n_701),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_772),
.A2(n_455),
.B1(n_459),
.B2(n_429),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_803),
.B(n_666),
.Y(n_884)
);

OAI22xp33_ASAP7_75t_L g885 ( 
.A1(n_798),
.A2(n_459),
.B1(n_461),
.B2(n_455),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_803),
.B(n_639),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_832),
.B(n_365),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_788),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_708),
.A2(n_467),
.B(n_474),
.C(n_461),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_788),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_832),
.B(n_365),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_710),
.B(n_293),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_712),
.A2(n_474),
.B(n_467),
.C(n_639),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_797),
.B(n_640),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_707),
.B(n_641),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_842),
.B(n_641),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_718),
.A2(n_410),
.B1(n_417),
.B2(n_371),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_734),
.A2(n_344),
.B1(n_349),
.B2(n_343),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_793),
.Y(n_899)
);

BUFx10_ASAP7_75t_L g900 ( 
.A(n_776),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_832),
.A2(n_264),
.B1(n_277),
.B2(n_253),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_842),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_732),
.A2(n_390),
.B1(n_420),
.B2(n_419),
.C(n_425),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_848),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_756),
.B(n_365),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_848),
.B(n_642),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_849),
.B(n_642),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_859),
.B(n_643),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_859),
.B(n_643),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_821),
.B(n_726),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_759),
.B(n_453),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_811),
.B(n_646),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_784),
.A2(n_351),
.B1(n_353),
.B2(n_350),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_769),
.B(n_297),
.C(n_296),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_762),
.B(n_354),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_837),
.A2(n_572),
.B(n_571),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_808),
.B(n_300),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_780),
.B(n_646),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_746),
.B(n_453),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_721),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_793),
.B(n_648),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_723),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_831),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_731),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_762),
.B(n_648),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_729),
.B(n_571),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_731),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_862),
.B(n_356),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_741),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_751),
.B(n_729),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_784),
.A2(n_366),
.B1(n_368),
.B2(n_357),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_764),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_763),
.B(n_301),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_741),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_764),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_745),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_838),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_838),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_829),
.B(n_653),
.Y(n_940)
);

AND2x2_ASAP7_75t_SL g941 ( 
.A(n_792),
.B(n_277),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_722),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_763),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_825),
.A2(n_298),
.B1(n_302),
.B2(n_291),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_829),
.B(n_653),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_830),
.B(n_655),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_825),
.A2(n_747),
.B1(n_850),
.B2(n_852),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_L g948 ( 
.A(n_736),
.B(n_373),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_717),
.B(n_572),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_844),
.Y(n_950)
);

BUFx6f_ASAP7_75t_SL g951 ( 
.A(n_714),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_747),
.A2(n_298),
.B1(n_302),
.B2(n_291),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_720),
.B(n_306),
.C(n_304),
.Y(n_953)
);

INVxp33_ASAP7_75t_L g954 ( 
.A(n_847),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_814),
.B(n_609),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_844),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_745),
.Y(n_957)
);

OAI221xp5_ASAP7_75t_L g958 ( 
.A1(n_836),
.A2(n_441),
.B1(n_307),
.B2(n_327),
.C(n_334),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_SL g959 ( 
.A(n_735),
.B(n_374),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_736),
.B(n_376),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_862),
.B(n_377),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_795),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_850),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_751),
.B(n_309),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_854),
.Y(n_965)
);

BUFx8_ASAP7_75t_L g966 ( 
.A(n_795),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_715),
.B(n_380),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_847),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_830),
.B(n_655),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_794),
.B(n_667),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_854),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_857),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_852),
.B(n_855),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_857),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_852),
.B(n_667),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_861),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_715),
.B(n_383),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_715),
.B(n_809),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_L g979 ( 
.A1(n_737),
.A2(n_327),
.B1(n_334),
.B2(n_307),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_767),
.B(n_669),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_861),
.B(n_864),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_864),
.B(n_669),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_870),
.B(n_774),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_766),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_817),
.B(n_573),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_806),
.B(n_573),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_766),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_870),
.B(n_312),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_768),
.B(n_674),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_768),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_715),
.B(n_385),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_750),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_786),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_SL g994 ( 
.A(n_800),
.B(n_316),
.C(n_314),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_740),
.A2(n_765),
.B(n_834),
.C(n_760),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_786),
.B(n_676),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_787),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_801),
.B(n_676),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_750),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_801),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_736),
.B(n_386),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_784),
.A2(n_392),
.B1(n_393),
.B2(n_396),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_810),
.B(n_679),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_739),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_820),
.B(n_824),
.Y(n_1005)
);

INVx8_ASAP7_75t_L g1006 ( 
.A(n_778),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_822),
.A2(n_379),
.B1(n_382),
.B2(n_446),
.C(n_444),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_820),
.B(n_611),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_816),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_824),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_715),
.B(n_404),
.Y(n_1011)
);

AND2x6_ASAP7_75t_SL g1012 ( 
.A(n_778),
.B(n_576),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_809),
.B(n_827),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_809),
.B(n_827),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_775),
.B(n_858),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_714),
.B(n_576),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_753),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_809),
.B(n_405),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_754),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_860),
.A2(n_633),
.B(n_631),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_714),
.B(n_577),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_809),
.B(n_416),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_845),
.B(n_611),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_753),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_865),
.B(n_319),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_841),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_709),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_783),
.B(n_733),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_706),
.B(n_623),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_739),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_709),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_783),
.B(n_577),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_835),
.A2(n_633),
.B(n_631),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_827),
.B(n_422),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_827),
.B(n_706),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_866),
.A2(n_631),
.B(n_633),
.C(n_397),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_747),
.A2(n_345),
.B1(n_452),
.B2(n_441),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_867),
.A2(n_442),
.B1(n_424),
.B2(n_426),
.Y(n_1038)
);

AND2x6_ASAP7_75t_L g1039 ( 
.A(n_716),
.B(n_345),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_L g1040 ( 
.A(n_901),
.B(n_827),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_931),
.B(n_778),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_938),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_L g1043 ( 
.A(n_901),
.B(n_736),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_939),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_942),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_875),
.B(n_735),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_950),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_956),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_875),
.B(n_963),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1015),
.B(n_716),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_931),
.B(n_778),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_892),
.A2(n_804),
.B1(n_853),
.B2(n_819),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_895),
.B(n_724),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_SL g1054 ( 
.A1(n_968),
.A2(n_781),
.B1(n_744),
.B2(n_785),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_883),
.A2(n_747),
.B1(n_397),
.B2(n_400),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_1004),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_879),
.Y(n_1058)
);

CKINVDCx6p67_ASAP7_75t_R g1059 ( 
.A(n_951),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_892),
.A2(n_736),
.B1(n_787),
.B2(n_730),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_918),
.B(n_911),
.C(n_903),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_971),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_881),
.A2(n_736),
.B1(n_787),
.B2(n_730),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_899),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_873),
.B(n_727),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_972),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_963),
.B(n_783),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_974),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_899),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_918),
.B(n_724),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_911),
.B(n_785),
.C(n_781),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_899),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_949),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_902),
.B(n_904),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_742),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_899),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_963),
.B(n_835),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_985),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_951),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_1016),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_L g1082 ( 
.A(n_983),
.B(n_744),
.C(n_400),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_963),
.Y(n_1083)
);

BUFx4f_ASAP7_75t_L g1084 ( 
.A(n_1006),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_923),
.B(n_375),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_874),
.B(n_835),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_888),
.B(n_375),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_944),
.B(n_742),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_883),
.A2(n_944),
.B1(n_877),
.B2(n_952),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1021),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_927),
.B(n_743),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1032),
.B(n_727),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_873),
.B(n_880),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_976),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_984),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_1030),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_913),
.B(n_755),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_987),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_997),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_934),
.B(n_738),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1025),
.A2(n_421),
.B(n_415),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1027),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_947),
.B(n_727),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_990),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_924),
.B(n_755),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_993),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_933),
.B(n_758),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1000),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_943),
.B(n_868),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1031),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_880),
.B(n_728),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_994),
.B(n_757),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_872),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_890),
.B(n_816),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1010),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_936),
.B(n_988),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_934),
.B(n_816),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1019),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_886),
.B(n_758),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_997),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_986),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1005),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_981),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_1006),
.B(n_791),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_975),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_922),
.Y(n_1126)
);

BUFx8_ASAP7_75t_L g1127 ( 
.A(n_1028),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_947),
.B(n_728),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_896),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_882),
.B(n_728),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_926),
.B(n_761),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_954),
.A2(n_338),
.B1(n_346),
.B2(n_335),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_997),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_997),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_878),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_1006),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_906),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_973),
.Y(n_1138)
);

AND2x6_ASAP7_75t_SL g1139 ( 
.A(n_988),
.B(n_578),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_962),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_966),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_1012),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_921),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_925),
.Y(n_1144)
);

NOR2x2_ASAP7_75t_L g1145 ( 
.A(n_979),
.B(n_757),
.Y(n_1145)
);

NAND2x1p5_ASAP7_75t_L g1146 ( 
.A(n_1035),
.B(n_770),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1026),
.B(n_770),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_955),
.A2(n_961),
.B1(n_929),
.B2(n_1025),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_928),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_966),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_887),
.B(n_770),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_983),
.A2(n_413),
.B1(n_348),
.B2(n_362),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1039),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_877),
.A2(n_415),
.B1(n_452),
.B2(n_439),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_930),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_900),
.B(n_761),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_959),
.B(n_431),
.Y(n_1158)
);

CKINVDCx6p67_ASAP7_75t_R g1159 ( 
.A(n_900),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_919),
.B(n_749),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_908),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_941),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_909),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1037),
.A2(n_434),
.B1(n_439),
.B2(n_458),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_887),
.B(n_790),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_935),
.Y(n_1166)
);

BUFx4f_ASAP7_75t_L g1167 ( 
.A(n_941),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_937),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_891),
.B(n_790),
.Y(n_1169)
);

AND3x1_ASAP7_75t_L g1170 ( 
.A(n_1007),
.B(n_582),
.C(n_578),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1039),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_916),
.B(n_432),
.Y(n_1172)
);

AND2x6_ASAP7_75t_SL g1173 ( 
.A(n_964),
.B(n_582),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_957),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_884),
.B(n_749),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_1039),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_910),
.B(n_752),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_929),
.B(n_435),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_894),
.B(n_752),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_992),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_1039),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_982),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_891),
.A2(n_713),
.B(n_771),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_999),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1008),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1037),
.A2(n_435),
.B1(n_834),
.B2(n_760),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_961),
.A2(n_787),
.B1(n_790),
.B2(n_856),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_964),
.A2(n_807),
.B1(n_813),
.B2(n_856),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1017),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1024),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_989),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1039),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_970),
.B(n_782),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_885),
.A2(n_713),
.B1(n_833),
.B2(n_826),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1035),
.B(n_807),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_979),
.B(n_807),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1020),
.A2(n_876),
.B(n_1033),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_940),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_885),
.A2(n_789),
.B1(n_833),
.B2(n_826),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_945),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_871),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_953),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_779),
.B1(n_805),
.B2(n_796),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_978),
.B(n_813),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_946),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_980),
.B(n_996),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_969),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_998),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_898),
.B(n_586),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_978),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1003),
.B(n_782),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_917),
.B(n_586),
.Y(n_1212)
);

INVxp67_ASAP7_75t_SL g1213 ( 
.A(n_1029),
.Y(n_1213)
);

AO22x1_ASAP7_75t_L g1214 ( 
.A1(n_915),
.A2(n_364),
.B1(n_369),
.B2(n_372),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_920),
.A2(n_839),
.B1(n_813),
.B2(n_856),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_897),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_889),
.B(n_839),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_SL g1218 ( 
.A1(n_948),
.A2(n_347),
.B1(n_388),
.B2(n_394),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_995),
.B(n_893),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1023),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_920),
.B(n_799),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_912),
.A2(n_839),
.B1(n_863),
.B2(n_851),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1036),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_905),
.Y(n_1224)
);

BUFx8_ASAP7_75t_SL g1225 ( 
.A(n_914),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_SL g1226 ( 
.A(n_932),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1013),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_912),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1061),
.B(n_1002),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1040),
.A2(n_1014),
.B(n_1013),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1101),
.A2(n_905),
.B(n_960),
.C(n_1001),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1129),
.B(n_1038),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1056),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1116),
.A2(n_1034),
.B(n_1022),
.C(n_1018),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1081),
.B(n_1117),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_L g1236 ( 
.A(n_1069),
.B(n_1034),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1167),
.B(n_967),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1090),
.A2(n_398),
.B1(n_472),
.B2(n_470),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1046),
.A2(n_1022),
.B(n_1018),
.C(n_967),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1046),
.A2(n_977),
.B(n_1011),
.C(n_991),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1040),
.A2(n_1014),
.B(n_991),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1043),
.A2(n_1011),
.B(n_977),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1162),
.B(n_401),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1089),
.A2(n_402),
.B1(n_406),
.B2(n_407),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1045),
.B(n_433),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1183),
.A2(n_1197),
.B(n_1221),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1137),
.B(n_771),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1086),
.A2(n_777),
.B(n_773),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1161),
.B(n_773),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1095),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1163),
.B(n_777),
.Y(n_1251)
);

BUFx4f_ASAP7_75t_L g1252 ( 
.A(n_1070),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1122),
.B(n_779),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1167),
.B(n_447),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1098),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1191),
.B(n_789),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_R g1257 ( 
.A(n_1045),
.B(n_448),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1125),
.B(n_796),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1202),
.A2(n_589),
.B(n_592),
.C(n_587),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_R g1260 ( 
.A(n_1072),
.B(n_449),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1216),
.A2(n_589),
.B(n_592),
.C(n_587),
.Y(n_1261)
);

CKINVDCx6p67_ASAP7_75t_R g1262 ( 
.A(n_1070),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1185),
.B(n_805),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1209),
.A2(n_597),
.B(n_598),
.C(n_599),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_L g1265 ( 
.A(n_1089),
.B(n_450),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1135),
.Y(n_1266)
);

AND2x6_ASAP7_75t_L g1267 ( 
.A(n_1192),
.B(n_799),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1136),
.B(n_597),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1104),
.Y(n_1269)
);

NOR3xp33_ASAP7_75t_L g1270 ( 
.A(n_1100),
.B(n_414),
.C(n_409),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1136),
.B(n_451),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1052),
.B(n_456),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1148),
.A2(n_869),
.B(n_863),
.C(n_851),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1074),
.B(n_428),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1079),
.B(n_598),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1096),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1106),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1219),
.A2(n_599),
.B(n_604),
.C(n_530),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1135),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1178),
.A2(n_466),
.B1(n_465),
.B2(n_851),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1113),
.Y(n_1281)
);

AO22x1_ASAP7_75t_L g1282 ( 
.A1(n_1082),
.A2(n_430),
.B1(n_457),
.B2(n_462),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1064),
.B(n_799),
.Y(n_1283)
);

NAND2x1_ASAP7_75t_SL g1284 ( 
.A(n_1041),
.B(n_604),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1069),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_SL g1286 ( 
.A(n_1084),
.B(n_1154),
.Y(n_1286)
);

AO32x1_ASAP7_75t_L g1287 ( 
.A1(n_1047),
.A2(n_528),
.A3(n_554),
.B1(n_530),
.B2(n_532),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1164),
.A2(n_464),
.B1(n_469),
.B2(n_528),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1164),
.A2(n_535),
.B1(n_553),
.B2(n_552),
.Y(n_1289)
);

NOR3xp33_ASAP7_75t_L g1290 ( 
.A(n_1153),
.B(n_554),
.C(n_532),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1108),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1143),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1155),
.A2(n_535),
.B1(n_552),
.B2(n_549),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1201),
.B(n_802),
.Y(n_1294)
);

OR2x6_ASAP7_75t_SL g1295 ( 
.A(n_1080),
.B(n_537),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1043),
.A2(n_869),
.B(n_863),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1049),
.A2(n_869),
.B(n_846),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1155),
.A2(n_1055),
.B1(n_1186),
.B2(n_1196),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1056),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1182),
.B(n_802),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1115),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1121),
.B(n_802),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_SL g1303 ( 
.A(n_1158),
.B(n_549),
.C(n_537),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1118),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1138),
.B(n_812),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1208),
.B(n_812),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1055),
.A2(n_553),
.B1(n_548),
.B2(n_547),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1196),
.A2(n_846),
.B1(n_840),
.B2(n_823),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1099),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1058),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1041),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1118),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1178),
.A2(n_840),
.B(n_823),
.C(n_815),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1178),
.A2(n_823),
.B(n_815),
.C(n_812),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1186),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1219),
.A2(n_529),
.B(n_539),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1157),
.B(n_815),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1157),
.B(n_0),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1041),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1050),
.A2(n_546),
.B1(n_539),
.B2(n_591),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1099),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1051),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1218),
.B(n_550),
.C(n_590),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1114),
.B(n_1),
.Y(n_1324)
);

OAI22x1_ASAP7_75t_L g1325 ( 
.A1(n_1114),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1130),
.A2(n_1086),
.B(n_1152),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1138),
.B(n_664),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_L g1328 ( 
.A1(n_1217),
.A2(n_595),
.B(n_630),
.C(n_623),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_L g1329 ( 
.A1(n_1217),
.A2(n_630),
.B(n_623),
.C(n_237),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1138),
.B(n_664),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1165),
.A2(n_1169),
.B(n_1206),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1075),
.A2(n_9),
.B(n_17),
.C(n_18),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1143),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1126),
.B(n_17),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1208),
.B(n_1200),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1088),
.A2(n_618),
.B1(n_670),
.B2(n_664),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1165),
.A2(n_675),
.B(n_670),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1169),
.A2(n_675),
.B(n_670),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1099),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1200),
.A2(n_618),
.B1(n_670),
.B2(n_664),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1138),
.B(n_1198),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1224),
.A2(n_675),
.B(n_20),
.C(n_21),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1205),
.B(n_650),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_SL g1344 ( 
.A(n_1176),
.B(n_618),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1123),
.A2(n_675),
.B(n_21),
.C(n_22),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1151),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1087),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1149),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1205),
.B(n_675),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1085),
.B(n_1132),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_SL g1351 ( 
.A(n_1176),
.B(n_675),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1071),
.A2(n_618),
.B(n_235),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1198),
.B(n_18),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1124),
.B(n_100),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1207),
.B(n_24),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1099),
.Y(n_1356)
);

INVx8_ASAP7_75t_L g1357 ( 
.A(n_1151),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1051),
.B(n_103),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1085),
.B(n_24),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1051),
.B(n_223),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1207),
.B(n_215),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1220),
.B(n_26),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1092),
.A2(n_1112),
.B1(n_1226),
.B2(n_1067),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1173),
.B(n_28),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1176),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1078),
.A2(n_211),
.B(n_209),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1220),
.B(n_31),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1228),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1078),
.A2(n_206),
.B(n_205),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1149),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1156),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1092),
.A2(n_204),
.B1(n_202),
.B2(n_199),
.Y(n_1372)
);

AND2x2_ASAP7_75t_SL g1373 ( 
.A(n_1084),
.B(n_38),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1087),
.B(n_198),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1193),
.A2(n_195),
.B(n_184),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1091),
.A2(n_173),
.B(n_169),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1156),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1067),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1053),
.A2(n_166),
.B(n_163),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1073),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1103),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1107),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1127),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1127),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1213),
.A2(n_158),
.B(n_156),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1059),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1175),
.A2(n_150),
.B(n_145),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1047),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1160),
.A2(n_143),
.B(n_134),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1103),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1248),
.A2(n_1093),
.B(n_1223),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1270),
.A2(n_1109),
.B1(n_1054),
.B2(n_1127),
.Y(n_1392)
);

AND2x2_ASAP7_75t_SL g1393 ( 
.A(n_1373),
.B(n_1150),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_R g1394 ( 
.A(n_1257),
.B(n_1080),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1276),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_L g1396 ( 
.A(n_1310),
.B(n_1109),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1331),
.A2(n_1176),
.B(n_1128),
.Y(n_1397)
);

AOI221xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1244),
.A2(n_1318),
.B1(n_1324),
.B2(n_1390),
.C(n_1381),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1231),
.A2(n_1128),
.B(n_1097),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1229),
.B(n_1214),
.C(n_1170),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1309),
.Y(n_1401)
);

AOI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1298),
.A2(n_1147),
.B(n_1212),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1232),
.A2(n_1147),
.B(n_1063),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1273),
.A2(n_1179),
.A3(n_1177),
.B(n_1211),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1119),
.B(n_1083),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1276),
.B(n_1139),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1267),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1358),
.B(n_1087),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1235),
.B(n_1225),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1365),
.A2(n_1131),
.B(n_1105),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1246),
.A2(n_1093),
.B(n_1223),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1363),
.B(n_1172),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1328),
.A2(n_1076),
.B(n_1060),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1233),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1297),
.A2(n_1111),
.B(n_1065),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1282),
.B(n_1142),
.C(n_1181),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1335),
.B(n_1298),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1281),
.B(n_1172),
.Y(n_1418)
);

OR2x2_ASAP7_75t_SL g1419 ( 
.A(n_1311),
.B(n_1225),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1275),
.B(n_1085),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1279),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1292),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1374),
.B(n_1192),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1365),
.A2(n_1181),
.B(n_1154),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1299),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1341),
.B(n_1042),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1296),
.A2(n_1062),
.B(n_1066),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1304),
.Y(n_1428)
);

O2A1O1Ixp5_ASAP7_75t_L g1429 ( 
.A1(n_1272),
.A2(n_1171),
.B(n_1073),
.C(n_1077),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1334),
.B(n_1044),
.Y(n_1430)
);

NAND2x1_ASAP7_75t_L g1431 ( 
.A(n_1267),
.B(n_1064),
.Y(n_1431)
);

AO31x2_ASAP7_75t_L g1432 ( 
.A1(n_1336),
.A2(n_1171),
.A3(n_1057),
.B(n_1068),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1359),
.B(n_1048),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1329),
.A2(n_1203),
.B(n_1199),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1312),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1250),
.B(n_1094),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1319),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1347),
.A2(n_1227),
.B1(n_1188),
.B2(n_1210),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1242),
.A2(n_1215),
.B(n_1187),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1234),
.A2(n_1240),
.B(n_1239),
.Y(n_1440)
);

NAND2x1_ASAP7_75t_L g1441 ( 
.A(n_1267),
.B(n_1134),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1350),
.A2(n_1159),
.B1(n_1124),
.B2(n_1142),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1255),
.B(n_1102),
.Y(n_1443)
);

AOI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1265),
.A2(n_1102),
.B(n_1110),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1269),
.B(n_1110),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1285),
.B(n_1077),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1241),
.A2(n_1222),
.B(n_1190),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1357),
.B(n_1124),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1374),
.A2(n_1210),
.B(n_1204),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1243),
.B(n_1174),
.Y(n_1450)
);

BUFx12f_ASAP7_75t_L g1451 ( 
.A(n_1386),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1353),
.A2(n_1174),
.B(n_1144),
.C(n_1184),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_SL g1453 ( 
.A(n_1361),
.B(n_1227),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1262),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1337),
.A2(n_1146),
.B(n_1195),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1358),
.B(n_1140),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1322),
.B(n_1168),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1230),
.A2(n_1227),
.B(n_1204),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1381),
.A2(n_1199),
.B(n_1194),
.Y(n_1459)
);

AO32x2_ASAP7_75t_L g1460 ( 
.A1(n_1390),
.A2(n_1145),
.A3(n_1134),
.B1(n_1194),
.B2(n_1203),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1378),
.A2(n_1144),
.B(n_1184),
.C(n_1189),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1277),
.A2(n_1227),
.B1(n_1146),
.B2(n_1189),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1336),
.A2(n_1190),
.A3(n_1180),
.B(n_1168),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1357),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1327),
.A2(n_1180),
.B(n_1166),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1244),
.A2(n_1141),
.B1(n_1140),
.B2(n_1145),
.C(n_1166),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1268),
.B(n_1133),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1388),
.Y(n_1468)
);

AO31x2_ASAP7_75t_L g1469 ( 
.A1(n_1313),
.A2(n_1133),
.A3(n_1120),
.B(n_63),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1333),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1360),
.A2(n_1254),
.B1(n_1237),
.B2(n_1245),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1314),
.A2(n_1120),
.A3(n_60),
.B(n_64),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1348),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1291),
.B(n_1141),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1338),
.A2(n_131),
.B(n_127),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1301),
.B(n_59),
.Y(n_1476)
);

AOI21xp33_ASAP7_75t_L g1477 ( 
.A1(n_1274),
.A2(n_64),
.B(n_67),
.Y(n_1477)
);

AOI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1330),
.A2(n_123),
.B(n_118),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1317),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1236),
.A2(n_110),
.B(n_104),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1349),
.A2(n_68),
.B(n_70),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1370),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1342),
.A2(n_74),
.A3(n_76),
.B(n_77),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1371),
.Y(n_1484)
);

AO31x2_ASAP7_75t_L g1485 ( 
.A1(n_1345),
.A2(n_74),
.A3(n_76),
.B(n_78),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1286),
.A2(n_1253),
.B(n_1263),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1352),
.A2(n_80),
.A3(n_82),
.B(n_84),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1316),
.A2(n_82),
.B(n_84),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1364),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1286),
.A2(n_85),
.B(n_86),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_SL g1491 ( 
.A1(n_1366),
.A2(n_85),
.B(n_86),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1377),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1247),
.A2(n_1249),
.B(n_1251),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1290),
.B(n_1368),
.C(n_1332),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1309),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1355),
.B(n_1256),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1258),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1278),
.Y(n_1499)
);

AOI21x1_ASAP7_75t_SL g1500 ( 
.A1(n_1268),
.A2(n_1300),
.B(n_1343),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1238),
.B(n_1302),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1261),
.Y(n_1503)
);

AO22x2_ASAP7_75t_L g1504 ( 
.A1(n_1325),
.A2(n_1288),
.B1(n_1303),
.B2(n_1305),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1316),
.A2(n_1306),
.B(n_1340),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1351),
.A2(n_1385),
.B(n_1379),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1376),
.A2(n_1389),
.B(n_1375),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1387),
.A2(n_1369),
.B(n_1271),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1271),
.A2(n_1308),
.B(n_1294),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1323),
.A2(n_1280),
.B(n_1283),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1383),
.A2(n_1354),
.B1(n_1372),
.B2(n_1288),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1283),
.A2(n_1340),
.B(n_1287),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1382),
.B(n_1264),
.C(n_1259),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1320),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1309),
.Y(n_1515)
);

AOI221x1_ASAP7_75t_L g1516 ( 
.A1(n_1320),
.A2(n_1307),
.B1(n_1315),
.B2(n_1289),
.C(n_1287),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1284),
.B(n_1380),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1321),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1339),
.A2(n_1356),
.B1(n_1321),
.B2(n_1354),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1260),
.B(n_1321),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1346),
.Y(n_1521)
);

OR2x6_ASAP7_75t_SL g1522 ( 
.A(n_1307),
.B(n_1315),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1267),
.A2(n_1344),
.B(n_1289),
.Y(n_1523)
);

AO31x2_ASAP7_75t_L g1524 ( 
.A1(n_1287),
.A2(n_1293),
.A3(n_1354),
.B(n_1295),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1293),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1357),
.B(n_1252),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1252),
.B(n_480),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1335),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1331),
.A2(n_1040),
.B(n_1043),
.Y(n_1529)
);

INVx6_ASAP7_75t_SL g1530 ( 
.A(n_1354),
.Y(n_1530)
);

AOI221x1_ASAP7_75t_L g1531 ( 
.A1(n_1381),
.A2(n_1101),
.B1(n_1061),
.B2(n_1390),
.C(n_1298),
.Y(n_1531)
);

AO31x2_ASAP7_75t_L g1532 ( 
.A1(n_1273),
.A2(n_1326),
.A3(n_1336),
.B(n_1313),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1309),
.Y(n_1533)
);

AOI221x1_ASAP7_75t_L g1534 ( 
.A1(n_1381),
.A2(n_1101),
.B1(n_1061),
.B2(n_1390),
.C(n_1298),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1276),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1197),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1197),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1197),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1262),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1233),
.Y(n_1540)
);

AOI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1248),
.A2(n_1086),
.B(n_1049),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1331),
.A2(n_1040),
.B(n_1043),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1335),
.B(n_1129),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1331),
.A2(n_1040),
.B(n_1043),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1335),
.B(n_1129),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1273),
.A2(n_1326),
.A3(n_1336),
.B(n_1313),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1331),
.A2(n_1061),
.B(n_892),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1335),
.B(n_1129),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1276),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1331),
.A2(n_1040),
.B(n_1043),
.Y(n_1550)
);

NAND2x1_ASAP7_75t_L g1551 ( 
.A(n_1267),
.B(n_1064),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1310),
.Y(n_1552)
);

XNOR2xp5_ASAP7_75t_L g1553 ( 
.A(n_1383),
.B(n_629),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1335),
.B(n_1129),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1324),
.A2(n_1061),
.B(n_892),
.C(n_1148),
.Y(n_1555)
);

AOI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1248),
.A2(n_1086),
.B(n_1049),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1197),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1266),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1273),
.A2(n_1326),
.A3(n_1336),
.B(n_1313),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1324),
.B(n_892),
.C(n_1061),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1331),
.A2(n_1061),
.B(n_892),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1335),
.B(n_1129),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1373),
.A2(n_911),
.B1(n_954),
.B2(n_1004),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1335),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_SL g1565 ( 
.A1(n_1453),
.A2(n_1491),
.B(n_1459),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1470),
.Y(n_1566)
);

NOR2xp67_ASAP7_75t_L g1567 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1560),
.A2(n_1555),
.B1(n_1430),
.B2(n_1400),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1394),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1414),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_SL g1571 ( 
.A1(n_1480),
.A2(n_1471),
.B(n_1496),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1545),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1398),
.A2(n_1477),
.B1(n_1494),
.B2(n_1402),
.C(n_1479),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1393),
.A2(n_1563),
.B1(n_1504),
.B2(n_1502),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1511),
.A2(n_1420),
.B1(n_1408),
.B2(n_1466),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1440),
.A2(n_1561),
.B(n_1547),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1557),
.A2(n_1411),
.B(n_1415),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1391),
.A2(n_1455),
.B(n_1500),
.Y(n_1578)
);

BUFx2_ASAP7_75t_SL g1579 ( 
.A(n_1540),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1512),
.A2(n_1505),
.B(n_1439),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1458),
.A2(n_1427),
.B(n_1541),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1473),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1504),
.A2(n_1513),
.B1(n_1412),
.B2(n_1490),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1531),
.A2(n_1534),
.B(n_1403),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1522),
.A2(n_1489),
.B1(n_1476),
.B2(n_1554),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1433),
.B(n_1437),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_L g1587 ( 
.A(n_1539),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1548),
.B(n_1562),
.Y(n_1588)
);

BUFx8_ASAP7_75t_SL g1589 ( 
.A(n_1451),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1556),
.A2(n_1397),
.B(n_1550),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1535),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1450),
.B(n_1417),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1447),
.A2(n_1544),
.B(n_1529),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1428),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1435),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1542),
.A2(n_1506),
.B(n_1507),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1395),
.B(n_1457),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1528),
.B(n_1564),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1425),
.B(n_1419),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1407),
.Y(n_1601)
);

AO22x2_ASAP7_75t_L g1602 ( 
.A1(n_1516),
.A2(n_1503),
.B1(n_1399),
.B2(n_1499),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1486),
.A2(n_1497),
.B(n_1410),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1408),
.B(n_1423),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1488),
.A2(n_1475),
.B(n_1508),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1423),
.B(n_1467),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1510),
.A2(n_1509),
.B(n_1462),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1449),
.A2(n_1493),
.B(n_1405),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1469),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1461),
.A2(n_1452),
.B(n_1523),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1406),
.B(n_1426),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1444),
.A2(n_1438),
.B(n_1514),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1429),
.A2(n_1465),
.B(n_1424),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1478),
.A2(n_1413),
.B(n_1434),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1407),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1484),
.B(n_1492),
.Y(n_1616)
);

CKINVDCx11_ASAP7_75t_R g1617 ( 
.A(n_1448),
.Y(n_1617)
);

BUFx12f_ASAP7_75t_L g1618 ( 
.A(n_1454),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1481),
.A2(n_1498),
.B(n_1418),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1528),
.B(n_1564),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1423),
.B(n_1467),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1401),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1413),
.A2(n_1434),
.B(n_1431),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1551),
.A2(n_1441),
.B(n_1468),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1401),
.Y(n_1625)
);

OAI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1392),
.A2(n_1527),
.B1(n_1396),
.B2(n_1442),
.C(n_1409),
.Y(n_1626)
);

AO22x2_ASAP7_75t_L g1627 ( 
.A1(n_1519),
.A2(n_1460),
.B1(n_1468),
.B2(n_1525),
.Y(n_1627)
);

AO31x2_ASAP7_75t_L g1628 ( 
.A1(n_1432),
.A2(n_1463),
.A3(n_1559),
.B(n_1532),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1517),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1553),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1456),
.B(n_1474),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1464),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1436),
.A2(n_1460),
.B(n_1416),
.C(n_1558),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1401),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1530),
.A2(n_1423),
.B1(n_1421),
.B2(n_1422),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1482),
.A2(n_1446),
.B(n_1518),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1521),
.A2(n_1501),
.B1(n_1526),
.B2(n_1460),
.C(n_1483),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1464),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1463),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1530),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1518),
.A2(n_1559),
.B(n_1546),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1532),
.A2(n_1559),
.B(n_1546),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1448),
.A2(n_1404),
.B(n_1469),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1495),
.A2(n_1533),
.B1(n_1515),
.B2(n_1483),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1432),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1495),
.A2(n_1533),
.B1(n_1515),
.B2(n_1483),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1485),
.A2(n_1533),
.B1(n_1515),
.B2(n_1495),
.C(n_1487),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1485),
.A2(n_1487),
.B(n_1524),
.Y(n_1648)
);

INVx5_ASAP7_75t_L g1649 ( 
.A(n_1472),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1524),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1432),
.A2(n_1463),
.B(n_1404),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1472),
.A2(n_1485),
.B(n_1487),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1539),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1654)
);

OA21x2_ASAP7_75t_L g1655 ( 
.A1(n_1440),
.A2(n_1561),
.B(n_1547),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1470),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1394),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_SL g1658 ( 
.A1(n_1453),
.A2(n_1491),
.B(n_1459),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1407),
.B(n_1365),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1543),
.B(n_911),
.Y(n_1660)
);

CKINVDCx11_ASAP7_75t_R g1661 ( 
.A(n_1539),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1395),
.B(n_1535),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1407),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1552),
.B(n_1045),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1547),
.A2(n_1561),
.B(n_1507),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1393),
.A2(n_657),
.B1(n_1100),
.B2(n_1563),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1470),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1668)
);

AOI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1560),
.A2(n_892),
.B(n_881),
.C(n_732),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1469),
.Y(n_1670)
);

AO31x2_ASAP7_75t_L g1671 ( 
.A1(n_1531),
.A2(n_1534),
.A3(n_1512),
.B(n_1555),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1440),
.A2(n_1561),
.B(n_1547),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1560),
.B(n_1061),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1555),
.A2(n_1298),
.B(n_1089),
.C(n_1560),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1555),
.A2(n_1298),
.B(n_1089),
.C(n_1560),
.Y(n_1677)
);

AO31x2_ASAP7_75t_L g1678 ( 
.A1(n_1531),
.A2(n_1534),
.A3(n_1512),
.B(n_1555),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_SL g1680 ( 
.A1(n_1453),
.A2(n_1491),
.B(n_1459),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1560),
.A2(n_1089),
.B1(n_1061),
.B2(n_911),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1547),
.A2(n_1561),
.B(n_1507),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1683)
);

INVx6_ASAP7_75t_SL g1684 ( 
.A(n_1448),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1543),
.B(n_911),
.Y(n_1685)
);

AO31x2_ASAP7_75t_L g1686 ( 
.A1(n_1531),
.A2(n_1534),
.A3(n_1512),
.B(n_1555),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1543),
.B(n_911),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1552),
.B(n_1045),
.Y(n_1688)
);

INVx6_ASAP7_75t_L g1689 ( 
.A(n_1464),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1433),
.B(n_1016),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1560),
.A2(n_1061),
.B1(n_1494),
.B2(n_881),
.Y(n_1692)
);

INVx8_ASAP7_75t_L g1693 ( 
.A(n_1423),
.Y(n_1693)
);

CKINVDCx16_ASAP7_75t_R g1694 ( 
.A(n_1394),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1543),
.B(n_911),
.Y(n_1695)
);

AO21x1_ASAP7_75t_L g1696 ( 
.A1(n_1547),
.A2(n_1390),
.B(n_1381),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1560),
.A2(n_1061),
.B(n_1555),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1469),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_L g1699 ( 
.A(n_1552),
.B(n_1045),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1560),
.A2(n_1061),
.B(n_1555),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1555),
.A2(n_1298),
.B(n_1089),
.C(n_1560),
.Y(n_1701)
);

AOI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1412),
.A2(n_1512),
.B(n_1458),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1414),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1543),
.B(n_911),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1560),
.A2(n_1061),
.B1(n_1494),
.B2(n_881),
.Y(n_1705)
);

INVx6_ASAP7_75t_L g1706 ( 
.A(n_1464),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1535),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1543),
.B(n_911),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1407),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1449),
.B(n_1448),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1470),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1560),
.A2(n_1061),
.B1(n_1494),
.B2(n_881),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1560),
.A2(n_1061),
.B(n_1555),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_SL g1716 ( 
.A(n_1414),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1560),
.A2(n_1061),
.B1(n_1494),
.B2(n_881),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1535),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1464),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1560),
.B(n_1061),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1470),
.Y(n_1722)
);

CKINVDCx8_ASAP7_75t_R g1723 ( 
.A(n_1454),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1560),
.A2(n_1061),
.B(n_1555),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1464),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1407),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1408),
.B(n_1423),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1393),
.A2(n_657),
.B1(n_1100),
.B2(n_1563),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1547),
.A2(n_1561),
.B(n_1507),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1470),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_SL g1732 ( 
.A(n_1560),
.B(n_657),
.C(n_892),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_L g1733 ( 
.A1(n_1560),
.A2(n_892),
.B(n_911),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1408),
.B(n_1423),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1537),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1681),
.A2(n_1685),
.B(n_1660),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1574),
.A2(n_1729),
.B1(n_1666),
.B2(n_1611),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1616),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1570),
.Y(n_1740)
);

INVx4_ASAP7_75t_SL g1741 ( 
.A(n_1712),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1595),
.Y(n_1742)
);

OA21x2_ASAP7_75t_L g1743 ( 
.A1(n_1614),
.A2(n_1603),
.B(n_1652),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1611),
.A2(n_1692),
.B1(n_1714),
.B2(n_1705),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1687),
.B(n_1695),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1712),
.B(n_1604),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1598),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1596),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1692),
.A2(n_1705),
.B1(n_1714),
.B2(n_1717),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1665),
.A2(n_1730),
.B(n_1682),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1608),
.A2(n_1597),
.B(n_1588),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1733),
.A2(n_1669),
.B(n_1732),
.C(n_1568),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1572),
.A2(n_1677),
.B(n_1676),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1676),
.A2(n_1701),
.B(n_1677),
.Y(n_1755)
);

OA21x2_ASAP7_75t_L g1756 ( 
.A1(n_1581),
.A2(n_1590),
.B(n_1623),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1704),
.B(n_1710),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1717),
.A2(n_1583),
.B1(n_1631),
.B2(n_1626),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1701),
.A2(n_1655),
.B(n_1576),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1609),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1576),
.A2(n_1672),
.B(n_1655),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1675),
.B(n_1721),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1675),
.B(n_1721),
.Y(n_1763)
);

BUFx2_ASAP7_75t_SL g1764 ( 
.A(n_1716),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1576),
.A2(n_1672),
.B(n_1655),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_L g1766 ( 
.A(n_1638),
.B(n_1720),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1583),
.A2(n_1631),
.B1(n_1567),
.B2(n_1635),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1585),
.B(n_1619),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1712),
.A2(n_1700),
.B(n_1697),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1592),
.B(n_1599),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1594),
.B(n_1591),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1635),
.A2(n_1657),
.B1(n_1569),
.B2(n_1694),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1715),
.A2(n_1724),
.B(n_1573),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1566),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1604),
.B(n_1728),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1709),
.B(n_1718),
.Y(n_1776)
);

NOR2xp67_ASAP7_75t_L g1777 ( 
.A(n_1638),
.B(n_1726),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1569),
.A2(n_1657),
.B1(n_1585),
.B2(n_1600),
.Y(n_1778)
);

AOI221x1_ASAP7_75t_SL g1779 ( 
.A1(n_1648),
.A2(n_1699),
.B1(n_1688),
.B2(n_1664),
.C(n_1575),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1571),
.A2(n_1584),
.B(n_1592),
.C(n_1696),
.Y(n_1780)
);

O2A1O1Ixp5_ASAP7_75t_L g1781 ( 
.A1(n_1702),
.A2(n_1643),
.B(n_1633),
.C(n_1650),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1734),
.B(n_1606),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1633),
.A2(n_1637),
.B(n_1593),
.C(n_1693),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1606),
.B(n_1621),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1630),
.A2(n_1684),
.B1(n_1620),
.B2(n_1689),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1582),
.B(n_1656),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1630),
.A2(n_1684),
.B1(n_1689),
.B2(n_1706),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1684),
.A2(n_1689),
.B1(n_1706),
.B2(n_1640),
.Y(n_1788)
);

AOI21x1_ASAP7_75t_SL g1789 ( 
.A1(n_1670),
.A2(n_1698),
.B(n_1645),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_L g1790 ( 
.A(n_1587),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1670),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1645),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1590),
.A2(n_1623),
.B(n_1642),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_SL g1794 ( 
.A1(n_1621),
.A2(n_1602),
.B(n_1671),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1731),
.B(n_1667),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1607),
.A2(n_1605),
.B(n_1610),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1713),
.B(n_1722),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_SL g1798 ( 
.A1(n_1602),
.A2(n_1678),
.B(n_1671),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1625),
.B(n_1634),
.Y(n_1799)
);

O2A1O1Ixp5_ASAP7_75t_L g1800 ( 
.A1(n_1650),
.A2(n_1639),
.B(n_1727),
.C(n_1615),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1659),
.A2(n_1601),
.B(n_1727),
.Y(n_1801)
);

AOI21x1_ASAP7_75t_SL g1802 ( 
.A1(n_1671),
.A2(n_1678),
.B(n_1686),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1706),
.A2(n_1632),
.B1(n_1703),
.B2(n_1579),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1671),
.B(n_1678),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1632),
.B(n_1663),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1629),
.B(n_1627),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1641),
.Y(n_1807)
);

OA21x2_ASAP7_75t_L g1808 ( 
.A1(n_1578),
.A2(n_1613),
.B(n_1673),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1629),
.B(n_1627),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1580),
.A2(n_1693),
.B(n_1578),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1627),
.B(n_1686),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1622),
.B(n_1617),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1647),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1723),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1617),
.Y(n_1815)
);

O2A1O1Ixp5_ASAP7_75t_L g1816 ( 
.A1(n_1639),
.A2(n_1615),
.B(n_1711),
.C(n_1601),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1693),
.A2(n_1716),
.B1(n_1644),
.B2(n_1646),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1678),
.B(n_1686),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1636),
.B(n_1622),
.Y(n_1819)
);

NOR2xp67_ASAP7_75t_L g1820 ( 
.A(n_1618),
.B(n_1711),
.Y(n_1820)
);

OA22x2_ASAP7_75t_L g1821 ( 
.A1(n_1565),
.A2(n_1658),
.B1(n_1680),
.B2(n_1624),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1622),
.B(n_1624),
.Y(n_1822)
);

AOI21x1_ASAP7_75t_SL g1823 ( 
.A1(n_1686),
.A2(n_1649),
.B(n_1644),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1622),
.B(n_1646),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1612),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1612),
.A2(n_1659),
.B(n_1651),
.C(n_1580),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1628),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1628),
.B(n_1651),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1661),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1649),
.B(n_1577),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1653),
.A2(n_1587),
.B1(n_1589),
.B2(n_1654),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1653),
.A2(n_1668),
.B(n_1735),
.Y(n_1833)
);

OA22x2_ASAP7_75t_L g1834 ( 
.A1(n_1673),
.A2(n_1674),
.B1(n_1679),
.B2(n_1683),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1691),
.B(n_1708),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1683),
.A2(n_1707),
.B1(n_1719),
.B2(n_1725),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1707),
.B(n_1719),
.Y(n_1837)
);

NOR2xp67_ASAP7_75t_L g1838 ( 
.A(n_1725),
.B(n_1736),
.Y(n_1838)
);

A2O1A1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1733),
.A2(n_1560),
.B(n_1669),
.C(n_1061),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1660),
.B(n_1685),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1841)
);

AOI21x1_ASAP7_75t_SL g1842 ( 
.A1(n_1660),
.A2(n_1687),
.B(n_1685),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1843)
);

AOI21x1_ASAP7_75t_SL g1844 ( 
.A1(n_1660),
.A2(n_1687),
.B(n_1685),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1574),
.A2(n_1729),
.B1(n_1666),
.B2(n_1611),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1847)
);

AND2x2_ASAP7_75t_SL g1848 ( 
.A(n_1576),
.B(n_1655),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1849)
);

O2A1O1Ixp5_ASAP7_75t_L g1850 ( 
.A1(n_1584),
.A2(n_1696),
.B(n_1555),
.C(n_1561),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1614),
.A2(n_1440),
.B(n_1603),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1661),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1598),
.B(n_1662),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1595),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1586),
.B(n_1690),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1660),
.B(n_1685),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1614),
.A2(n_1440),
.B(n_1603),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1609),
.Y(n_1858)
);

O2A1O1Ixp5_ASAP7_75t_L g1859 ( 
.A1(n_1584),
.A2(n_1696),
.B(n_1555),
.C(n_1561),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1609),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1616),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1570),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1591),
.Y(n_1863)
);

AOI21x1_ASAP7_75t_SL g1864 ( 
.A1(n_1660),
.A2(n_1687),
.B(n_1685),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1574),
.A2(n_1729),
.B1(n_1666),
.B2(n_1611),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1660),
.B(n_1685),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1712),
.B(n_1604),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1574),
.A2(n_1729),
.B1(n_1666),
.B2(n_1611),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1660),
.B(n_1685),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1748),
.Y(n_1870)
);

OR2x6_ASAP7_75t_L g1871 ( 
.A(n_1833),
.B(n_1752),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1742),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1750),
.A2(n_1744),
.B1(n_1758),
.B2(n_1738),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1806),
.B(n_1809),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1822),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1749),
.Y(n_1876)
);

AOI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1768),
.A2(n_1838),
.B(n_1796),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1748),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1848),
.B(n_1828),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1739),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1752),
.B(n_1751),
.Y(n_1881)
);

CKINVDCx16_ASAP7_75t_R g1882 ( 
.A(n_1812),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1762),
.B(n_1745),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1780),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1741),
.B(n_1830),
.Y(n_1885)
);

OR2x6_ASAP7_75t_L g1886 ( 
.A(n_1751),
.B(n_1769),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1834),
.A2(n_1810),
.B(n_1836),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1763),
.B(n_1854),
.Y(n_1888)
);

AOI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1835),
.A2(n_1765),
.B(n_1761),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_L g1890 ( 
.A1(n_1834),
.A2(n_1810),
.B(n_1821),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1811),
.B(n_1774),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1804),
.B(n_1818),
.Y(n_1892)
);

AO21x2_ASAP7_75t_L g1893 ( 
.A1(n_1759),
.A2(n_1825),
.B(n_1837),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1808),
.Y(n_1894)
);

AO31x2_ASAP7_75t_L g1895 ( 
.A1(n_1759),
.A2(n_1827),
.A3(n_1783),
.B(n_1755),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1830),
.Y(n_1896)
);

BUFx12f_ASAP7_75t_L g1897 ( 
.A(n_1829),
.Y(n_1897)
);

INVxp67_ASAP7_75t_SL g1898 ( 
.A(n_1780),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1792),
.B(n_1760),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1754),
.B(n_1770),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1754),
.B(n_1755),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1793),
.Y(n_1902)
);

OA21x2_ASAP7_75t_L g1903 ( 
.A1(n_1781),
.A2(n_1859),
.B(n_1850),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1792),
.B(n_1791),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1850),
.A2(n_1859),
.B(n_1800),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1851),
.B(n_1857),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1852),
.Y(n_1907)
);

AO21x2_ASAP7_75t_L g1908 ( 
.A1(n_1826),
.A2(n_1807),
.B(n_1773),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1800),
.A2(n_1813),
.B(n_1807),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1813),
.B(n_1737),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1858),
.B(n_1860),
.Y(n_1911)
);

CKINVDCx10_ASAP7_75t_R g1912 ( 
.A(n_1790),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1853),
.B(n_1757),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1851),
.B(n_1857),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1795),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1861),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1753),
.A2(n_1845),
.B1(n_1868),
.B2(n_1865),
.C(n_1839),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1746),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1756),
.Y(n_1919)
);

AO21x2_ASAP7_75t_L g1920 ( 
.A1(n_1753),
.A2(n_1797),
.B(n_1786),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1863),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1743),
.B(n_1776),
.Y(n_1922)
);

NAND4xp25_ASAP7_75t_L g1923 ( 
.A(n_1840),
.B(n_1869),
.C(n_1856),
.D(n_1866),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1819),
.Y(n_1924)
);

OA21x2_ASAP7_75t_L g1925 ( 
.A1(n_1816),
.A2(n_1798),
.B(n_1824),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1767),
.A2(n_1778),
.B(n_1772),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1831),
.B(n_1771),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1821),
.Y(n_1928)
);

BUFx2_ASAP7_75t_L g1929 ( 
.A(n_1824),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1741),
.Y(n_1930)
);

OA21x2_ASAP7_75t_L g1931 ( 
.A1(n_1798),
.A2(n_1802),
.B(n_1823),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1867),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1741),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1867),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1779),
.B(n_1849),
.Y(n_1935)
);

AOI21x1_ASAP7_75t_L g1936 ( 
.A1(n_1817),
.A2(n_1832),
.B(n_1785),
.Y(n_1936)
);

NOR2xp67_ASAP7_75t_L g1937 ( 
.A(n_1775),
.B(n_1803),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1747),
.B(n_1841),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1899),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1920),
.B(n_1843),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1874),
.B(n_1855),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1920),
.B(n_1846),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1874),
.B(n_1847),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1920),
.B(n_1799),
.Y(n_1944)
);

OAI222xp33_ASAP7_75t_L g1945 ( 
.A1(n_1873),
.A2(n_1815),
.B1(n_1787),
.B2(n_1788),
.C1(n_1782),
.C2(n_1784),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1875),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1920),
.B(n_1740),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1922),
.B(n_1802),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1879),
.B(n_1906),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1906),
.B(n_1914),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1894),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1922),
.B(n_1794),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1914),
.B(n_1794),
.Y(n_1953)
);

OR2x6_ASAP7_75t_L g1954 ( 
.A(n_1871),
.B(n_1801),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1899),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1900),
.B(n_1740),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1904),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1917),
.A2(n_1764),
.B1(n_1790),
.B2(n_1814),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1890),
.B(n_1895),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1896),
.B(n_1805),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1872),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1892),
.B(n_1789),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1872),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1895),
.B(n_1893),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1876),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1911),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1884),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1929),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1891),
.B(n_1862),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1921),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1915),
.B(n_1820),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1915),
.B(n_1842),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1893),
.B(n_1766),
.Y(n_1973)
);

OAI31xp33_ASAP7_75t_L g1974 ( 
.A1(n_1910),
.A2(n_1842),
.A3(n_1844),
.B(n_1864),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1893),
.B(n_1777),
.Y(n_1975)
);

OAI221xp5_ASAP7_75t_L g1976 ( 
.A1(n_1958),
.A2(n_1910),
.B1(n_1926),
.B2(n_1901),
.C(n_1898),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1951),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1967),
.A2(n_1926),
.B1(n_1901),
.B2(n_1882),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1949),
.B(n_1929),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1967),
.A2(n_1886),
.B1(n_1923),
.B2(n_1937),
.Y(n_1980)
);

OAI222xp33_ASAP7_75t_L g1981 ( 
.A1(n_1970),
.A2(n_1936),
.B1(n_1886),
.B2(n_1935),
.C1(n_1882),
.C2(n_1871),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1954),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1941),
.A2(n_1935),
.B1(n_1937),
.B2(n_1886),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1961),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1949),
.B(n_1924),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1939),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1961),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1963),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_R g1989 ( 
.A(n_1973),
.B(n_1903),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1963),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_SL g1991 ( 
.A1(n_1972),
.A2(n_1936),
.B(n_1934),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_L g1992 ( 
.A(n_1974),
.B(n_1947),
.C(n_1942),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1945),
.A2(n_1923),
.B(n_1886),
.Y(n_1993)
);

OAI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1974),
.A2(n_1886),
.B1(n_1871),
.B2(n_1883),
.C(n_1913),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1956),
.B(n_1870),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1940),
.B(n_1892),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1954),
.A2(n_1871),
.B1(n_1928),
.B2(n_1932),
.Y(n_1997)
);

OR2x6_ASAP7_75t_L g1998 ( 
.A(n_1954),
.B(n_1885),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_L g1999 ( 
.A(n_1947),
.B(n_1903),
.C(n_1881),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1940),
.B(n_1909),
.Y(n_2000)
);

OAI21xp33_ASAP7_75t_L g2001 ( 
.A1(n_1959),
.A2(n_1881),
.B(n_1888),
.Y(n_2001)
);

OR2x6_ASAP7_75t_L g2002 ( 
.A(n_1954),
.B(n_1885),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1965),
.Y(n_2003)
);

AND2x6_ASAP7_75t_SL g2004 ( 
.A(n_1969),
.B(n_1912),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1942),
.A2(n_1928),
.B1(n_1932),
.B2(n_1903),
.Y(n_2005)
);

OA21x2_ASAP7_75t_L g2006 ( 
.A1(n_1959),
.A2(n_1887),
.B(n_1902),
.Y(n_2006)
);

AOI222xp33_ASAP7_75t_L g2007 ( 
.A1(n_1945),
.A2(n_1878),
.B1(n_1938),
.B2(n_1888),
.C1(n_1916),
.C2(n_1880),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1968),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1950),
.B(n_1925),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1960),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1941),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1972),
.A2(n_1933),
.B1(n_1930),
.B2(n_1918),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1950),
.B(n_1925),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1941),
.B(n_1943),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1939),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1971),
.B(n_1927),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_L g2017 ( 
.A(n_1971),
.B(n_1877),
.C(n_1930),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1943),
.B(n_1907),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1973),
.B(n_1975),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1946),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_1943),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_SL g2022 ( 
.A1(n_1959),
.A2(n_1905),
.B1(n_1908),
.B2(n_1931),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1977),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_SL g2024 ( 
.A(n_1993),
.B(n_1952),
.C(n_1944),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1984),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2019),
.B(n_1950),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2000),
.Y(n_2027)
);

INVx4_ASAP7_75t_SL g2028 ( 
.A(n_1998),
.Y(n_2028)
);

BUFx8_ASAP7_75t_L g2029 ( 
.A(n_2008),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1998),
.Y(n_2030)
);

INVx4_ASAP7_75t_SL g2031 ( 
.A(n_1998),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1987),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_2002),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1996),
.B(n_1955),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2009),
.B(n_1953),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1988),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1996),
.B(n_1952),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_2018),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1990),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_SL g2040 ( 
.A1(n_1994),
.A2(n_1905),
.B(n_1973),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1992),
.B(n_1952),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2013),
.B(n_1953),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2003),
.Y(n_2043)
);

INVx5_ASAP7_75t_L g2044 ( 
.A(n_2002),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1986),
.Y(n_2045)
);

INVx4_ASAP7_75t_L g2046 ( 
.A(n_2004),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2015),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2014),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2011),
.Y(n_2049)
);

OAI21x1_ASAP7_75t_L g2050 ( 
.A1(n_2006),
.A2(n_1889),
.B(n_1919),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2021),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2000),
.B(n_1948),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1979),
.B(n_2010),
.Y(n_2053)
);

INVxp67_ASAP7_75t_SL g2054 ( 
.A(n_1989),
.Y(n_2054)
);

NAND4xp25_ASAP7_75t_L g2055 ( 
.A(n_1976),
.B(n_1964),
.C(n_1944),
.D(n_1962),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2041),
.B(n_2037),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_2044),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_2041),
.B(n_1955),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2049),
.B(n_2016),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2050),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2054),
.B(n_2020),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2054),
.B(n_2022),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2025),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2025),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2049),
.B(n_2016),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_2038),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2026),
.B(n_1979),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2026),
.B(n_1953),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2055),
.A2(n_1978),
.B1(n_2018),
.B2(n_2007),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2051),
.B(n_2017),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2034),
.B(n_1957),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_2044),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2032),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2028),
.B(n_2002),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2034),
.B(n_1966),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2036),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2036),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2035),
.B(n_2006),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2051),
.B(n_1995),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2050),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2028),
.B(n_1982),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2052),
.B(n_1966),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_2039),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2028),
.B(n_1982),
.Y(n_2084)
);

NAND2x1_ASAP7_75t_L g2085 ( 
.A(n_2040),
.B(n_1991),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2052),
.B(n_1948),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2035),
.B(n_1985),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2042),
.B(n_1985),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_2055),
.A2(n_2001),
.B1(n_1983),
.B2(n_1982),
.Y(n_2089)
);

NAND2x1p5_ASAP7_75t_L g2090 ( 
.A(n_2044),
.B(n_1905),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2050),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2024),
.A2(n_1980),
.B1(n_1881),
.B2(n_1997),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2030),
.B(n_2033),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2023),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2043),
.Y(n_2095)
);

INVx3_ASAP7_75t_SL g2096 ( 
.A(n_2046),
.Y(n_2096)
);

INVx1_ASAP7_75t_SL g2097 ( 
.A(n_2096),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2074),
.B(n_2030),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2056),
.B(n_2052),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2066),
.B(n_2038),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2074),
.B(n_2028),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2077),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2061),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2093),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2066),
.B(n_2046),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2093),
.B(n_2046),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2077),
.Y(n_2107)
);

CKINVDCx16_ASAP7_75t_R g2108 ( 
.A(n_2081),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2083),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2093),
.B(n_2046),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2056),
.B(n_2045),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_SL g2112 ( 
.A(n_2096),
.B(n_1981),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2083),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2081),
.B(n_2084),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2058),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2084),
.B(n_2033),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_2072),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2096),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2061),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2058),
.B(n_2045),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2067),
.B(n_2028),
.Y(n_2121)
);

NOR3xp33_ASAP7_75t_L g2122 ( 
.A(n_2085),
.B(n_2024),
.C(n_1999),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2070),
.B(n_2047),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2067),
.B(n_2028),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2071),
.B(n_2047),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2063),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2067),
.B(n_2031),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2063),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2070),
.B(n_2059),
.Y(n_2129)
);

A2O1A1Ixp33_ASAP7_75t_L g2130 ( 
.A1(n_2085),
.A2(n_2027),
.B(n_2044),
.C(n_2005),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2061),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2059),
.B(n_2065),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2065),
.B(n_2048),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2078),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2069),
.B(n_2048),
.Y(n_2135)
);

O2A1O1Ixp33_ASAP7_75t_SL g2136 ( 
.A1(n_2057),
.A2(n_2012),
.B(n_2027),
.C(n_2029),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2079),
.B(n_2053),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2079),
.B(n_2053),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2078),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2064),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2113),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2114),
.B(n_2087),
.Y(n_2142)
);

INVx4_ASAP7_75t_L g2143 ( 
.A(n_2108),
.Y(n_2143)
);

NAND3xp33_ASAP7_75t_L g2144 ( 
.A(n_2122),
.B(n_2062),
.C(n_2089),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2103),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_2121),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2114),
.B(n_2087),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2103),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2108),
.B(n_2087),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2103),
.B(n_2071),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_L g2151 ( 
.A(n_2106),
.B(n_1897),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2112),
.B(n_2044),
.Y(n_2152)
);

NOR2x1_ASAP7_75t_L g2153 ( 
.A(n_2097),
.B(n_2072),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2119),
.B(n_2075),
.Y(n_2154)
);

INVx1_ASAP7_75t_SL g2155 ( 
.A(n_2105),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2097),
.B(n_2062),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2121),
.B(n_2088),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2115),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_2118),
.Y(n_2159)
);

INVx1_ASAP7_75t_SL g2160 ( 
.A(n_2118),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2104),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2124),
.B(n_2088),
.Y(n_2162)
);

AO21x1_ASAP7_75t_L g2163 ( 
.A1(n_2112),
.A2(n_2062),
.B(n_2090),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2116),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_2116),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2110),
.B(n_1897),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2119),
.B(n_2075),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2098),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2119),
.B(n_2082),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2131),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2143),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2168),
.B(n_2129),
.Y(n_2172)
);

OA22x2_ASAP7_75t_L g2173 ( 
.A1(n_2143),
.A2(n_2135),
.B1(n_2100),
.B2(n_2123),
.Y(n_2173)
);

NAND3xp33_ASAP7_75t_SL g2174 ( 
.A(n_2163),
.B(n_2144),
.C(n_2152),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2161),
.Y(n_2175)
);

AOI32xp33_ASAP7_75t_L g2176 ( 
.A1(n_2143),
.A2(n_2098),
.A3(n_2127),
.B1(n_2124),
.B2(n_2132),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2164),
.B(n_2131),
.Y(n_2177)
);

AOI322xp5_ASAP7_75t_L g2178 ( 
.A1(n_2159),
.A2(n_2130),
.A3(n_2138),
.B1(n_2137),
.B2(n_2068),
.C1(n_2092),
.C2(n_2102),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2161),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2165),
.B(n_2131),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2160),
.B(n_2133),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2158),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_2151),
.B(n_2101),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2158),
.Y(n_2184)
);

AOI211xp5_ASAP7_75t_SL g2185 ( 
.A1(n_2156),
.A2(n_2136),
.B(n_2072),
.C(n_2101),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_L g2186 ( 
.A(n_2153),
.B(n_2102),
.Y(n_2186)
);

O2A1O1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_2163),
.A2(n_2109),
.B(n_2107),
.C(n_2057),
.Y(n_2187)
);

OAI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2144),
.A2(n_2101),
.B(n_2057),
.Y(n_2188)
);

XNOR2x1_ASAP7_75t_L g2189 ( 
.A(n_2155),
.B(n_2101),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2145),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2146),
.B(n_2111),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_2153),
.Y(n_2192)
);

NAND3xp33_ASAP7_75t_L g2193 ( 
.A(n_2141),
.B(n_2109),
.C(n_2107),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2145),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2186),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2194),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2192),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_2187),
.B(n_2146),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2174),
.A2(n_2149),
.B1(n_2166),
.B2(n_2162),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2192),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2171),
.B(n_1897),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2190),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2191),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2176),
.B(n_2149),
.Y(n_2204)
);

NOR2x1_ASAP7_75t_L g2205 ( 
.A(n_2193),
.B(n_2141),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2189),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2185),
.B(n_2157),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2185),
.B(n_2157),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2175),
.Y(n_2209)
);

AOI21xp33_ASAP7_75t_L g2210 ( 
.A1(n_2205),
.A2(n_2173),
.B(n_2183),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2199),
.A2(n_2206),
.B1(n_2195),
.B2(n_2198),
.Y(n_2211)
);

O2A1O1Ixp33_ASAP7_75t_L g2212 ( 
.A1(n_2198),
.A2(n_2188),
.B(n_2184),
.C(n_2182),
.Y(n_2212)
);

NAND4xp25_ASAP7_75t_L g2213 ( 
.A(n_2204),
.B(n_2178),
.C(n_2181),
.D(n_2172),
.Y(n_2213)
);

AOI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2195),
.A2(n_2173),
.B(n_2177),
.Y(n_2214)
);

AOI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2207),
.A2(n_2179),
.B1(n_2180),
.B2(n_2162),
.C(n_2142),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2207),
.B(n_2142),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2208),
.A2(n_2117),
.B(n_2148),
.Y(n_2217)
);

AOI322xp5_ASAP7_75t_L g2218 ( 
.A1(n_2206),
.A2(n_2147),
.A3(n_2127),
.B1(n_2068),
.B2(n_2078),
.C1(n_2134),
.C2(n_2139),
.Y(n_2218)
);

OAI211xp5_ASAP7_75t_L g2219 ( 
.A1(n_2208),
.A2(n_2072),
.B(n_2170),
.C(n_2148),
.Y(n_2219)
);

NAND3xp33_ASAP7_75t_L g2220 ( 
.A(n_2200),
.B(n_2170),
.C(n_2154),
.Y(n_2220)
);

AOI21xp33_ASAP7_75t_SL g2221 ( 
.A1(n_2201),
.A2(n_2154),
.B(n_2150),
.Y(n_2221)
);

AOI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2197),
.A2(n_2117),
.B(n_2150),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2216),
.Y(n_2223)
);

AOI222xp33_ASAP7_75t_L g2224 ( 
.A1(n_2211),
.A2(n_2197),
.B1(n_2203),
.B2(n_2209),
.C1(n_2202),
.C2(n_2196),
.Y(n_2224)
);

AOI221xp5_ASAP7_75t_L g2225 ( 
.A1(n_2210),
.A2(n_2147),
.B1(n_2167),
.B2(n_2140),
.C(n_2126),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2220),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2214),
.B(n_2167),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2213),
.A2(n_2126),
.B1(n_2140),
.B2(n_2128),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2219),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2223),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_2229),
.B(n_2217),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2227),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2226),
.B(n_2222),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2225),
.A2(n_2212),
.B(n_2215),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2224),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2228),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2223),
.B(n_2221),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2234),
.A2(n_2218),
.B(n_2128),
.C(n_2169),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2237),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2232),
.A2(n_2235),
.B(n_2233),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_L g2241 ( 
.A(n_2236),
.B(n_2169),
.C(n_2099),
.Y(n_2241)
);

NOR2x1_ASAP7_75t_SL g2242 ( 
.A(n_2230),
.B(n_2111),
.Y(n_2242)
);

XNOR2xp5_ASAP7_75t_L g2243 ( 
.A(n_2231),
.B(n_1912),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2231),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_2239),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2242),
.B(n_2120),
.Y(n_2246)
);

NOR3x1_ASAP7_75t_L g2247 ( 
.A(n_2241),
.B(n_2099),
.C(n_2120),
.Y(n_2247)
);

INVxp67_ASAP7_75t_SL g2248 ( 
.A(n_2243),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2244),
.B(n_2125),
.Y(n_2249)
);

INVxp67_ASAP7_75t_L g2250 ( 
.A(n_2249),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2248),
.B(n_2240),
.Y(n_2251)
);

NOR4xp25_ASAP7_75t_L g2252 ( 
.A(n_2246),
.B(n_2238),
.C(n_2139),
.D(n_2134),
.Y(n_2252)
);

OAI221xp5_ASAP7_75t_L g2253 ( 
.A1(n_2252),
.A2(n_2245),
.B1(n_2247),
.B2(n_2125),
.C(n_2134),
.Y(n_2253)
);

AOI322xp5_ASAP7_75t_L g2254 ( 
.A1(n_2251),
.A2(n_2250),
.A3(n_2139),
.B1(n_2060),
.B2(n_2080),
.C1(n_2091),
.C2(n_2068),
.Y(n_2254)
);

OAI22x1_ASAP7_75t_L g2255 ( 
.A1(n_2253),
.A2(n_2090),
.B1(n_2044),
.B2(n_2094),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_2254),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_L g2257 ( 
.A(n_2253),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2257),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2256),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_L g2260 ( 
.A(n_2255),
.B(n_2086),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2259),
.B(n_2086),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_SL g2262 ( 
.A1(n_2261),
.A2(n_2258),
.B1(n_2260),
.B2(n_2090),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2262),
.A2(n_2080),
.B1(n_2060),
.B2(n_2091),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_2263),
.B(n_2060),
.Y(n_2264)
);

AOI221x1_ASAP7_75t_L g2265 ( 
.A1(n_2264),
.A2(n_2080),
.B1(n_2091),
.B2(n_2094),
.C(n_2064),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2265),
.A2(n_2094),
.B1(n_2095),
.B2(n_2076),
.Y(n_2266)
);

AOI211xp5_ASAP7_75t_L g2267 ( 
.A1(n_2266),
.A2(n_2095),
.B(n_2073),
.C(n_2076),
.Y(n_2267)
);


endmodule