module real_jpeg_5959_n_31 (n_17, n_8, n_0, n_21, n_2, n_185, n_29, n_180, n_10, n_178, n_9, n_12, n_24, n_176, n_6, n_28, n_183, n_177, n_179, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_30, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_185;
input n_29;
input n_180;
input n_10;
input n_178;
input n_9;
input n_12;
input n_24;
input n_176;
input n_6;
input n_28;
input n_183;
input n_177;
input n_179;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_1),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_51),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_48),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_5),
.B(n_143),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_104),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_74),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_13),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_15),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_18),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_18),
.B(n_160),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_19),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_19),
.B(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_21),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_22),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_23),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_120),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_25),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_28),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_29),
.B(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_30),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_62),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_169),
.Y(n_31)
);

AO21x1_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_41),
.B(n_167),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_35),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_72),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_37),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_37),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_40),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_166),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_43),
.B(n_48),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_45),
.B(n_144),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_48),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_165),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_53),
.B(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_155),
.B(n_162),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_136),
.B(n_149),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_76),
.B(n_124),
.C(n_133),
.Y(n_59)
);

NOR4xp25_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.C(n_70),
.D(n_73),
.Y(n_60)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_90),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_119),
.B(n_123),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_112),
.B(n_118),
.Y(n_77)
);

AO221x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_86),
.B1(n_109),
.B2(n_110),
.C(n_111),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B(n_108),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_103),
.B(n_107),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_102),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_101),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_117),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_130),
.C(n_131),
.D(n_132),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_145),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_145),
.B(n_150),
.C(n_153),
.D(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_176),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_177),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_178),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_179),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_180),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_181),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_182),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_183),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_184),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_185),
.Y(n_121)
);


endmodule