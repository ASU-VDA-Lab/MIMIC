module real_jpeg_7450_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_1),
.A2(n_35),
.B1(n_48),
.B2(n_57),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_2),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_2),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_2),
.A2(n_41),
.B1(n_255),
.B2(n_274),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_2),
.A2(n_255),
.B1(n_308),
.B2(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_2),
.A2(n_109),
.B1(n_194),
.B2(n_255),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_47),
.B1(n_149),
.B2(n_153),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_4),
.A2(n_47),
.B1(n_234),
.B2(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_5),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_57),
.B1(n_108),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_5),
.A2(n_108),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_5),
.A2(n_108),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_7),
.Y(n_322)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_7),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_8),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_8),
.A2(n_164),
.B1(n_182),
.B2(n_241),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_8),
.A2(n_182),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_8),
.A2(n_182),
.B1(n_342),
.B2(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_9),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_10),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_89),
.B1(n_131),
.B2(n_176),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_10),
.A2(n_89),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_10),
.A2(n_89),
.B1(n_223),
.B2(n_254),
.Y(n_402)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_12),
.Y(n_181)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_12),
.Y(n_378)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_12),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_144),
.B1(n_148),
.B2(n_151),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_13),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_151),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_151),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_13),
.A2(n_151),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_14),
.A2(n_82),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_14),
.B(n_67),
.C(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_14),
.B(n_136),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_14),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_14),
.B(n_83),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_14),
.B(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_16),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_16),
.A2(n_70),
.B1(n_78),
.B2(n_164),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_16),
.A2(n_78),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_213),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_211),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_186),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_20),
.B(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_121),
.C(n_160),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_21),
.A2(n_22),
.B1(n_121),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_84),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_23),
.A2(n_24),
.B(n_86),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B1(n_86),
.B2(n_120),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_24),
.A2(n_45),
.B1(n_120),
.B2(n_411),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_25),
.A2(n_34),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_25),
.A2(n_240),
.B(n_244),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_25),
.A2(n_225),
.B(n_244),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_25),
.A2(n_267),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_26),
.B(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_26),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_26),
.A2(n_32),
.B1(n_319),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_26),
.A2(n_383),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_27),
.Y(n_166)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_28),
.Y(n_321)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_30),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_37),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_38),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_44),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_45),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_55),
.B1(n_77),
.B2(n_83),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_46),
.A2(n_55),
.B1(n_83),
.B2(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_51),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_51),
.Y(n_257)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_55),
.A2(n_77),
.B1(n_83),
.B2(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_55),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_55),
.B(n_227),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_56)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

INVx5_ASAP7_75t_SL g301 ( 
.A(n_63),
.Y(n_301)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_64),
.Y(n_224)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_66),
.A2(n_158),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_66),
.A2(n_252),
.B(n_258),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_66),
.A2(n_258),
.B(n_402),
.Y(n_401)
);

AOI22x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_71),
.Y(n_248)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g329 ( 
.A(n_82),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_83),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_83),
.Y(n_297)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_106),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_88),
.Y(n_191)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_94),
.B(n_225),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_94),
.A2(n_179),
.B1(n_180),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_101),
.B2(n_104),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_95),
.A2(n_365),
.A3(n_368),
.B1(n_370),
.B2(n_375),
.Y(n_364)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_99),
.Y(n_205)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_100),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_100),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_100),
.Y(n_315)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_106),
.A2(n_192),
.B(n_424),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_110),
.Y(n_369)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_114),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_114),
.A2(n_391),
.B(n_394),
.Y(n_390)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_121),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_155),
.B(n_159),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_156),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_136),
.B1(n_142),
.B2(n_152),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_124),
.A2(n_304),
.B(n_310),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_124),
.B(n_346),
.Y(n_345)
);

AOI22x1_ASAP7_75t_L g425 ( 
.A1(n_124),
.A2(n_136),
.B1(n_346),
.B2(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_124),
.A2(n_310),
.B(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_143),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_125),
.A2(n_177),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_125),
.A2(n_177),
.B1(n_341),
.B2(n_397),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_126)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_127),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_130),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_135),
.Y(n_305)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_135),
.Y(n_367)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_135),
.Y(n_374)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_136)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g323 ( 
.A1(n_148),
.A2(n_307),
.A3(n_324),
.B1(n_325),
.B2(n_329),
.Y(n_323)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_150),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_187),
.CI(n_188),
.CON(n_186),
.SN(n_186)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_160),
.B(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_174),
.C(n_178),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_161),
.B(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_162),
.B(n_167),
.Y(n_436)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_163),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_165),
.Y(n_286)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_168),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g324 ( 
.A(n_170),
.Y(n_324)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_174),
.B(n_178),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_175),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_177),
.B(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_177),
.A2(n_341),
.B(n_345),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B(n_185),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_185),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_186),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_210),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_209),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_222),
.B(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_199),
.A2(n_252),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_199),
.A2(n_226),
.B(n_298),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_199),
.A2(n_297),
.B1(n_402),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI311xp33_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_405),
.A3(n_444),
.B1(n_462),
.C1(n_467),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_358),
.B(n_404),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_332),
.B(n_357),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_291),
.B(n_331),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_261),
.B(n_290),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_238),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_220),
.B(n_238),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_221),
.A2(n_229),
.B1(n_230),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_225),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_225),
.B(n_376),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_SL g391 ( 
.A1(n_225),
.A2(n_375),
.B(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_249),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_250),
.C(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_259),
.B2(n_260),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_282),
.B(n_289),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_271),
.B(n_281),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_280),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_280),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_277),
.B(n_279),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_318),
.B(n_322),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_287),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_293),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_316),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_302),
.B2(n_303),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_302),
.C(n_316),
.Y(n_333)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_323),
.Y(n_338)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_333),
.B(n_334),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_339),
.B2(n_356),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_338),
.C(n_356),
.Y(n_359)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_347),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_348),
.C(n_349),
.Y(n_385)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_359),
.B(n_360),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_388),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_361)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_379),
.B2(n_380),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_364),
.B(n_379),
.Y(n_440)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_385),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_385),
.B(n_386),
.C(n_388),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_395),
.B2(n_403),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_396),
.C(n_401),
.Y(n_453)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_430),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g462 ( 
.A1(n_406),
.A2(n_430),
.B(n_463),
.C(n_466),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_427),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_407),
.B(n_427),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.C(n_412),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g443 ( 
.A(n_408),
.B(n_410),
.CI(n_412),
.CON(n_443),
.SN(n_443)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_422),
.C(n_425),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_416),
.Y(n_452)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_422),
.A2(n_423),
.B1(n_425),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_425),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_443),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_436),
.C(n_437),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_432),
.A2(n_433),
.B1(n_436),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.C(n_441),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_438),
.A2(n_439),
.B1(n_441),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_443),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_457),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_464),
.B(n_465),
.Y(n_463)
);

NOR2x1_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_454),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_454),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_451),
.C(n_453),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_453),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_459),
.Y(n_464)
);


endmodule