module fake_aes_2895_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVxp33_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_5), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
AOI211xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_0), .B(n_1), .C(n_2), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_12), .B(n_0), .Y(n_21) );
AND2x6_ASAP7_75t_L g22 ( .A(n_11), .B(n_7), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx3_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
INVx3_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_28), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_29), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_31), .Y(n_34) );
OAI222xp33_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_23), .B1(n_28), .B2(n_18), .C1(n_17), .C2(n_29), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
BUFx2_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
OAI221xp5_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_29), .B1(n_28), .B2(n_3), .C(n_1), .Y(n_38) );
BUFx2_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
AOI322xp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_10), .A3(n_28), .B1(n_29), .B2(n_34), .C1(n_35), .C2(n_40), .Y(n_41) );
endmodule