module fake_ariane_2159_n_1541 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1541);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1541;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_137;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_136;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_135;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_138;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_134;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_140;
wire n_725;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_139;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_2),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_33),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_79),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_71),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_63),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_60),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_38),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_37),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_78),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_56),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_107),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_22),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_45),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_14),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_55),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_35),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_64),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_57),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_87),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_38),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_88),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_68),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_9),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_35),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_43),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_10),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_82),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_46),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_12),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_118),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_100),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_20),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_52),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_20),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_33),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_22),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_12),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_67),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_34),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_39),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_25),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_90),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_51),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_31),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_36),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_61),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_17),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_99),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_23),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_24),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_9),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_121),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_115),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_84),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_70),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_123),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_52),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_105),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_120),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_24),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_177),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_142),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_152),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_185),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVxp33_ASAP7_75t_SL g285 ( 
.A(n_269),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_196),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_168),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_135),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_169),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_135),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_207),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_157),
.B(n_0),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_260),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_153),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_224),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_257),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_182),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_219),
.B(n_0),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_198),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_208),
.B(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_158),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_257),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_182),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_158),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_179),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_180),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_188),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_153),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_191),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_162),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_194),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_200),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_202),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_200),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_198),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_227),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_239),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_239),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_227),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_233),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_139),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_211),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_148),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_212),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_214),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_174),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_216),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_240),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_240),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_279),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_283),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_299),
.B(n_178),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_296),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_278),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_195),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_286),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_145),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_277),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_312),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_287),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_280),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_288),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_282),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_284),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_289),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_304),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_289),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_304),
.B(n_293),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_305),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_319),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_320),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_321),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_290),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_325),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_290),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_330),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_292),
.B(n_146),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_292),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_312),
.A2(n_155),
.B(n_147),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_295),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_298),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_337),
.B(n_134),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_340),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_313),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_315),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_342),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_315),
.B(n_156),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_328),
.B(n_159),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_347),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_316),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_350),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_R g422 ( 
.A(n_275),
.B(n_276),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_387),
.B(n_164),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_332),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_394),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_362),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

BUFx4f_ASAP7_75t_L g441 ( 
.A(n_419),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_364),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_364),
.B(n_165),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_360),
.A2(n_285),
.B1(n_310),
.B2(n_314),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_422),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_341),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_366),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_366),
.A2(n_301),
.B1(n_324),
.B2(n_178),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_366),
.A2(n_317),
.B1(n_176),
.B2(n_183),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NOR2x1p5_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_241),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_365),
.B(n_333),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_412),
.A2(n_258),
.B1(n_204),
.B2(n_217),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_369),
.B(n_166),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_421),
.A2(n_218),
.B1(n_221),
.B2(n_223),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_369),
.B(n_336),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_362),
.A2(n_199),
.B1(n_259),
.B2(n_256),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_356),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_SL g475 ( 
.A1(n_380),
.A2(n_346),
.B(n_343),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_423),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_382),
.B(n_384),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_368),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_372),
.B(n_336),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_385),
.A2(n_386),
.B1(n_390),
.B2(n_388),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_372),
.B(n_172),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_403),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_376),
.B(n_377),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_377),
.B(n_338),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_378),
.B(n_184),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVxp33_ASAP7_75t_SL g491 ( 
.A(n_406),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_379),
.B(n_201),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_379),
.B(n_338),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_361),
.B(n_339),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_393),
.B(n_149),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_353),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_391),
.B(n_205),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_363),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_339),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_353),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_408),
.B(n_343),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_353),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_409),
.A2(n_163),
.B1(n_231),
.B2(n_252),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_416),
.B(n_170),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx4_ASAP7_75t_SL g512 ( 
.A(n_353),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_351),
.A2(n_248),
.B1(n_266),
.B2(n_244),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_353),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_408),
.A2(n_245),
.B1(n_259),
.B2(n_266),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_352),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_359),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_420),
.B(n_345),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_418),
.A2(n_253),
.B1(n_242),
.B2(n_237),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_373),
.B(n_322),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_345),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_397),
.B(n_149),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_392),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_363),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_358),
.B(n_206),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_354),
.B(n_346),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_407),
.B(n_241),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_400),
.A2(n_271),
.B1(n_226),
.B2(n_267),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_400),
.B(n_149),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_367),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_367),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_374),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_383),
.B(n_149),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_417),
.B(n_273),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_355),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_419),
.B(n_149),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_355),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_419),
.B(n_270),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_355),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_355),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_371),
.B(n_134),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_362),
.A2(n_249),
.B1(n_248),
.B2(n_252),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_419),
.B(n_326),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_419),
.B(n_303),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_371),
.B(n_137),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_371),
.B(n_137),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_387),
.B(n_238),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_506),
.B(n_138),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_451),
.B(n_244),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_506),
.B(n_140),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_498),
.B1(n_445),
.B2(n_448),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_483),
.B(n_140),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_141),
.Y(n_564)
);

O2A1O1Ixp5_ASAP7_75t_L g565 ( 
.A1(n_426),
.A2(n_251),
.B(n_262),
.C(n_263),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_490),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_441),
.B(n_220),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_526),
.B(n_141),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_498),
.B(n_143),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_490),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_498),
.B(n_144),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_222),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_454),
.B(n_144),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_434),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_454),
.B(n_150),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_546),
.A2(n_445),
.B1(n_448),
.B2(n_437),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_444),
.B(n_154),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_435),
.B(n_225),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_475),
.A2(n_274),
.B(n_160),
.C(n_307),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_523),
.B(n_245),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_510),
.A2(n_439),
.B1(n_552),
.B2(n_544),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_481),
.B(n_256),
.C(n_246),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_327),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_486),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_532),
.B(n_161),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_303),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_518),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_491),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_552),
.B(n_228),
.Y(n_593)
);

BUFx8_ASAP7_75t_L g594 ( 
.A(n_520),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_495),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_432),
.B(n_232),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_431),
.B(n_209),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_528),
.B(n_246),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_451),
.B(n_209),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_551),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_432),
.B(n_436),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_478),
.B(n_243),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_542),
.B(n_249),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_525),
.B(n_306),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_533),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_511),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_453),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_549),
.A2(n_555),
.B1(n_554),
.B2(n_487),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_433),
.A2(n_268),
.B1(n_255),
.B2(n_235),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_456),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_436),
.B(n_236),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_456),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_517),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_436),
.B(n_255),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_440),
.B(n_254),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_494),
.B(n_264),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_540),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_450),
.B(n_268),
.C(n_265),
.Y(n_625)
);

NAND2x1p5_ASAP7_75t_L g626 ( 
.A(n_452),
.B(n_250),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_548),
.A2(n_470),
.B1(n_442),
.B2(n_447),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_550),
.B(n_264),
.C(n_265),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_461),
.B(n_462),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_466),
.B(n_272),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_468),
.B(n_261),
.Y(n_631)
);

AND2x4_ASAP7_75t_SL g632 ( 
.A(n_538),
.B(n_306),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_455),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_458),
.A2(n_457),
.B1(n_539),
.B2(n_473),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_460),
.B(n_307),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_464),
.B(n_308),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_541),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_424),
.B(n_3),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_167),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_502),
.B(n_173),
.Y(n_640)
);

OAI22x1_ASAP7_75t_L g641 ( 
.A1(n_479),
.A2(n_508),
.B1(n_513),
.B2(n_515),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_472),
.B(n_480),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_446),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_429),
.B(n_3),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_472),
.B(n_181),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_541),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_480),
.B(n_488),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_446),
.B(n_469),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_455),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_488),
.B(n_308),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_471),
.B(n_4),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_503),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_4),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_493),
.B(n_234),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_541),
.B(n_544),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_503),
.Y(n_660)
);

BUFx4_ASAP7_75t_L g661 ( 
.A(n_541),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_463),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_509),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_541),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_545),
.B(n_547),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_545),
.B(n_5),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_521),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_547),
.B(n_215),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_497),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_519),
.B(n_213),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_519),
.B(n_197),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_521),
.B(n_544),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_530),
.Y(n_676)
);

INVxp33_ASAP7_75t_L g677 ( 
.A(n_531),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_427),
.B(n_6),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_501),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_544),
.B(n_193),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_437),
.A2(n_190),
.B1(n_170),
.B2(n_189),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_452),
.B(n_190),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_544),
.B(n_192),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_529),
.B(n_170),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_437),
.A2(n_190),
.B1(n_170),
.B2(n_186),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_585),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_612),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_661),
.B(n_518),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_643),
.B(n_469),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_614),
.A2(n_449),
.B(n_448),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_583),
.B(n_482),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_558),
.A2(n_556),
.B(n_482),
.C(n_489),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_650),
.B(n_489),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_592),
.B(n_492),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_595),
.B(n_492),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_560),
.B(n_428),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_667),
.A2(n_484),
.B(n_465),
.Y(n_698)
);

AO22x1_ASAP7_75t_L g699 ( 
.A1(n_583),
.A2(n_499),
.B1(n_527),
.B2(n_537),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_557),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_564),
.B(n_430),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_610),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_683),
.A2(n_505),
.B(n_514),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_662),
.B(n_524),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_580),
.B(n_536),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_629),
.A2(n_459),
.B(n_485),
.C(n_467),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_669),
.A2(n_449),
.B(n_514),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_645),
.B(n_187),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_561),
.A2(n_529),
.B1(n_505),
.B2(n_514),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_679),
.A2(n_505),
.B(n_485),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_SL g711 ( 
.A1(n_638),
.A2(n_531),
.B(n_7),
.C(n_8),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_629),
.A2(n_507),
.B(n_443),
.C(n_190),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_SL g713 ( 
.A1(n_685),
.A2(n_537),
.B(n_527),
.C(n_499),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_576),
.B(n_477),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_576),
.B(n_477),
.Y(n_715)
);

AOI21x1_ASAP7_75t_L g716 ( 
.A1(n_685),
.A2(n_512),
.B(n_500),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_627),
.A2(n_443),
.B1(n_11),
.B2(n_18),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_679),
.A2(n_499),
.B(n_527),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_633),
.A2(n_512),
.B(n_499),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_588),
.B(n_499),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_633),
.A2(n_537),
.B(n_527),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_596),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_6),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_596),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_652),
.A2(n_537),
.B(n_527),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_594),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_573),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_575),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_578),
.B(n_620),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_651),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_620),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_578),
.B(n_30),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_644),
.A2(n_72),
.B(n_114),
.Y(n_733)
);

NOR2x1_ASAP7_75t_R g734 ( 
.A(n_611),
.B(n_32),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_619),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_632),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_638),
.A2(n_34),
.B(n_36),
.C(n_40),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_579),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_646),
.B(n_44),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_586),
.B(n_47),
.Y(n_740)
);

AOI21x1_ASAP7_75t_L g741 ( 
.A1(n_675),
.A2(n_83),
.B(n_93),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_648),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_658),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_581),
.B(n_74),
.Y(n_745)
);

O2A1O1Ixp5_ASAP7_75t_L g746 ( 
.A1(n_647),
.A2(n_75),
.B(n_85),
.C(n_89),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_664),
.A2(n_672),
.B(n_680),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_557),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_567),
.B(n_572),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_624),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_671),
.A2(n_673),
.B(n_674),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_598),
.A2(n_617),
.B(n_605),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_567),
.B(n_572),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_598),
.A2(n_617),
.B(n_605),
.Y(n_754)
);

OR2x4_ASAP7_75t_L g755 ( 
.A(n_593),
.B(n_603),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_677),
.B(n_566),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_682),
.A2(n_686),
.B(n_599),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_563),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_634),
.A2(n_655),
.B1(n_651),
.B2(n_642),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_589),
.B(n_632),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_563),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_623),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_574),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_654),
.B(n_569),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_624),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_635),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_570),
.B(n_625),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_571),
.B(n_600),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_651),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_647),
.A2(n_657),
.B(n_668),
.C(n_678),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_631),
.B(n_636),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_584),
.Y(n_772)
);

AOI221xp5_ASAP7_75t_SL g773 ( 
.A1(n_615),
.A2(n_622),
.B1(n_678),
.B2(n_630),
.C(n_621),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_559),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_668),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_657),
.B(n_602),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_593),
.B(n_609),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_604),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_584),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_608),
.B(n_582),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_683),
.A2(n_656),
.B(n_660),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_584),
.B(n_653),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_626),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_562),
.B(n_640),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_639),
.B(n_618),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_590),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_659),
.B(n_686),
.Y(n_788)
);

OA22x2_ASAP7_75t_L g789 ( 
.A1(n_641),
.A2(n_618),
.B1(n_587),
.B2(n_676),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_628),
.B(n_670),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_682),
.A2(n_613),
.B(n_587),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_591),
.A2(n_656),
.B(n_663),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_591),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_597),
.A2(n_660),
.B1(n_665),
.B2(n_601),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_590),
.Y(n_795)
);

AO21x1_ASAP7_75t_L g796 ( 
.A1(n_597),
.A2(n_616),
.B(n_665),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_601),
.A2(n_670),
.B1(n_663),
.B2(n_613),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_616),
.A2(n_676),
.B(n_653),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_590),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_653),
.A2(n_681),
.B(n_684),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_565),
.A2(n_637),
.B(n_649),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_666),
.Y(n_802)
);

CKINVDCx6p67_ASAP7_75t_R g803 ( 
.A(n_596),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_607),
.A2(n_667),
.B(n_650),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_577),
.B(n_441),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_643),
.B(n_650),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_643),
.B(n_650),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_584),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_577),
.B(n_441),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_595),
.Y(n_810)
);

OAI321xp33_ASAP7_75t_L g811 ( 
.A1(n_634),
.A2(n_508),
.A3(n_625),
.B1(n_655),
.B2(n_682),
.C(n_686),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_576),
.B(n_607),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_607),
.A2(n_667),
.B(n_650),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_607),
.A2(n_667),
.B(n_650),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_595),
.Y(n_815)
);

AND2x6_ASAP7_75t_L g816 ( 
.A(n_661),
.B(n_581),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_558),
.A2(n_491),
.B(n_560),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_643),
.B(n_650),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_558),
.A2(n_564),
.B(n_568),
.C(n_560),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_643),
.B(n_650),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_585),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_557),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_595),
.B(n_419),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_585),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_595),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_650),
.A2(n_643),
.B1(n_560),
.B2(n_564),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_650),
.A2(n_643),
.B1(n_560),
.B2(n_564),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_557),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_643),
.B(n_650),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_557),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_557),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_558),
.A2(n_564),
.B(n_568),
.C(n_560),
.Y(n_832)
);

OA22x2_ASAP7_75t_L g833 ( 
.A1(n_634),
.A2(n_641),
.B1(n_632),
.B2(n_552),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_557),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_643),
.A2(n_444),
.B(n_629),
.C(n_475),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_558),
.A2(n_564),
.B(n_568),
.C(n_560),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_596),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_771),
.B(n_702),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_779),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_803),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_775),
.A2(n_770),
.B1(n_729),
.B2(n_749),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_779),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_702),
.B(n_753),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_777),
.B(n_705),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_759),
.B(n_806),
.Y(n_845)
);

NOR2x1_ASAP7_75t_SL g846 ( 
.A(n_807),
.B(n_818),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_835),
.A2(n_819),
.B(n_836),
.C(n_832),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_817),
.B(n_820),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_810),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_759),
.B(n_829),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_779),
.Y(n_851)
);

AND2x2_ASAP7_75t_SL g852 ( 
.A(n_788),
.B(n_730),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_833),
.A2(n_788),
.B1(n_704),
.B2(n_757),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_795),
.B(n_772),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_689),
.Y(n_855)
);

AO31x2_ASAP7_75t_L g856 ( 
.A1(n_796),
.A2(n_706),
.A3(n_826),
.B(n_827),
.Y(n_856)
);

AOI21xp33_ASAP7_75t_L g857 ( 
.A1(n_811),
.A2(n_833),
.B(n_732),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_805),
.B(n_809),
.C(n_694),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_752),
.A2(n_791),
.B(n_798),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_823),
.B(n_810),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_748),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_812),
.A2(n_745),
.B(n_751),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_739),
.A2(n_809),
.B(n_805),
.C(n_738),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_722),
.Y(n_864)
);

AOI21xp33_ASAP7_75t_L g865 ( 
.A1(n_756),
.A2(n_767),
.B(n_766),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_812),
.A2(n_745),
.B(n_733),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_768),
.B(n_756),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_687),
.B(n_688),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_825),
.A2(n_724),
.B1(n_815),
.B2(n_760),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_735),
.B(n_762),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_821),
.B(n_824),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_692),
.B(n_825),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_769),
.B(n_736),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_792),
.A2(n_716),
.B(n_741),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_692),
.B(n_726),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_690),
.A2(n_693),
.B(n_740),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_710),
.A2(n_747),
.B(n_698),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_769),
.B(n_755),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_714),
.A2(n_715),
.B(n_783),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_692),
.B(n_837),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_837),
.B(n_723),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_723),
.B(n_781),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_781),
.B(n_784),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_695),
.B(n_696),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_785),
.A2(n_697),
.B1(n_701),
.B2(n_764),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_714),
.A2(n_715),
.B(n_783),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_L g887 ( 
.A1(n_767),
.A2(n_789),
.B(n_780),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_744),
.B(n_774),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_758),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_778),
.B(n_765),
.Y(n_890)
);

AO31x2_ASAP7_75t_L g891 ( 
.A1(n_709),
.A2(n_712),
.A3(n_786),
.B(n_717),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_772),
.B(n_808),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_761),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_784),
.B(n_778),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_737),
.B(n_731),
.C(n_743),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_816),
.B(n_755),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_790),
.B(n_787),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_816),
.B(n_689),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_746),
.A2(n_713),
.B(n_719),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_816),
.B(n_689),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_801),
.A2(n_718),
.B(n_794),
.Y(n_901)
);

AO31x2_ASAP7_75t_L g902 ( 
.A1(n_720),
.A2(n_763),
.A3(n_831),
.B(n_830),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_SL g903 ( 
.A1(n_727),
.A2(n_728),
.B1(n_742),
.B2(n_799),
.C(n_773),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_787),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_816),
.B(n_689),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_794),
.A2(n_797),
.B(n_828),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_793),
.A2(n_834),
.B(n_822),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_711),
.B(n_708),
.C(n_750),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_689),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_721),
.A2(n_725),
.B(n_711),
.C(n_802),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_816),
.B(n_789),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_SL g912 ( 
.A1(n_699),
.A2(n_770),
.B(n_775),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_734),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_771),
.B(n_702),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_771),
.B(n_702),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_782),
.A2(n_703),
.B(n_800),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_729),
.A2(n_491),
.B1(n_483),
.B2(n_481),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_779),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_823),
.B(n_439),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_825),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_804),
.A2(n_814),
.B(n_813),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_687),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_825),
.Y(n_923)
);

OAI21x1_ASAP7_75t_L g924 ( 
.A1(n_782),
.A2(n_707),
.B(n_691),
.Y(n_924)
);

AOI21xp33_ASAP7_75t_L g925 ( 
.A1(n_729),
.A2(n_775),
.B(n_283),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_803),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_702),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_782),
.A2(n_707),
.B(n_691),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_689),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_803),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_804),
.A2(n_814),
.B(n_813),
.Y(n_931)
);

AOI21x1_ASAP7_75t_L g932 ( 
.A1(n_752),
.A2(n_754),
.B(n_812),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_823),
.B(n_439),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_803),
.Y(n_934)
);

OAI22x1_ASAP7_75t_L g935 ( 
.A1(n_769),
.A2(n_583),
.B1(n_420),
.B2(n_730),
.Y(n_935)
);

AO31x2_ASAP7_75t_L g936 ( 
.A1(n_796),
.A2(n_770),
.A3(n_706),
.B(n_826),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_707),
.B(n_691),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_729),
.A2(n_491),
.B1(n_483),
.B2(n_481),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_810),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_700),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_782),
.A2(n_703),
.B(n_800),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_722),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_803),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_771),
.B(n_702),
.Y(n_944)
);

BUFx8_ASAP7_75t_L g945 ( 
.A(n_726),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_771),
.B(n_702),
.Y(n_946)
);

INVx8_ASAP7_75t_L g947 ( 
.A(n_689),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_771),
.B(n_702),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_771),
.B(n_702),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_803),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_782),
.A2(n_703),
.B(n_800),
.Y(n_951)
);

AOI21x1_ASAP7_75t_SL g952 ( 
.A1(n_729),
.A2(n_775),
.B(n_776),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_752),
.A2(n_754),
.B(n_812),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_770),
.A2(n_796),
.B(n_707),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_823),
.B(n_439),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_749),
.B(n_753),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_803),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_SL g958 ( 
.A1(n_729),
.A2(n_481),
.B(n_380),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_771),
.B(n_702),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_SL g960 ( 
.A1(n_770),
.A2(n_775),
.B(n_753),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_933),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_841),
.A2(n_925),
.B(n_958),
.C(n_956),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_860),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_921),
.A2(n_931),
.B(n_960),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_922),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_868),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_920),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_870),
.Y(n_968)
);

AND2x2_ASAP7_75t_SL g969 ( 
.A(n_900),
.B(n_852),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_844),
.B(n_843),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_956),
.A2(n_858),
.B1(n_863),
.B2(n_912),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_845),
.B(n_850),
.Y(n_972)
);

INVx3_ASAP7_75t_SL g973 ( 
.A(n_840),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_863),
.A2(n_858),
.B(n_847),
.C(n_895),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_900),
.B(n_929),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_943),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_929),
.B(n_855),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_871),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_855),
.Y(n_979)
);

INVxp33_ASAP7_75t_L g980 ( 
.A(n_923),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_867),
.B(n_838),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_890),
.Y(n_982)
);

AO32x2_ASAP7_75t_L g983 ( 
.A1(n_885),
.A2(n_952),
.A3(n_857),
.B1(n_936),
.B2(n_853),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_840),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_914),
.B(n_915),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_957),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_939),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_917),
.B(n_938),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_L g989 ( 
.A1(n_847),
.A2(n_848),
.B(n_895),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_849),
.B(n_939),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_927),
.B(n_944),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_946),
.B(n_948),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_853),
.A2(n_852),
.B1(n_887),
.B2(n_935),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_872),
.B(n_875),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_889),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_949),
.B(n_959),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_893),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_864),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_861),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_875),
.B(n_942),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_930),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_909),
.B(n_880),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_882),
.B(n_848),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_940),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_883),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_897),
.B(n_846),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_930),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_947),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_878),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_897),
.B(n_876),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_888),
.Y(n_1011)
);

CKINVDCx8_ASAP7_75t_R g1012 ( 
.A(n_950),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_865),
.B(n_906),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_950),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_904),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_911),
.B(n_903),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_894),
.Y(n_1017)
);

CKINVDCx11_ASAP7_75t_R g1018 ( 
.A(n_839),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_878),
.B(n_913),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_898),
.B(n_905),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_945),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_873),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_908),
.B(n_896),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_884),
.A2(n_910),
.B(n_901),
.C(n_877),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_869),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_936),
.B(n_892),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_910),
.A2(n_928),
.B(n_937),
.C(n_924),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_862),
.A2(n_932),
.B1(n_953),
.B2(n_918),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_839),
.B(n_851),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_851),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_913),
.B(n_934),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_851),
.B(n_842),
.Y(n_1032)
);

BUFx4f_ASAP7_75t_SL g1033 ( 
.A(n_945),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_851),
.Y(n_1034)
);

AOI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_954),
.A2(n_907),
.B(n_859),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_926),
.B(n_945),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_936),
.B(n_892),
.Y(n_1037)
);

INVx2_ASAP7_75t_R g1038 ( 
.A(n_879),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_842),
.B(n_918),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_854),
.B(n_856),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_854),
.B(n_856),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_886),
.B(n_952),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_899),
.A2(n_874),
.B1(n_916),
.B2(n_941),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_899),
.A2(n_951),
.B(n_856),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_856),
.A2(n_891),
.B(n_902),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_891),
.A2(n_813),
.B(n_804),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_891),
.B(n_844),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_852),
.A2(n_833),
.B1(n_280),
.B2(n_300),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_849),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_840),
.Y(n_1050)
);

AO21x1_ASAP7_75t_L g1051 ( 
.A1(n_841),
.A2(n_775),
.B(n_729),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_855),
.B(n_929),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_956),
.B(n_841),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_919),
.B(n_933),
.Y(n_1054)
);

AO21x1_ASAP7_75t_L g1055 ( 
.A1(n_841),
.A2(n_775),
.B(n_729),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_956),
.B(n_841),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_864),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_864),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_956),
.B(n_841),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_947),
.B(n_900),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_943),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_947),
.B(n_900),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_900),
.B(n_929),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_919),
.B(n_933),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_921),
.A2(n_813),
.B(n_804),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_841),
.A2(n_925),
.B(n_958),
.C(n_729),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_956),
.B(n_841),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_956),
.B(n_841),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_956),
.A2(n_775),
.B(n_960),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_956),
.A2(n_775),
.B(n_753),
.C(n_749),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_920),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_841),
.A2(n_925),
.B(n_958),
.C(n_729),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_L g1073 ( 
.A(n_841),
.B(n_775),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_956),
.B(n_841),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_943),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_866),
.A2(n_770),
.B(n_729),
.C(n_775),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_956),
.B(n_867),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_922),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_956),
.A2(n_775),
.B1(n_770),
.B2(n_841),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_943),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_956),
.B(n_841),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_988),
.A2(n_971),
.B1(n_1079),
.B2(n_1025),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_990),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_1036),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1041),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_1034),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_SL g1087 ( 
.A1(n_971),
.A2(n_1079),
.B1(n_969),
.B2(n_1067),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_998),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_979),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_1040),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_984),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1053),
.A2(n_1081),
.B1(n_1056),
.B2(n_1059),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1026),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_964),
.B(n_1065),
.Y(n_1094)
);

BUFx8_ASAP7_75t_L g1095 ( 
.A(n_1014),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1053),
.A2(n_1081),
.B1(n_1056),
.B2(n_1059),
.Y(n_1096)
);

AO21x1_ASAP7_75t_L g1097 ( 
.A1(n_974),
.A2(n_1072),
.B(n_1066),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_1021),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_SL g1099 ( 
.A1(n_1067),
.A2(n_1068),
.B1(n_1074),
.B2(n_1013),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1069),
.A2(n_989),
.B1(n_1009),
.B2(n_1077),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1078),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1068),
.A2(n_1074),
.B1(n_1013),
.B2(n_1048),
.Y(n_1102)
);

BUFx8_ASAP7_75t_L g1103 ( 
.A(n_982),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_993),
.A2(n_961),
.B1(n_1064),
.B2(n_1054),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_972),
.A2(n_1047),
.B1(n_963),
.B2(n_1020),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

BUFx2_ASAP7_75t_R g1107 ( 
.A(n_1012),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_1033),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_997),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_1050),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1017),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_998),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_987),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1037),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_SL g1115 ( 
.A(n_1007),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_SL g1116 ( 
.A1(n_1010),
.A2(n_1016),
.B(n_1023),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_967),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_999),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1020),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1070),
.A2(n_962),
.B1(n_1010),
.B2(n_1016),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1004),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_983),
.B(n_966),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1046),
.A2(n_1051),
.B(n_1055),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_972),
.A2(n_1005),
.B1(n_981),
.B2(n_1003),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1005),
.A2(n_1006),
.B1(n_968),
.B2(n_978),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1022),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1037),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1049),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1006),
.A2(n_970),
.B1(n_1000),
.B2(n_996),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_1001),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_980),
.A2(n_992),
.B1(n_991),
.B2(n_985),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1057),
.A2(n_1058),
.B1(n_975),
.B2(n_1063),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_SL g1133 ( 
.A(n_976),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1015),
.B(n_1071),
.Y(n_1134)
);

AO22x1_ASAP7_75t_L g1135 ( 
.A1(n_1011),
.A2(n_994),
.B1(n_1002),
.B2(n_1015),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_977),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1019),
.A2(n_1031),
.B1(n_1002),
.B2(n_1080),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_1035),
.A2(n_1045),
.B(n_1044),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1052),
.A2(n_986),
.B1(n_1075),
.B2(n_1061),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1076),
.A2(n_1042),
.B(n_1024),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1028),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1027),
.A2(n_1044),
.B(n_1035),
.Y(n_1142)
);

OA21x2_ASAP7_75t_L g1143 ( 
.A1(n_1043),
.A2(n_1028),
.B(n_1038),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1032),
.B(n_1039),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1060),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1034),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1052),
.A2(n_1062),
.B1(n_1060),
.B2(n_1008),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

OAI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_1039),
.A2(n_1032),
.B(n_1029),
.Y(n_1149)
);

BUFx4f_ASAP7_75t_SL g1150 ( 
.A(n_973),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1030),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1030),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1048),
.A2(n_833),
.B1(n_857),
.B2(n_988),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_965),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_987),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_965),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1018),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_965),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_965),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_965),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_965),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1041),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_988),
.A2(n_833),
.B1(n_280),
.B2(n_300),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_1007),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1041),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_965),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_987),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_965),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1048),
.A2(n_833),
.B1(n_857),
.B2(n_988),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_R g1171 ( 
.A(n_984),
.B(n_592),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1033),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_965),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1077),
.B(n_981),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_965),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1073),
.A2(n_770),
.B(n_729),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_SL g1177 ( 
.A1(n_974),
.A2(n_1056),
.B(n_1053),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_988),
.A2(n_833),
.B1(n_280),
.B2(n_300),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1018),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1018),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_965),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1122),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1138),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1140),
.A2(n_1094),
.B(n_1123),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1083),
.B(n_1174),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1138),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1093),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1085),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1093),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1099),
.B(n_1131),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1113),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1155),
.B(n_1168),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1138),
.Y(n_1193)
);

BUFx2_ASAP7_75t_R g1194 ( 
.A(n_1084),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1163),
.B(n_1166),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1156),
.B(n_1090),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1134),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1128),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1156),
.B(n_1090),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1163),
.B(n_1166),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1114),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1127),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1118),
.Y(n_1203)
);

INVxp33_ASAP7_75t_L g1204 ( 
.A(n_1171),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1121),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1116),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1177),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1087),
.B(n_1082),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1177),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_1092),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1096),
.B(n_1141),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1124),
.B(n_1100),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1143),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1119),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1101),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1084),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1154),
.B(n_1157),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1159),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1160),
.B(n_1161),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1162),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1167),
.Y(n_1221)
);

NAND4xp25_ASAP7_75t_L g1222 ( 
.A(n_1176),
.B(n_1120),
.C(n_1117),
.D(n_1102),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1169),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1115),
.B(n_1165),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1173),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1175),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1181),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1106),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1109),
.B(n_1142),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1111),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1097),
.A2(n_1126),
.B(n_1139),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1143),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1105),
.A2(n_1125),
.B(n_1148),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1088),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1112),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_1170),
.B(n_1153),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1135),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1137),
.B(n_1104),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1091),
.B(n_1107),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1103),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1195),
.B(n_1180),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1206),
.B(n_1145),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1203),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1203),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1206),
.B(n_1136),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1205),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1208),
.A2(n_1178),
.B1(n_1164),
.B2(n_1133),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1232),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1229),
.Y(n_1250)
);

AOI221xp5_ASAP7_75t_L g1251 ( 
.A1(n_1208),
.A2(n_1133),
.B1(n_1179),
.B2(n_1158),
.C(n_1180),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1210),
.B(n_1103),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1229),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1211),
.B(n_1089),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1182),
.B(n_1179),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1211),
.B(n_1146),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1195),
.B(n_1158),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1184),
.A2(n_1147),
.B(n_1086),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1187),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1188),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1204),
.B(n_1091),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1233),
.A2(n_1149),
.B(n_1144),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1187),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1189),
.Y(n_1264)
);

CKINVDCx6p67_ASAP7_75t_R g1265 ( 
.A(n_1216),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1200),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1196),
.B(n_1152),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1200),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1185),
.B(n_1152),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1196),
.B(n_1132),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1253),
.B(n_1199),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1251),
.B(n_1222),
.C(n_1190),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1248),
.A2(n_1237),
.B1(n_1212),
.B2(n_1238),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1253),
.B(n_1199),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1266),
.B(n_1191),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1266),
.B(n_1197),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1250),
.B(n_1188),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1248),
.A2(n_1237),
.B1(n_1238),
.B2(n_1234),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1268),
.B(n_1192),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1268),
.B(n_1198),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1251),
.B(n_1209),
.C(n_1207),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1256),
.B(n_1235),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1252),
.A2(n_1207),
.B1(n_1209),
.B2(n_1237),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1250),
.B(n_1189),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_L g1285 ( 
.A(n_1269),
.B(n_1230),
.C(n_1227),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1254),
.B(n_1236),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1254),
.B(n_1215),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1252),
.B(n_1186),
.C(n_1193),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1249),
.A2(n_1220),
.B1(n_1225),
.B2(n_1221),
.C(n_1226),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1242),
.A2(n_1239),
.B1(n_1151),
.B2(n_1241),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1255),
.B(n_1215),
.Y(n_1291)
);

OAI221xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1270),
.A2(n_1213),
.B1(n_1183),
.B2(n_1193),
.C(n_1186),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1259),
.B(n_1183),
.C(n_1186),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1258),
.A2(n_1213),
.B(n_1232),
.Y(n_1294)
);

NAND2x1_ASAP7_75t_L g1295 ( 
.A(n_1246),
.B(n_1201),
.Y(n_1295)
);

AOI21xp33_ASAP7_75t_L g1296 ( 
.A1(n_1262),
.A2(n_1231),
.B(n_1184),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1267),
.B(n_1202),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1259),
.B(n_1202),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1263),
.B(n_1193),
.C(n_1183),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1267),
.B(n_1214),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1261),
.A2(n_1240),
.B(n_1224),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1264),
.B(n_1217),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1264),
.B(n_1219),
.Y(n_1303)
);

OAI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1257),
.A2(n_1225),
.B1(n_1223),
.B2(n_1221),
.C(n_1228),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1244),
.B(n_1232),
.C(n_1218),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1305),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1295),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1305),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1293),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1298),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1272),
.A2(n_1243),
.B(n_1246),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1292),
.B(n_1243),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1277),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1289),
.B(n_1244),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1293),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1272),
.A2(n_1243),
.B(n_1246),
.Y(n_1317)
);

NAND3x1_ASAP7_75t_SL g1318 ( 
.A(n_1294),
.B(n_1265),
.C(n_1194),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1299),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1299),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1285),
.B(n_1245),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1284),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1302),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1285),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1303),
.B(n_1245),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1283),
.B(n_1247),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1280),
.B(n_1260),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1277),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1287),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1304),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1288),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1327),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1314),
.B(n_1297),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1330),
.B(n_1275),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1306),
.B(n_1286),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1321),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1282),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1308),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1308),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1314),
.B(n_1300),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1321),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1324),
.B(n_1291),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1315),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1307),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1314),
.B(n_1300),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1330),
.B(n_1279),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1315),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1307),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1322),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1322),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1328),
.B(n_1257),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1307),
.B(n_1288),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1330),
.B(n_1265),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1328),
.B(n_1312),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1324),
.B(n_1247),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1325),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1308),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1325),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_L g1359 ( 
.A(n_1319),
.B(n_1281),
.C(n_1296),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1326),
.B(n_1276),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1310),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1310),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1310),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1361),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1365)
);

INVxp67_ASAP7_75t_SL g1366 ( 
.A(n_1359),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1337),
.B(n_1326),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1343),
.B(n_1308),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1343),
.A2(n_1331),
.B(n_1319),
.C(n_1316),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1347),
.B(n_1329),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1347),
.B(n_1329),
.Y(n_1371)
);

BUFx2_ASAP7_75t_R g1372 ( 
.A(n_1337),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1360),
.B(n_1329),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1334),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1360),
.B(n_1309),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1338),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1352),
.B(n_1331),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1361),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1338),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1338),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1359),
.B(n_1336),
.Y(n_1382)
);

NOR2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1339),
.B(n_1265),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_1357),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1339),
.A2(n_1319),
.B(n_1316),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1362),
.Y(n_1386)
);

OAI32xp33_ASAP7_75t_L g1387 ( 
.A1(n_1357),
.A2(n_1331),
.A3(n_1309),
.B1(n_1320),
.B2(n_1316),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1336),
.B(n_1309),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1341),
.B(n_1309),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1351),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1341),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1362),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1332),
.B(n_1316),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1355),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1363),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1353),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1333),
.B(n_1312),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1332),
.B(n_1320),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1352),
.Y(n_1399)
);

AOI32xp33_ASAP7_75t_L g1400 ( 
.A1(n_1342),
.A2(n_1331),
.A3(n_1320),
.B1(n_1313),
.B2(n_1273),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1363),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1351),
.B(n_1216),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1334),
.A2(n_1313),
.B1(n_1320),
.B2(n_1317),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1349),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1344),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1323),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1364),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1364),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1383),
.B(n_1352),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1379),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1383),
.B(n_1352),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1372),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1378),
.B(n_1333),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1387),
.A2(n_1294),
.B1(n_1311),
.B2(n_1317),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1378),
.B(n_1340),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1387),
.A2(n_1369),
.B(n_1382),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1391),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1378),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1374),
.B(n_1356),
.Y(n_1421)
);

NOR2x1_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1301),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1386),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1367),
.B(n_1356),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1386),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1405),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1405),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1358),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1394),
.B(n_1358),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1392),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1397),
.B(n_1340),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_1345),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1392),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1376),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1396),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1399),
.B(n_1345),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1395),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1395),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1399),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1370),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1401),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1436),
.B(n_1373),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1407),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_1402),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1407),
.Y(n_1446)
);

OAI221xp5_ASAP7_75t_L g1447 ( 
.A1(n_1417),
.A2(n_1400),
.B1(n_1389),
.B2(n_1388),
.C(n_1398),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1411),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1408),
.Y(n_1449)
);

AO22x1_ASAP7_75t_L g1450 ( 
.A1(n_1422),
.A2(n_1384),
.B1(n_1393),
.B2(n_1344),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1411),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1419),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1440),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1390),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1415),
.A2(n_1403),
.B1(n_1346),
.B2(n_1278),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1440),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1408),
.A2(n_1371),
.B(n_1355),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1420),
.A2(n_1406),
.B(n_1380),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1419),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1436),
.B(n_1301),
.Y(n_1460)
);

AOI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1429),
.A2(n_1381),
.B1(n_1380),
.B2(n_1376),
.C(n_1401),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1424),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1418),
.B(n_1390),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1416),
.B(n_1365),
.Y(n_1464)
);

NOR4xp25_ASAP7_75t_SL g1465 ( 
.A(n_1424),
.B(n_1404),
.C(n_1318),
.D(n_1350),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1423),
.B(n_1346),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1420),
.A2(n_1441),
.B(n_1423),
.C(n_1421),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1444),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1427),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1446),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1453),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1420),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1456),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1460),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1448),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1451),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1457),
.B(n_1428),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1455),
.A2(n_1435),
.B1(n_1412),
.B2(n_1410),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1450),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1445),
.B(n_1428),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1445),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1463),
.B(n_1425),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1480),
.A2(n_1447),
.B(n_1465),
.Y(n_1489)
);

NAND4xp75_ASAP7_75t_L g1490 ( 
.A(n_1477),
.B(n_1443),
.C(n_1458),
.D(n_1461),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1485),
.A2(n_1468),
.B1(n_1484),
.B2(n_1487),
.C(n_1483),
.Y(n_1491)
);

AOI211xp5_ASAP7_75t_L g1492 ( 
.A1(n_1485),
.A2(n_1412),
.B(n_1410),
.C(n_1452),
.Y(n_1492)
);

AOI32xp33_ASAP7_75t_L g1493 ( 
.A1(n_1477),
.A2(n_1410),
.A3(n_1412),
.B1(n_1462),
.B2(n_1459),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1473),
.B(n_1464),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1486),
.B(n_1464),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1469),
.B(n_1430),
.Y(n_1496)
);

OAI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1473),
.A2(n_1437),
.B(n_1409),
.Y(n_1497)
);

AOI211x1_ASAP7_75t_L g1498 ( 
.A1(n_1474),
.A2(n_1467),
.B(n_1437),
.C(n_1433),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1469),
.A2(n_1431),
.B(n_1426),
.Y(n_1499)
);

NAND4xp25_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1476),
.C(n_1479),
.D(n_1488),
.Y(n_1500)
);

AOI211xp5_ASAP7_75t_L g1501 ( 
.A1(n_1491),
.A2(n_1478),
.B(n_1475),
.C(n_1479),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1489),
.B(n_1481),
.C(n_1470),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1490),
.A2(n_1476),
.B1(n_1488),
.B2(n_1435),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1494),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1496),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1495),
.B(n_1150),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1508)
);

AO22x2_ASAP7_75t_L g1509 ( 
.A1(n_1499),
.A2(n_1482),
.B1(n_1481),
.B2(n_1438),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1492),
.B(n_1432),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1501),
.A2(n_1482),
.B(n_1497),
.C(n_1442),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_SL g1512 ( 
.A(n_1503),
.B(n_1493),
.C(n_1172),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1504),
.B(n_1506),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1432),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1507),
.A2(n_1442),
.B(n_1439),
.C(n_1431),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1514),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1515),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1511),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1512),
.A2(n_1502),
.B1(n_1509),
.B2(n_1510),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1513),
.A2(n_1509),
.B1(n_1508),
.B2(n_1381),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1514),
.Y(n_1521)
);

AO21x1_ASAP7_75t_L g1522 ( 
.A1(n_1517),
.A2(n_1438),
.B(n_1434),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1516),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1518),
.A2(n_1439),
.B1(n_1434),
.B2(n_1404),
.C(n_1433),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1521),
.Y(n_1525)
);

XNOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1519),
.B(n_1108),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1526),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1523),
.B(n_1520),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1525),
.B(n_1344),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1529),
.Y(n_1530)
);

NOR2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1530),
.B(n_1527),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1531),
.B(n_1528),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1531),
.Y(n_1533)
);

AOI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1532),
.A2(n_1522),
.B(n_1524),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1533),
.A2(n_1172),
.B1(n_1108),
.B2(n_1348),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1535),
.A2(n_1534),
.B1(n_1110),
.B2(n_1130),
.C1(n_1095),
.C2(n_1098),
.Y(n_1536)
);

AOI222xp33_ASAP7_75t_L g1537 ( 
.A1(n_1535),
.A2(n_1130),
.B1(n_1098),
.B2(n_1133),
.C1(n_1110),
.C2(n_1348),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1537),
.B(n_1365),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1538),
.A2(n_1536),
.B1(n_1110),
.B2(n_1098),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_R g1540 ( 
.A1(n_1539),
.A2(n_1095),
.B1(n_1348),
.B2(n_1318),
.C(n_1377),
.Y(n_1540)
);

AOI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1540),
.A2(n_1095),
.B(n_1377),
.C(n_1290),
.Y(n_1541)
);


endmodule