module fake_jpeg_24544_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_49),
.B1(n_21),
.B2(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_63),
.B1(n_65),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_29),
.B2(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_20),
.B1(n_27),
.B2(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_73),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_83),
.B1(n_84),
.B2(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_22),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_21),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_16),
.B1(n_19),
.B2(n_10),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_63),
.B1(n_61),
.B2(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_44),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_92),
.C(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_91),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_88),
.B1(n_69),
.B2(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_105),
.B1(n_108),
.B2(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_59),
.B(n_48),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_105),
.B(n_92),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_19),
.B1(n_78),
.B2(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_82),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_50),
.B1(n_55),
.B2(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_89),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_73),
.B1(n_75),
.B2(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_123),
.B1(n_137),
.B2(n_1),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_74),
.B1(n_70),
.B2(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_131),
.B1(n_22),
.B2(n_24),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_76),
.B(n_71),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_135),
.B(n_94),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_62),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_62),
.B1(n_76),
.B2(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_142),
.Y(n_168)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_148),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_104),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_0),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_2),
.B(n_3),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_30),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_95),
.B1(n_101),
.B2(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_101),
.B1(n_91),
.B2(n_100),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_31),
.B1(n_24),
.B2(n_22),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_7),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_114),
.C(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_0),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_0),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_126),
.B1(n_131),
.B2(n_127),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_8),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_9),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_115),
.B1(n_114),
.B2(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_176),
.C(n_186),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_172),
.B1(n_181),
.B2(n_164),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_178),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_115),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_183),
.B(n_143),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_117),
.B1(n_138),
.B2(n_133),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_117),
.C(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_7),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_142),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_196),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_170),
.B(n_171),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_194),
.B1(n_199),
.B2(n_183),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_148),
.B1(n_164),
.B2(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_166),
.B1(n_187),
.B2(n_175),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_140),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_144),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_150),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_173),
.C(n_177),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_156),
.B1(n_161),
.B2(n_4),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_9),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_207),
.Y(n_215)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_185),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_6),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_167),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_223),
.B1(n_225),
.B2(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_15),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_190),
.C(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_221),
.C(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_199),
.B1(n_195),
.B2(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_218),
.B1(n_225),
.B2(n_226),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_194),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_215),
.C(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_215),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_197),
.C(n_10),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_11),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_247),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_228),
.C(n_234),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_238),
.B1(n_237),
.B2(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_248),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_256),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_227),
.B1(n_210),
.B2(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_212),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_11),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_5),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_241),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_258),
.C(n_253),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

OAI31xp67_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_259),
.A3(n_3),
.B(n_4),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_5),
.B(n_13),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_15),
.C(n_270),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_271),
.B(n_267),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_276),
.B1(n_2),
.B2(n_3),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_263),
.B(n_3),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_2),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_273),
.Y(n_280)
);


endmodule