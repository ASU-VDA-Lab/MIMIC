module fake_jpeg_13225_n_350 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_43),
.Y(n_90)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_56),
.Y(n_92)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_59),
.Y(n_97)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_8),
.B(n_13),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_31),
.Y(n_95)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_23),
.B1(n_36),
.B2(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_91),
.B1(n_93),
.B2(n_101),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_30),
.B1(n_41),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_86),
.B1(n_113),
.B2(n_37),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_75),
.B(n_79),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_42),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_41),
.B1(n_33),
.B2(n_32),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_100),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_22),
.B1(n_38),
.B2(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_38),
.B1(n_31),
.B2(n_27),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_R g150 ( 
.A(n_95),
.B(n_37),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_26),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_16),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_25),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_54),
.B1(n_64),
.B2(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_33),
.B1(n_34),
.B2(n_29),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_25),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_60),
.B(n_27),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_38),
.B1(n_24),
.B2(n_41),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_110),
.B1(n_21),
.B2(n_2),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_41),
.B1(n_30),
.B2(n_32),
.Y(n_112)
);

OA22x2_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_21),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_33),
.B1(n_34),
.B2(n_29),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_12),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_125),
.A2(n_152),
.B1(n_153),
.B2(n_113),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_128),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_0),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_143),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_37),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_108),
.C(n_97),
.Y(n_170)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_144),
.Y(n_167)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_0),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_80),
.Y(n_144)
);

AND2x4_ASAP7_75t_SL g145 ( 
.A(n_79),
.B(n_37),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_117),
.Y(n_156)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_82),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_112),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_37),
.B1(n_21),
.B2(n_9),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_151),
.A2(n_154),
.B1(n_100),
.B2(n_83),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_95),
.A2(n_21),
.B1(n_15),
.B2(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_155),
.A2(n_178),
.B1(n_153),
.B2(n_151),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_120),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_92),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_75),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_95),
.B1(n_111),
.B2(n_86),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_190),
.B1(n_156),
.B2(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_179),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_172),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_111),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_180),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_97),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_188),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_186),
.Y(n_210)
);

O2A1O1Ixp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_112),
.B(n_118),
.C(n_82),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_119),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_119),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_187),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_115),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_189),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_104),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_133),
.B(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_145),
.C(n_127),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_204),
.C(n_156),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_121),
.B1(n_144),
.B2(n_109),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_109),
.B1(n_160),
.B2(n_76),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_154),
.B1(n_125),
.B2(n_131),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_221),
.B1(n_203),
.B2(n_216),
.Y(n_228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_150),
.B(n_145),
.C(n_127),
.D(n_129),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_198),
.A2(n_202),
.B(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_222),
.B(n_182),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_123),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_217),
.B1(n_156),
.B2(n_177),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_213),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_153),
.B(n_129),
.C(n_112),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_215),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_140),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_158),
.A2(n_190),
.B1(n_168),
.B2(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_134),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_175),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_153),
.B(n_84),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_159),
.B(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_158),
.A2(n_167),
.B1(n_187),
.B2(n_181),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_159),
.B(n_124),
.C(n_130),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_242),
.C(n_203),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_231),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_244),
.B(n_246),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_205),
.B1(n_208),
.B2(n_211),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_194),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_234),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_199),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_243),
.B1(n_196),
.B2(n_221),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_245),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_163),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_217),
.A2(n_169),
.B1(n_94),
.B2(n_96),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_166),
.B(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_166),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_198),
.B(n_202),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_239),
.B(n_227),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_254),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_258),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_243),
.B1(n_225),
.B2(n_226),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_193),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_262),
.C(n_263),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_259),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_236),
.B(n_235),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_248),
.C(n_241),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_233),
.B1(n_214),
.B2(n_160),
.Y(n_283)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_212),
.B1(n_220),
.B2(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_200),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_270),
.C(n_235),
.Y(n_280)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_269),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_191),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_289),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_225),
.B(n_244),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_284),
.B(n_269),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_231),
.A3(n_226),
.B1(n_225),
.B2(n_212),
.C1(n_240),
.C2(n_232),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_267),
.C(n_251),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_287),
.B(n_288),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_233),
.C(n_215),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_266),
.B1(n_252),
.B2(n_103),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_84),
.B(n_147),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_174),
.B(n_87),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_174),
.B(n_87),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_251),
.CI(n_260),
.CON(n_291),
.SN(n_291)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_302),
.B(n_306),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_295),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_260),
.C(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_265),
.B(n_263),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_257),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_277),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_287),
.B1(n_94),
.B2(n_185),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_286),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_278),
.A2(n_281),
.B(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_313),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_281),
.B1(n_282),
.B2(n_273),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_249),
.B1(n_288),
.B2(n_265),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_303),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_265),
.B1(n_273),
.B2(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_317),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_304),
.B1(n_296),
.B2(n_291),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_254),
.B1(n_185),
.B2(n_94),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_298),
.Y(n_324)
);

AOI21x1_ASAP7_75t_SL g321 ( 
.A1(n_307),
.A2(n_302),
.B(n_306),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_309),
.B(n_314),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_295),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_323),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_291),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_313),
.B1(n_315),
.B2(n_311),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_141),
.C(n_149),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_96),
.Y(n_334)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_308),
.B(n_320),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_333),
.B(n_327),
.Y(n_338)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_76),
.B(n_15),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_1),
.C(n_2),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_338),
.A2(n_334),
.B(n_4),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_81),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_340),
.B(n_337),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_344),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_345),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_2),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_347),
.A2(n_346),
.B1(n_343),
.B2(n_342),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_348),
.Y(n_350)
);


endmodule