module fake_aes_12073_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx4_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_2), .B(n_1), .Y(n_4) );
O2A1O1Ixp33_ASAP7_75t_SL g5 ( .A1(n_4), .A2(n_0), .B(n_1), .C(n_2), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
NOR2x1p5_ASAP7_75t_L g7 ( .A(n_6), .B(n_3), .Y(n_7) );
AOI222xp33_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_0), .B1(n_1), .B2(n_4), .C1(n_3), .C2(n_5), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
OAI22xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_11), .B1(n_7), .B2(n_8), .Y(n_13) );
endmodule