module real_aes_6390_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g257 ( .A1(n_0), .A2(n_258), .B(n_259), .C(n_262), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_1), .B(n_246), .Y(n_263) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_91), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g459 ( .A(n_2), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_3), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_4), .A2(n_135), .B(n_138), .C(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_5), .A2(n_130), .B(n_577), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_6), .A2(n_130), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_7), .B(n_246), .Y(n_583) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_8), .A2(n_165), .B(n_202), .Y(n_201) );
AND2x6_ASAP7_75t_L g135 ( .A(n_9), .B(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_10), .A2(n_135), .B(n_138), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g521 ( .A(n_11), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_12), .B(n_41), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_13), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_13), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_14), .B(n_222), .Y(n_555) );
INVx1_ASAP7_75t_L g156 ( .A(n_15), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_16), .B(n_174), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_17), .A2(n_175), .B(n_539), .C(n_541), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_18), .B(n_246), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_19), .B(n_150), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_20), .A2(n_138), .B(n_141), .C(n_149), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_21), .A2(n_210), .B(n_261), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_22), .B(n_222), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_23), .A2(n_57), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_23), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_24), .B(n_222), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g568 ( .A(n_25), .Y(n_568) );
INVx1_ASAP7_75t_L g493 ( .A(n_26), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_27), .A2(n_138), .B(n_149), .C(n_205), .Y(n_204) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_28), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_29), .Y(n_551) );
INVx1_ASAP7_75t_L g509 ( .A(n_30), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_31), .A2(n_130), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_33), .A2(n_178), .B(n_187), .C(n_189), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_34), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_35), .A2(n_261), .B(n_580), .C(n_582), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_36), .A2(n_105), .B1(n_114), .B2(n_766), .Y(n_104) );
INVxp67_ASAP7_75t_L g510 ( .A(n_37), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_38), .B(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_39), .A2(n_138), .B(n_149), .C(n_492), .Y(n_491) );
CKINVDCx14_ASAP7_75t_R g578 ( .A(n_40), .Y(n_578) );
INVx1_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_42), .A2(n_262), .B(n_519), .C(n_520), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_43), .B(n_129), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_44), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_45), .B(n_174), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_46), .B(n_130), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_47), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_48), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_49), .A2(n_178), .B(n_187), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_50), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g260 ( .A(n_51), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_52), .A2(n_447), .B1(n_448), .B2(n_451), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_52), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_53), .A2(n_466), .B1(n_467), .B2(n_476), .C1(n_756), .C2(n_760), .Y(n_465) );
INVx1_ASAP7_75t_L g232 ( .A(n_54), .Y(n_232) );
INVx1_ASAP7_75t_L g527 ( .A(n_55), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_56), .B(n_130), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_57), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_58), .Y(n_158) );
CKINVDCx14_ASAP7_75t_R g517 ( .A(n_59), .Y(n_517) );
INVx1_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_61), .B(n_130), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_62), .B(n_246), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_63), .A2(n_148), .B(n_171), .C(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g155 ( .A(n_64), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_65), .A2(n_103), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_65), .Y(n_473) );
INVx1_ASAP7_75t_SL g581 ( .A(n_66), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_67), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_68), .B(n_174), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_69), .B(n_246), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_70), .B(n_175), .Y(n_220) );
INVx1_ASAP7_75t_L g571 ( .A(n_71), .Y(n_571) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_72), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_73), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_74), .A2(n_138), .B(n_169), .C(n_178), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_75), .Y(n_241) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_77), .A2(n_130), .B(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_78), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_79), .A2(n_130), .B(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_80), .A2(n_129), .B(n_505), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_81), .Y(n_490) );
INVx1_ASAP7_75t_L g537 ( .A(n_82), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_83), .B(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_84), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_85), .A2(n_130), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g540 ( .A(n_86), .Y(n_540) );
INVx2_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx1_ASAP7_75t_L g554 ( .A(n_88), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_89), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_90), .B(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g456 ( .A(n_91), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g479 ( .A(n_91), .B(n_458), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_91), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_92), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_92), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_93), .A2(n_138), .B(n_178), .C(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_94), .B(n_130), .Y(n_185) );
INVx1_ASAP7_75t_L g190 ( .A(n_95), .Y(n_190) );
INVxp67_ASAP7_75t_L g244 ( .A(n_96), .Y(n_244) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_97), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_97), .B(n_165), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g170 ( .A(n_99), .Y(n_170) );
INVx1_ASAP7_75t_L g216 ( .A(n_100), .Y(n_216) );
INVx2_ASAP7_75t_L g530 ( .A(n_101), .Y(n_530) );
AND2x2_ASAP7_75t_L g234 ( .A(n_102), .B(n_152), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_103), .Y(n_472) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g766 ( .A(n_106), .Y(n_766) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_117), .B(n_464), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g765 ( .A(n_116), .Y(n_765) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_453), .B(n_461), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_445), .B1(n_446), .B2(n_452), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_120), .A2(n_483), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g452 ( .A(n_121), .Y(n_452) );
AND3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_349), .C(n_406), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_294), .C(n_330), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_196), .B(n_248), .C(n_281), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g251 ( .A(n_126), .B(n_252), .Y(n_251) );
INVx5_ASAP7_75t_L g280 ( .A(n_126), .Y(n_280) );
AND2x2_ASAP7_75t_L g353 ( .A(n_126), .B(n_269), .Y(n_353) );
AND2x2_ASAP7_75t_L g391 ( .A(n_126), .B(n_297), .Y(n_391) );
AND2x2_ASAP7_75t_L g411 ( .A(n_126), .B(n_253), .Y(n_411) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_157), .Y(n_126) );
AOI21xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_137), .B(n_150), .Y(n_127) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_131), .B(n_135), .Y(n_217) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_134), .Y(n_144) );
INVx3_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_134), .Y(n_222) );
BUFx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx4_ASAP7_75t_SL g179 ( .A(n_135), .Y(n_179) );
INVx5_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
BUFx3_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_147), .Y(n_141) );
INVx2_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_146), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_146), .A2(n_192), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g553 ( .A1(n_146), .A2(n_554), .B(n_555), .C(n_556), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_146), .A2(n_556), .B(n_571), .C(n_572), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_147), .A2(n_174), .B(n_493), .C(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_148), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_151), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_152), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_152), .A2(n_229), .B(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_152), .A2(n_217), .B(n_490), .C(n_491), .Y(n_489) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_152), .A2(n_515), .B(n_522), .Y(n_514) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g166 ( .A(n_153), .B(n_154), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_159), .A2(n_550), .B(n_557), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_160), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_183), .Y(n_160) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_161), .Y(n_292) );
AND2x2_ASAP7_75t_L g306 ( .A(n_161), .B(n_252), .Y(n_306) );
INVx1_ASAP7_75t_L g329 ( .A(n_161), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_161), .B(n_280), .Y(n_368) );
OR2x2_ASAP7_75t_L g405 ( .A(n_161), .B(n_250), .Y(n_405) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_162), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_162), .B(n_253), .Y(n_348) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g269 ( .A(n_163), .B(n_253), .Y(n_269) );
BUFx2_ASAP7_75t_L g297 ( .A(n_163), .Y(n_297) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_181), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_164), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_164), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_164), .A2(n_215), .B(n_223), .Y(n_214) );
INVx3_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_164), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_164), .B(n_558), .Y(n_557) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_164), .A2(n_567), .B(n_573), .Y(n_566) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_165), .A2(n_203), .B(n_204), .Y(n_202) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_165), .Y(n_238) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_173), .C(n_176), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_172), .A2(n_174), .B1(n_509), .B2(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_172), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_172), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_174), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g258 ( .A(n_174), .Y(n_258) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_175), .B(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g582 ( .A(n_177), .Y(n_582) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_179), .A2(n_188), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_179), .A2(n_188), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_179), .A2(n_188), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_179), .A2(n_188), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g526 ( .A1(n_179), .A2(n_188), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_179), .A2(n_188), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g577 ( .A1(n_179), .A2(n_188), .B(n_578), .C(n_579), .Y(n_577) );
INVx5_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
BUFx2_ASAP7_75t_L g273 ( .A(n_183), .Y(n_273) );
AND2x2_ASAP7_75t_L g430 ( .A(n_183), .B(n_284), .Y(n_430) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_194), .Y(n_183) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g262 ( .A(n_193), .Y(n_262) );
INVx1_ASAP7_75t_L g541 ( .A(n_193), .Y(n_541) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_235), .Y(n_197) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_198), .A2(n_331), .B1(n_338), .B2(n_339), .C(n_342), .Y(n_330) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_212), .Y(n_198) );
AND2x2_ASAP7_75t_L g236 ( .A(n_199), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_199), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g265 ( .A(n_200), .B(n_213), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_200), .B(n_214), .Y(n_275) );
OR2x2_ASAP7_75t_L g286 ( .A(n_200), .B(n_237), .Y(n_286) );
AND2x2_ASAP7_75t_L g289 ( .A(n_200), .B(n_277), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_200), .B(n_226), .Y(n_305) );
OR2x2_ASAP7_75t_L g321 ( .A(n_200), .B(n_214), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_200), .B(n_237), .Y(n_383) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_201), .B(n_226), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_201), .B(n_214), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B(n_209), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g299 ( .A(n_212), .B(n_286), .Y(n_299) );
INVx2_ASAP7_75t_L g325 ( .A(n_212), .Y(n_325) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
AND2x2_ASAP7_75t_L g247 ( .A(n_213), .B(n_227), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_213), .B(n_237), .Y(n_304) );
OR2x2_ASAP7_75t_L g315 ( .A(n_213), .B(n_227), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_213), .B(n_277), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_213), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_407) );
INVx5_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_214), .B(n_237), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_217), .A2(n_551), .B(n_552), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_217), .A2(n_568), .B(n_569), .Y(n_567) );
INVx4_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
INVx2_ASAP7_75t_L g519 ( .A(n_222), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g502 ( .A(n_225), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_226), .B(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_226), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g293 ( .A(n_226), .B(n_265), .Y(n_293) );
OR2x2_ASAP7_75t_L g337 ( .A(n_226), .B(n_237), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_226), .B(n_289), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_226), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_226), .B(n_403), .Y(n_402) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_227), .B(n_236), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_227), .A2(n_271), .B(n_274), .C(n_278), .Y(n_270) );
OR2x2_ASAP7_75t_L g308 ( .A(n_227), .B(n_304), .Y(n_308) );
OR2x2_ASAP7_75t_L g344 ( .A(n_227), .B(n_286), .Y(n_344) );
OAI311xp33_ASAP7_75t_L g350 ( .A1(n_227), .A2(n_289), .A3(n_351), .B1(n_354), .C1(n_361), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_227), .B(n_237), .Y(n_401) );
AND2x2_ASAP7_75t_L g409 ( .A(n_227), .B(n_264), .Y(n_409) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_227), .Y(n_427) );
AND2x2_ASAP7_75t_L g444 ( .A(n_227), .B(n_265), .Y(n_444) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_247), .Y(n_235) );
AND2x2_ASAP7_75t_L g272 ( .A(n_236), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g428 ( .A(n_236), .Y(n_428) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g277 ( .A(n_237), .Y(n_277) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
INVxp67_ASAP7_75t_L g359 ( .A(n_237), .Y(n_359) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_245), .Y(n_237) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_238), .A2(n_525), .B(n_531), .Y(n_524) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_238), .A2(n_535), .B(n_542), .Y(n_534) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_238), .A2(n_576), .B(n_583), .Y(n_575) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_246), .A2(n_254), .B(n_263), .Y(n_253) );
AND2x2_ASAP7_75t_L g437 ( .A(n_247), .B(n_285), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_264), .B1(n_266), .B2(n_267), .C(n_270), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_250), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g290 ( .A(n_250), .B(n_280), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_250), .B(n_252), .Y(n_298) );
OR2x2_ASAP7_75t_L g310 ( .A(n_250), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_250), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g352 ( .A(n_250), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_250), .Y(n_372) );
AND2x2_ASAP7_75t_L g424 ( .A(n_250), .B(n_348), .Y(n_424) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_250), .A2(n_301), .A3(n_400), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_251), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g396 ( .A(n_251), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_251), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g284 ( .A(n_252), .B(n_280), .Y(n_284) );
INVx1_ASAP7_75t_L g371 ( .A(n_252), .Y(n_371) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g421 ( .A(n_253), .B(n_280), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_261), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g556 ( .A(n_262), .Y(n_556) );
INVx1_ASAP7_75t_SL g431 ( .A(n_264), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_265), .B(n_336), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_266), .A2(n_378), .B1(n_416), .B2(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_269), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_269), .B(n_290), .Y(n_443) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g413 ( .A(n_272), .B(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_273), .A2(n_332), .B(n_334), .Y(n_331) );
OR2x2_ASAP7_75t_L g339 ( .A(n_273), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g360 ( .A(n_273), .B(n_348), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_273), .B(n_371), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_273), .B(n_411), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g387 ( .A1(n_274), .A2(n_388), .B1(n_393), .B2(n_396), .C(n_397), .Y(n_387) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g364 ( .A(n_275), .B(n_337), .Y(n_364) );
INVx1_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
INVx2_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_280), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g347 ( .A(n_280), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g435 ( .A(n_280), .B(n_405), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B1(n_287), .B2(n_290), .C1(n_291), .C2(n_293), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_284), .A2(n_334), .B1(n_362), .B2(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_284), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OAI21xp33_ASAP7_75t_SL g322 ( .A1(n_293), .A2(n_323), .B(n_326), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_299), .B(n_300), .C(n_322), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_298), .A2(n_301), .B1(n_306), .B2(n_307), .C(n_309), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_298), .B(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g392 ( .A(n_298), .Y(n_392) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
AND2x2_ASAP7_75t_L g394 ( .A(n_303), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g311 ( .A(n_306), .Y(n_311) );
AND2x2_ASAP7_75t_L g317 ( .A(n_306), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_316), .B2(n_319), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_313), .B(n_325), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_314), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g414 ( .A(n_318), .Y(n_414) );
AND2x2_ASAP7_75t_L g433 ( .A(n_318), .B(n_348), .Y(n_433) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_325), .B(n_382), .Y(n_441) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_328), .B(n_396), .Y(n_439) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
BUFx2_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
OAI21xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_345), .B(n_347), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_365), .C(n_387), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_369), .B(n_373), .C(n_376), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_366), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp67_ASAP7_75t_SL g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g395 ( .A(n_375), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B(n_384), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g400 ( .A(n_378), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_402), .B2(n_404), .Y(n_397) );
INVx2_ASAP7_75t_SL g418 ( .A(n_405), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_422), .C(n_434), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_418), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_429), .B2(n_431), .C(n_432), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_423), .A2(n_435), .B(n_436), .C(n_438), .Y(n_434) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_442), .B2(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_452), .A2(n_477), .B1(n_480), .B2(n_482), .Y(n_476) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_456), .Y(n_463) );
NOR2x2_ASAP7_75t_L g762 ( .A(n_457), .B(n_481), .Y(n_762) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g480 ( .A(n_458), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_461), .B(n_465), .C(n_763), .Y(n_464) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_471), .Y(n_474) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g757 ( .A(n_478), .Y(n_757) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g759 ( .A(n_480), .Y(n_759) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
OR5x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_650), .C(n_714), .D(n_730), .E(n_745), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_485), .B(n_584), .C(n_611), .D(n_634), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_532), .B(n_543), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_497), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_SL g563 ( .A(n_488), .Y(n_563) );
AND2x4_ASAP7_75t_L g597 ( .A(n_488), .B(n_586), .Y(n_597) );
OR2x2_ASAP7_75t_L g607 ( .A(n_488), .B(n_565), .Y(n_607) );
OR2x2_ASAP7_75t_L g653 ( .A(n_488), .B(n_500), .Y(n_653) );
AND2x2_ASAP7_75t_L g667 ( .A(n_488), .B(n_564), .Y(n_667) );
AND2x2_ASAP7_75t_L g710 ( .A(n_488), .B(n_600), .Y(n_710) );
AND2x2_ASAP7_75t_L g717 ( .A(n_488), .B(n_575), .Y(n_717) );
AND2x2_ASAP7_75t_L g736 ( .A(n_488), .B(n_626), .Y(n_736) );
AND2x2_ASAP7_75t_L g754 ( .A(n_488), .B(n_596), .Y(n_754) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g719 ( .A(n_497), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_513), .Y(n_497) );
AND2x2_ASAP7_75t_L g629 ( .A(n_498), .B(n_564), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_498), .B(n_649), .Y(n_648) );
AOI32xp33_ASAP7_75t_L g662 ( .A1(n_498), .A2(n_663), .A3(n_666), .B1(n_668), .B2(n_672), .Y(n_662) );
AND2x2_ASAP7_75t_L g732 ( .A(n_498), .B(n_626), .Y(n_732) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g596 ( .A(n_500), .B(n_565), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_500), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g638 ( .A(n_500), .B(n_585), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_500), .B(n_717), .Y(n_716) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_503), .B(n_511), .Y(n_500) );
INVx1_ASAP7_75t_L g601 ( .A(n_501), .Y(n_601) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_504), .A2(n_512), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g603 ( .A(n_513), .B(n_547), .Y(n_603) );
AND2x2_ASAP7_75t_L g679 ( .A(n_513), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g751 ( .A(n_513), .Y(n_751) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
OR2x2_ASAP7_75t_L g546 ( .A(n_514), .B(n_524), .Y(n_546) );
AND2x2_ASAP7_75t_L g560 ( .A(n_514), .B(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_514), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g610 ( .A(n_514), .Y(n_610) );
AND2x2_ASAP7_75t_L g637 ( .A(n_514), .B(n_524), .Y(n_637) );
BUFx3_ASAP7_75t_L g640 ( .A(n_514), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_514), .B(n_615), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_514), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g591 ( .A(n_523), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_523), .B(n_589), .Y(n_609) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g620 ( .A(n_524), .B(n_534), .Y(n_620) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_524), .Y(n_633) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_533), .B(n_640), .Y(n_690) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_SL g561 ( .A(n_534), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_534), .B(n_609), .C(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g616 ( .A(n_534), .B(n_589), .Y(n_616) );
AND2x2_ASAP7_75t_L g636 ( .A(n_534), .B(n_589), .Y(n_636) );
AND2x2_ASAP7_75t_L g680 ( .A(n_534), .B(n_549), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_559), .B(n_562), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_547), .Y(n_544) );
AND2x2_ASAP7_75t_L g755 ( .A(n_545), .B(n_680), .Y(n_755) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_546), .A2(n_653), .B1(n_695), .B2(n_697), .Y(n_694) );
OR2x2_ASAP7_75t_L g701 ( .A(n_546), .B(n_616), .Y(n_701) );
OR2x2_ASAP7_75t_L g725 ( .A(n_546), .B(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_546), .B(n_645), .Y(n_738) );
AND2x2_ASAP7_75t_L g631 ( .A(n_547), .B(n_632), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_547), .A2(n_704), .B(n_719), .Y(n_718) );
AOI32xp33_ASAP7_75t_L g739 ( .A1(n_547), .A2(n_629), .A3(n_740), .B1(n_742), .B2(n_743), .Y(n_739) );
OR2x2_ASAP7_75t_L g750 ( .A(n_547), .B(n_751), .Y(n_750) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_548), .B(n_632), .Y(n_697) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g589 ( .A(n_549), .Y(n_589) );
AND2x2_ASAP7_75t_L g655 ( .A(n_549), .B(n_620), .Y(n_655) );
AND3x2_ASAP7_75t_L g664 ( .A(n_549), .B(n_560), .C(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g590 ( .A(n_561), .B(n_591), .Y(n_590) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_561), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_561), .B(n_589), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g585 ( .A(n_563), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g625 ( .A(n_563), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g643 ( .A(n_563), .B(n_575), .Y(n_643) );
AND2x2_ASAP7_75t_L g661 ( .A(n_563), .B(n_565), .Y(n_661) );
OR2x2_ASAP7_75t_L g675 ( .A(n_563), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g721 ( .A(n_563), .B(n_649), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_564), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_575), .Y(n_564) );
AND2x2_ASAP7_75t_L g622 ( .A(n_565), .B(n_600), .Y(n_622) );
OR2x2_ASAP7_75t_L g676 ( .A(n_565), .B(n_600), .Y(n_676) );
AND2x2_ASAP7_75t_L g729 ( .A(n_565), .B(n_586), .Y(n_729) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g627 ( .A(n_566), .Y(n_627) );
AND2x2_ASAP7_75t_L g649 ( .A(n_566), .B(n_575), .Y(n_649) );
INVx2_ASAP7_75t_L g586 ( .A(n_575), .Y(n_586) );
INVx1_ASAP7_75t_L g606 ( .A(n_575), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B(n_592), .C(n_604), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_585), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g748 ( .A(n_585), .Y(n_748) );
AND2x2_ASAP7_75t_L g626 ( .A(n_586), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_589), .B(n_590), .Y(n_598) );
INVx1_ASAP7_75t_L g683 ( .A(n_589), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_589), .B(n_610), .Y(n_707) );
AND2x2_ASAP7_75t_L g723 ( .A(n_589), .B(n_637), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_590), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g614 ( .A(n_591), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_595), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_596), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g621 ( .A(n_597), .B(n_622), .Y(n_621) );
AOI221xp5_ASAP7_75t_SL g686 ( .A1(n_597), .A2(n_639), .B1(n_687), .B2(n_692), .C(n_694), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_597), .B(n_660), .Y(n_693) );
INVx1_ASAP7_75t_L g753 ( .A(n_599), .Y(n_753) );
BUFx3_ASAP7_75t_L g660 ( .A(n_600), .Y(n_660) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_608), .Y(n_604) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_606), .B(n_660), .Y(n_713) );
INVx1_ASAP7_75t_L g670 ( .A(n_607), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_607), .B(n_660), .Y(n_671) );
INVxp67_ASAP7_75t_L g691 ( .A(n_609), .Y(n_691) );
AND2x2_ASAP7_75t_L g632 ( .A(n_610), .B(n_633), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_617), .B(n_621), .C(n_623), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_SL g646 ( .A(n_614), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_615), .B(n_646), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_615), .B(n_637), .Y(n_688) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_618), .A2(n_624), .B1(n_628), .B2(n_630), .Y(n_623) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g639 ( .A(n_620), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g684 ( .A(n_620), .B(n_685), .Y(n_684) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_622), .A2(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_626), .A2(n_635), .B1(n_638), .B2(n_639), .C(n_641), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_626), .B(n_660), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_626), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g742 ( .A(n_632), .Y(n_742) );
INVxp67_ASAP7_75t_L g665 ( .A(n_633), .Y(n_665) );
INVx1_ASAP7_75t_L g672 ( .A(n_635), .Y(n_672) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g711 ( .A(n_636), .B(n_640), .Y(n_711) );
INVx1_ASAP7_75t_L g685 ( .A(n_640), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_640), .B(n_655), .Y(n_715) );
OAI32xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .A3(n_646), .B1(n_647), .B2(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g654 ( .A(n_649), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_649), .B(n_681), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_649), .B(n_710), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g749 ( .A(n_649), .B(n_660), .Y(n_749) );
NAND5xp2_ASAP7_75t_L g650 ( .A(n_651), .B(n_673), .C(n_686), .D(n_698), .E(n_699), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B1(n_656), .B2(n_658), .C(n_662), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp33_ASAP7_75t_SL g677 ( .A(n_657), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_660), .B(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_661), .A2(n_674), .B1(n_677), .B2(n_681), .Y(n_673) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_664), .A2(n_669), .B(n_670), .C(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g696 ( .A(n_676), .Y(n_696) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_685), .B(n_734), .Y(n_744) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_704), .B2(n_708), .C1(n_711), .C2(n_712), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_718), .B2(n_720), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_727), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g734 ( .A(n_726), .Y(n_734) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B1(n_735), .B2(n_737), .C(n_739), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B(n_750), .C(n_752), .Y(n_745) );
INVxp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_755), .Y(n_752) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
endmodule