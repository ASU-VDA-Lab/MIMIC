module fake_jpeg_17852_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_1),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_29),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_3),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_34),
.C(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_49),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_50),
.B(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_39),
.B1(n_38),
.B2(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

BUFx12f_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_59),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_64),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_14),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_51),
.C(n_16),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_15),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_17),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_64),
.B(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_76),
.A2(n_74),
.B1(n_71),
.B2(n_77),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_22),
.B(n_24),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_26),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_28),
.Y(n_83)
);


endmodule