module real_jpeg_29078_n_7 (n_46, n_5, n_4, n_43, n_0, n_1, n_47, n_2, n_45, n_6, n_42, n_44, n_3, n_7);

input n_46;
input n_5;
input n_4;
input n_43;
input n_0;
input n_1;
input n_47;
input n_2;
input n_45;
input n_6;
input n_42;
input n_44;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_0),
.B(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_3),
.B(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_5),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_11),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_15),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_14),
.Y(n_8)
);

CKINVDCx14_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_36),
.B(n_40),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_32),
.B(n_35),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_27),
.B(n_31),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_23),
.B(n_26),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_34),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_42),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_43),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_44),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_45),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_47),
.Y(n_39)
);


endmodule