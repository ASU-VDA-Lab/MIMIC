module fake_netlist_6_2904_n_1553 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1553);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1553;

wire n_992;
wire n_801;
wire n_1458;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_81),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_46),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_7),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_92),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_74),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_38),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_82),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

BUFx8_ASAP7_75t_SL g166 ( 
.A(n_122),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_34),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_91),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_109),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_23),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_1),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_67),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_61),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_103),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_142),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_105),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_59),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_136),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_60),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_52),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_43),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_94),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_141),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_133),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_24),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_8),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_139),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_22),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_15),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_18),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_131),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_58),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_16),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_57),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_134),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_51),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_49),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_106),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_73),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_43),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_56),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_79),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_29),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_1),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_85),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_119),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_117),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_25),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_72),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_127),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_16),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_53),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_26),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_44),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_19),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_108),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_30),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_101),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_146),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_97),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_34),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_100),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_19),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_36),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_27),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_40),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_86),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_54),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_4),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_123),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_36),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_66),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_38),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_30),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_29),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_197),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_197),
.Y(n_297)
);

BUFx2_ASAP7_75t_SL g298 ( 
.A(n_155),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_166),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_255),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_170),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_150),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_170),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_151),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_189),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_189),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_152),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_152),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_154),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_182),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_171),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_212),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_195),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_195),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_199),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_199),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_161),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_161),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_234),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_244),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_158),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_248),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_226),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_252),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_153),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_212),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_234),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_167),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_252),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_208),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_212),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_221),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_163),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_246),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_265),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_265),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_157),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_282),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_162),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_163),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_280),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_177),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_264),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_289),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_165),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_243),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_362),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_157),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_164),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_315),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_297),
.B(n_172),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_298),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_323),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_303),
.B(n_174),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_304),
.B(n_173),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_304),
.B(n_174),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_331),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_305),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_302),
.A2(n_294),
.B1(n_279),
.B2(n_257),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_348),
.A2(n_269),
.B1(n_268),
.B2(n_205),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_296),
.B(n_359),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_299),
.B(n_281),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_332),
.B(n_179),
.Y(n_410)
);

NOR2x1_ASAP7_75t_L g411 ( 
.A(n_333),
.B(n_218),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_354),
.B(n_251),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_251),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_311),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_321),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_313),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_353),
.A2(n_284),
.B1(n_289),
.B2(n_293),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_314),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_336),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_334),
.B(n_243),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_325),
.B(n_176),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_355),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_325),
.A2(n_168),
.B(n_165),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_327),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_365),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_SL g433 ( 
.A(n_418),
.B(n_286),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_382),
.B(n_341),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_382),
.B(n_339),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_343),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_369),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_384),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_428),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_282),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_368),
.B(n_361),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_376),
.B(n_306),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_364),
.C(n_349),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_370),
.B(n_346),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_432),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_370),
.B(n_373),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_386),
.B(n_352),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_392),
.B(n_296),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_R g457 ( 
.A(n_380),
.B(n_178),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_406),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_328),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_425),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_425),
.B(n_180),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_374),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_377),
.B(n_200),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_413),
.B(n_186),
.Y(n_471)
);

OR2x6_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_298),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_406),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_414),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_372),
.A2(n_218),
.B1(n_168),
.B2(n_233),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_413),
.B(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_380),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_377),
.B(n_213),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_388),
.A2(n_214),
.B1(n_224),
.B2(n_291),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_389),
.B(n_372),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_414),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_388),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_374),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_378),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_374),
.Y(n_492)
);

BUFx8_ASAP7_75t_SL g493 ( 
.A(n_395),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_417),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_427),
.B(n_176),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_389),
.B(n_228),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_375),
.A2(n_369),
.B1(n_426),
.B2(n_372),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_426),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_412),
.B(n_169),
.Y(n_505)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_411),
.C(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_379),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_395),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_429),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_398),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_381),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_381),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_416),
.A2(n_181),
.B(n_169),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_374),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_398),
.A2(n_259),
.B1(n_231),
.B2(n_236),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_422),
.B(n_329),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

AO21x2_ASAP7_75t_L g520 ( 
.A1(n_412),
.A2(n_185),
.B(n_183),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_385),
.B(n_187),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_429),
.A2(n_215),
.B1(n_277),
.B2(n_253),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_394),
.B(n_188),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_422),
.B(n_190),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_397),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_424),
.B(n_329),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_396),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_397),
.B(n_399),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

AND3x2_ASAP7_75t_L g534 ( 
.A(n_387),
.B(n_253),
.C(n_183),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_387),
.B(n_216),
.C(n_204),
.Y(n_535)
);

AND3x1_ASAP7_75t_L g536 ( 
.A(n_424),
.B(n_366),
.C(n_363),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_431),
.B(n_191),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_387),
.A2(n_277),
.B1(n_181),
.B2(n_184),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_396),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_396),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_387),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_390),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_400),
.Y(n_544)
);

BUFx6f_ASAP7_75t_SL g545 ( 
.A(n_390),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_390),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_400),
.Y(n_547)
);

OAI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_430),
.A2(n_184),
.B(n_194),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_430),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_431),
.B(n_192),
.Y(n_550)
);

INVx6_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_430),
.B(n_194),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_431),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_401),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_407),
.B(n_193),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_407),
.B(n_209),
.C(n_211),
.Y(n_557)
);

INVx6_ASAP7_75t_L g558 ( 
.A(n_391),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_401),
.A2(n_402),
.B(n_249),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_407),
.B(n_219),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_400),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_401),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_400),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_402),
.A2(n_196),
.B1(n_206),
.B2(n_215),
.Y(n_564)
);

BUFx6f_ASAP7_75t_SL g565 ( 
.A(n_427),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_415),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_391),
.B(n_415),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_391),
.B(n_198),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_427),
.B(n_176),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_453),
.B(n_206),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_439),
.B(n_176),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_450),
.B(n_217),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_483),
.B(n_217),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_487),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_524),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_542),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_439),
.B(n_176),
.Y(n_580)
);

NAND2x1_ASAP7_75t_L g581 ( 
.A(n_551),
.B(n_427),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_460),
.B(n_330),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_462),
.B(n_220),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_230),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_504),
.B(n_330),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_555),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_555),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_477),
.B(n_335),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_469),
.B(n_229),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_496),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_456),
.B(n_201),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_542),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_436),
.A2(n_241),
.B1(n_292),
.B2(n_287),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_232),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_456),
.B(n_202),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_456),
.B(n_203),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_518),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_502),
.B(n_232),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_436),
.B(n_233),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_503),
.B(n_235),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_460),
.B(n_245),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_476),
.B(n_335),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_445),
.B(n_249),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_533),
.A2(n_338),
.B1(n_337),
.B2(n_340),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_419),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_459),
.B(n_419),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_541),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_542),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_506),
.A2(n_225),
.B1(n_275),
.B2(n_274),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_533),
.A2(n_337),
.B1(n_338),
.B2(n_340),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_473),
.B(n_420),
.Y(n_615)
);

OAI221xp5_ASAP7_75t_L g616 ( 
.A1(n_475),
.A2(n_342),
.B1(n_347),
.B2(n_350),
.C(n_351),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_472),
.B(n_342),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_481),
.B(n_420),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_438),
.B(n_238),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_438),
.B(n_239),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_546),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_420),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_509),
.A2(n_391),
.B(n_423),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_488),
.B(n_347),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_443),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_435),
.B(n_250),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_488),
.B(n_350),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_451),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_509),
.B(n_207),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_449),
.B(n_256),
.Y(n_631)
);

AND2x6_ASAP7_75t_SL g632 ( 
.A(n_472),
.B(n_444),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_553),
.B(n_210),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_455),
.B(n_351),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_568),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_437),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_549),
.B(n_421),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_553),
.B(n_222),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_451),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_554),
.B(n_421),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_464),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_472),
.B(n_356),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_505),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_437),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_433),
.B(n_262),
.C(n_258),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_522),
.B(n_223),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_516),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_440),
.B(n_366),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_505),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_464),
.Y(n_652)
);

AO221x1_ASAP7_75t_L g653 ( 
.A1(n_479),
.A2(n_356),
.B1(n_357),
.B2(n_360),
.C(n_363),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_463),
.B(n_427),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_517),
.B(n_290),
.C(n_288),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_433),
.B(n_278),
.C(n_271),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_434),
.B(n_357),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_463),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_440),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_515),
.A2(n_360),
.B(n_263),
.C(n_285),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_458),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_465),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_491),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_498),
.B(n_260),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_R g666 ( 
.A(n_442),
.B(n_227),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_507),
.B(n_247),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_513),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_514),
.B(n_266),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_242),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_528),
.A2(n_283),
.B(n_276),
.C(n_272),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_519),
.B(n_240),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_516),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_471),
.B(n_237),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_474),
.B(n_391),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_148),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_525),
.B(n_145),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_564),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_508),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_474),
.B(n_135),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_545),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g683 ( 
.A(n_516),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_446),
.B(n_5),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_444),
.B(n_10),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_528),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_121),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_526),
.A2(n_112),
.B1(n_102),
.B2(n_93),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_468),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_510),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_470),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_559),
.B(n_83),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_566),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_461),
.B(n_80),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_566),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_461),
.B(n_77),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_461),
.B(n_75),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_480),
.B(n_70),
.Y(n_700)
);

BUFx6f_ASAP7_75t_SL g701 ( 
.A(n_472),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_516),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_482),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

OAI221xp5_ASAP7_75t_L g705 ( 
.A1(n_538),
.A2(n_557),
.B1(n_535),
.B2(n_548),
.C(n_510),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_467),
.B(n_69),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_466),
.B(n_13),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_484),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_467),
.B(n_63),
.Y(n_709)
);

AO22x2_ASAP7_75t_L g710 ( 
.A1(n_441),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_710)
);

INVxp33_ASAP7_75t_L g711 ( 
.A(n_454),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_537),
.B(n_14),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_467),
.B(n_50),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_489),
.B(n_48),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_588),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_574),
.B(n_520),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_624),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_572),
.B(n_583),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_628),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_650),
.B(n_458),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_590),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_686),
.B(n_520),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_672),
.A2(n_550),
.B(n_556),
.C(n_520),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_492),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_619),
.B(n_448),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_704),
.B(n_511),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_578),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_669),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_571),
.B(n_452),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_669),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_620),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_620),
.B(n_452),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_646),
.B(n_492),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_606),
.B(n_552),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_577),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_658),
.B(n_664),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_585),
.B(n_598),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_691),
.B(n_508),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_579),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_668),
.B(n_604),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_694),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_659),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_694),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_679),
.B(n_570),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_617),
.B(n_564),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_607),
.B(n_564),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_659),
.Y(n_747)
);

AO21x1_ASAP7_75t_L g748 ( 
.A1(n_630),
.A2(n_511),
.B(n_494),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_606),
.B(n_540),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_614),
.B(n_529),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_697),
.Y(n_751)
);

BUFx8_ASAP7_75t_SL g752 ( 
.A(n_701),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_608),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_608),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_633),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_614),
.B(n_552),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_529),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_679),
.A2(n_493),
.B1(n_565),
.B2(n_501),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_595),
.B(n_529),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_649),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_707),
.A2(n_493),
.B1(n_565),
.B2(n_570),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_633),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_582),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_661),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_611),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_682),
.B(n_534),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_621),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_584),
.B(n_523),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_666),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_576),
.Y(n_770)
);

NOR2x1p5_ASAP7_75t_L g771 ( 
.A(n_636),
.B(n_569),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_578),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_657),
.Y(n_773)
);

OAI21xp33_ASAP7_75t_SL g774 ( 
.A1(n_625),
.A2(n_600),
.B(n_603),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_696),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_599),
.A2(n_500),
.B1(n_494),
.B2(n_495),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_582),
.B(n_539),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_691),
.B(n_601),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_645),
.B(n_539),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_685),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_584),
.B(n_530),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_578),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_586),
.B(n_587),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_500),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_578),
.B(n_552),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_575),
.B(n_530),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_602),
.B(n_544),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_684),
.A2(n_565),
.B1(n_501),
.B2(n_552),
.Y(n_789)
);

CKINVDCx8_ASAP7_75t_R g790 ( 
.A(n_632),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_612),
.B(n_497),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_612),
.B(n_497),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_692),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_627),
.B(n_495),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_666),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_651),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_707),
.A2(n_499),
.B1(n_512),
.B2(n_523),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_612),
.B(n_499),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_649),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_617),
.B(n_512),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_677),
.B(n_543),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_675),
.B(n_547),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_591),
.A2(n_490),
.B(n_561),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_630),
.A2(n_563),
.B1(n_543),
.B2(n_544),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_563),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_609),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_678),
.B(n_547),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_675),
.B(n_561),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_591),
.A2(n_561),
.B(n_490),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_SL g811 ( 
.A(n_680),
.B(n_567),
.C(n_21),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_701),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_593),
.B(n_670),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_671),
.B(n_532),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_687),
.B(n_532),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_SL g816 ( 
.A(n_690),
.B(n_20),
.C(n_21),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_684),
.A2(n_532),
.B1(n_558),
.B2(n_551),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_711),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_596),
.A2(n_532),
.B(n_558),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_635),
.A2(n_558),
.B1(n_551),
.B2(n_27),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_592),
.Y(n_821)
);

AOI21xp33_ASAP7_75t_L g822 ( 
.A1(n_627),
.A2(n_24),
.B(n_25),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_644),
.B(n_32),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_644),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_665),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_610),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_597),
.A2(n_558),
.B(n_39),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_649),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_635),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_626),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_640),
.A2(n_35),
.B1(n_42),
.B2(n_45),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_673),
.B(n_45),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_615),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_597),
.A2(n_47),
.B(n_623),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_649),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_705),
.B(n_47),
.Y(n_836)
);

CKINVDCx11_ASAP7_75t_R g837 ( 
.A(n_647),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_640),
.A2(n_667),
.B1(n_665),
.B2(n_712),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_629),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_605),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_618),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_631),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_663),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_622),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_641),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_643),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_653),
.A2(n_710),
.B1(n_648),
.B2(n_693),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_631),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_663),
.B(n_674),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_660),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_656),
.B(n_655),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_652),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_639),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_594),
.B(n_672),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_710),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_710),
.A2(n_648),
.B1(n_616),
.B2(n_681),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_681),
.A2(n_700),
.B1(n_689),
.B2(n_662),
.Y(n_857)
);

NOR2x2_ASAP7_75t_L g858 ( 
.A(n_690),
.B(n_708),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_573),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_573),
.A2(n_580),
.B1(n_613),
.B2(n_654),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_688),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_642),
.B(n_683),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_663),
.B(n_702),
.Y(n_863)
);

INVxp33_ASAP7_75t_L g864 ( 
.A(n_580),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_581),
.B(n_700),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_842),
.B(n_663),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_848),
.B(n_703),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_809),
.A2(n_702),
.B(n_674),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_814),
.A2(n_702),
.B(n_674),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_717),
.B(n_660),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_721),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_779),
.B(n_676),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_779),
.A2(n_699),
.B(n_713),
.C(n_709),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_764),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_741),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_769),
.B(n_695),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_R g877 ( 
.A(n_747),
.B(n_698),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_819),
.A2(n_706),
.B(n_714),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_744),
.A2(n_634),
.B1(n_758),
.B2(n_861),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_728),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_837),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_741),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_843),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_SL g884 ( 
.A1(n_744),
.A2(n_634),
.B(n_758),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_725),
.B(n_634),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_SL g886 ( 
.A(n_824),
.B(n_738),
.C(n_729),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_720),
.B(n_715),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_719),
.B(n_818),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_763),
.B(n_740),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_742),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_763),
.B(n_825),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_727),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_742),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_836),
.A2(n_822),
.B(n_832),
.C(n_854),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_732),
.B(n_773),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_803),
.A2(n_810),
.B(n_804),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_729),
.B(n_795),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_718),
.B(n_853),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_788),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_807),
.B(n_826),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_727),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_836),
.A2(n_854),
.B1(n_850),
.B2(n_785),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_813),
.A2(n_862),
.B(n_787),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_840),
.A2(n_736),
.B(n_853),
.C(n_774),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_840),
.B(n_833),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_841),
.B(n_844),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_834),
.A2(n_855),
.B(n_765),
.C(n_767),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_838),
.A2(n_851),
.B1(n_781),
.B2(n_771),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_752),
.Y(n_909)
);

CKINVDCx11_ASAP7_75t_R g910 ( 
.A(n_790),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_766),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_768),
.B(n_775),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_727),
.B(n_772),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_743),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_738),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_784),
.B(n_806),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_727),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_856),
.A2(n_847),
.B1(n_746),
.B2(n_778),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_864),
.B(n_797),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_778),
.A2(n_794),
.B1(n_761),
.B2(n_797),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_772),
.B(n_783),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_801),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_772),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_751),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_864),
.B(n_770),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_858),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_823),
.B(n_859),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_723),
.A2(n_856),
.B(n_847),
.C(n_860),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_816),
.A2(n_811),
.B(n_716),
.C(n_722),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_R g930 ( 
.A(n_812),
.B(n_783),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_783),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_766),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_761),
.A2(n_829),
.B1(n_831),
.B2(n_750),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_749),
.A2(n_745),
.B1(n_820),
.B2(n_816),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_823),
.B(n_811),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_730),
.B(n_780),
.Y(n_936)
);

BUFx8_ASAP7_75t_SL g937 ( 
.A(n_801),
.Y(n_937)
);

AOI221x1_ASAP7_75t_L g938 ( 
.A1(n_827),
.A2(n_782),
.B1(n_805),
.B2(n_759),
.C(n_757),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_801),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_815),
.A2(n_756),
.B(n_734),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_SL g941 ( 
.A(n_800),
.B(n_730),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_791),
.A2(n_799),
.B(n_792),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_735),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_745),
.A2(n_789),
.B1(n_760),
.B2(n_756),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_835),
.B(n_865),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_815),
.A2(n_734),
.B(n_808),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_846),
.B(n_739),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_SL g948 ( 
.A(n_800),
.B(n_760),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_835),
.Y(n_949)
);

AOI22x1_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_762),
.B1(n_755),
.B2(n_793),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_828),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_726),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_776),
.A2(n_857),
.B(n_755),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_SL g954 ( 
.A(n_798),
.B(n_724),
.C(n_733),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_739),
.B(n_753),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_865),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_726),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_808),
.A2(n_802),
.B(n_799),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_726),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_776),
.A2(n_796),
.B(n_777),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_802),
.A2(n_792),
.B(n_791),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_849),
.B(n_863),
.C(n_786),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_726),
.A2(n_865),
.B1(n_845),
.B2(n_839),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_726),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_821),
.B(n_839),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_830),
.B(n_845),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_830),
.B(n_852),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_852),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_849),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_817),
.B(n_742),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_731),
.A2(n_779),
.B(n_450),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_842),
.B(n_848),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_731),
.B(n_737),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_731),
.B(n_842),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_720),
.B(n_588),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_842),
.B(n_848),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_943),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_975),
.B(n_926),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_958),
.A2(n_869),
.B(n_868),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_915),
.A2(n_897),
.B1(n_926),
.B2(n_974),
.Y(n_981)
);

CKINVDCx11_ASAP7_75t_R g982 ( 
.A(n_910),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_928),
.A2(n_902),
.B(n_903),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_898),
.B(n_973),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_953),
.A2(n_885),
.B(n_907),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_933),
.A2(n_953),
.B(n_866),
.C(n_946),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_887),
.B(n_895),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_959),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_940),
.A2(n_942),
.B(n_878),
.Y(n_989)
);

AO21x1_ASAP7_75t_L g990 ( 
.A1(n_933),
.A2(n_904),
.B(n_944),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_935),
.B(n_899),
.Y(n_991)
);

CKINVDCx11_ASAP7_75t_R g992 ( 
.A(n_874),
.Y(n_992)
);

NOR4xp25_ASAP7_75t_L g993 ( 
.A(n_929),
.B(n_934),
.C(n_879),
.D(n_918),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_970),
.B(n_945),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_SL g995 ( 
.A1(n_970),
.A2(n_879),
.B(n_944),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_956),
.A2(n_872),
.B1(n_927),
.B2(n_919),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_972),
.A2(n_976),
.B(n_870),
.C(n_900),
.Y(n_997)
);

AOI221x1_ASAP7_75t_L g998 ( 
.A1(n_934),
.A2(n_954),
.B1(n_960),
.B2(n_941),
.C(n_925),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_900),
.B(n_906),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_871),
.B(n_905),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_875),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_888),
.Y(n_1002)
);

AO31x2_ASAP7_75t_L g1003 ( 
.A1(n_969),
.A2(n_966),
.A3(n_967),
.B(n_947),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_889),
.A2(n_891),
.B(n_912),
.C(n_884),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_890),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_901),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_916),
.B(n_867),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_920),
.A2(n_963),
.B(n_962),
.C(n_886),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_892),
.A2(n_923),
.B(n_931),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_892),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_882),
.A2(n_924),
.B(n_914),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_913),
.A2(n_921),
.B(n_959),
.C(n_936),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_892),
.A2(n_923),
.B(n_931),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_880),
.A2(n_957),
.B(n_952),
.C(n_965),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_952),
.A2(n_965),
.B(n_964),
.C(n_968),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_911),
.B(n_893),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_SL g1017 ( 
.A(n_876),
.B(n_877),
.C(n_881),
.Y(n_1017)
);

AO21x2_ASAP7_75t_L g1018 ( 
.A1(n_955),
.A2(n_930),
.B(n_945),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_932),
.B(n_909),
.C(n_949),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_917),
.A2(n_937),
.B(n_968),
.C(n_883),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_931),
.A2(n_968),
.B(n_951),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_951),
.A2(n_931),
.A3(n_901),
.B(n_883),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_975),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_928),
.A2(n_748),
.A3(n_938),
.B(n_873),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.C(n_854),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_939),
.B(n_922),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_892),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_939),
.B(n_922),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_943),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_959),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_888),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_898),
.B(n_731),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_898),
.B(n_731),
.Y(n_1035)
);

AO32x2_ASAP7_75t_L g1036 ( 
.A1(n_933),
.A2(n_855),
.A3(n_934),
.B1(n_944),
.B2(n_879),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_898),
.B(n_731),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.C(n_854),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_874),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1041)
);

AOI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_898),
.B(n_731),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.C(n_854),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_971),
.A2(n_779),
.B1(n_731),
.B2(n_836),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_971),
.B(n_779),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_971),
.A2(n_779),
.B(n_731),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_895),
.B(n_725),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_910),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_L g1053 ( 
.A(n_971),
.B(n_861),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_874),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_928),
.A2(n_748),
.A3(n_938),
.B(n_873),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_971),
.B(n_779),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_898),
.B(n_731),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_890),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_894),
.A2(n_971),
.B(n_731),
.C(n_854),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_943),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_892),
.B(n_923),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_943),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_902),
.A2(n_744),
.B1(n_758),
.B2(n_928),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_943),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_971),
.B(n_731),
.C(n_732),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_SL g1068 ( 
.A1(n_928),
.A2(n_612),
.B(n_578),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_939),
.B(n_922),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_948),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_971),
.A2(n_779),
.B(n_731),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_898),
.B(n_731),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_898),
.B(n_731),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_939),
.B(n_922),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_898),
.B(n_731),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_928),
.A2(n_731),
.B(n_574),
.C(n_834),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_900),
.B(n_902),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_910),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_874),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_SL g1082 ( 
.A1(n_928),
.A2(n_612),
.B(n_578),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_928),
.A2(n_748),
.A3(n_938),
.B(n_873),
.Y(n_1083)
);

OAI22x1_ASAP7_75t_L g1084 ( 
.A1(n_908),
.A2(n_779),
.B1(n_855),
.B2(n_836),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_898),
.B(n_731),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_950),
.A2(n_961),
.B(n_896),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_928),
.A2(n_748),
.A3(n_938),
.B(n_873),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_943),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_928),
.A2(n_894),
.B(n_902),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_994),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1064),
.A2(n_1056),
.B1(n_1046),
.B2(n_1045),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_1033),
.B(n_1054),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_978),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_982),
.Y(n_1095)
);

AO21x1_ASAP7_75t_L g1096 ( 
.A1(n_1064),
.A2(n_1041),
.B(n_1037),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1026),
.A2(n_1044),
.B(n_1039),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_994),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1090),
.A2(n_1071),
.B(n_1037),
.C(n_1041),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1062),
.A2(n_1090),
.B1(n_1071),
.B2(n_1066),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1029),
.A2(n_1072),
.B(n_1086),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1047),
.A2(n_1050),
.B(n_980),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1084),
.A2(n_1007),
.B1(n_1002),
.B2(n_991),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_992),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1067),
.B(n_1059),
.C(n_1053),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_987),
.B(n_979),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1079),
.B(n_999),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1049),
.B(n_1073),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_994),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_1040),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_981),
.A2(n_1074),
.B1(n_1057),
.B2(n_1038),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_988),
.B(n_1032),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1010),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1023),
.B(n_1016),
.Y(n_1115)
);

AOI22x1_ASAP7_75t_L g1116 ( 
.A1(n_1062),
.A2(n_1066),
.B1(n_1070),
.B2(n_983),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_1052),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1080),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_990),
.A2(n_1008),
.A3(n_1014),
.B(n_1015),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1079),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_984),
.B(n_996),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_995),
.B(n_1020),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_1081),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1005),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1016),
.B(n_1076),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1034),
.A2(n_1075),
.B1(n_1035),
.B2(n_1085),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1004),
.B(n_997),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1078),
.A2(n_986),
.B(n_1042),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_1048),
.A2(n_1012),
.B(n_1049),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1031),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1051),
.B(n_1000),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1073),
.A2(n_1089),
.B(n_1060),
.C(n_1088),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1058),
.B(n_1017),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1061),
.B(n_1021),
.Y(n_1135)
);

BUFx2_ASAP7_75t_R g1136 ( 
.A(n_1018),
.Y(n_1136)
);

INVx5_ASAP7_75t_L g1137 ( 
.A(n_1028),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1024),
.A2(n_1087),
.A3(n_1083),
.B(n_1055),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1063),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1065),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1027),
.B(n_1076),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1011),
.A2(n_1009),
.B(n_1013),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_993),
.A2(n_1018),
.B(n_1083),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1030),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1069),
.A2(n_1019),
.B1(n_993),
.B2(n_1036),
.Y(n_1145)
);

CKINVDCx11_ASAP7_75t_R g1146 ( 
.A(n_1006),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1036),
.A2(n_1003),
.B(n_1022),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1022),
.B(n_1006),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1022),
.A2(n_971),
.B1(n_1064),
.B2(n_731),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1040),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1049),
.B(n_971),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1068),
.B(n_1082),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_978),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1005),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_978),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1064),
.A2(n_971),
.B1(n_731),
.B2(n_1046),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1078),
.A2(n_894),
.B(n_1026),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_990),
.A2(n_928),
.A3(n_998),
.B(n_985),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1064),
.A2(n_971),
.B1(n_731),
.B2(n_1046),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1053),
.A2(n_731),
.B1(n_324),
.B2(n_353),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1001),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1079),
.B(n_999),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1010),
.B(n_892),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_978),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1064),
.A2(n_971),
.B1(n_731),
.B2(n_1046),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1006),
.Y(n_1168)
);

AOI222xp33_ASAP7_75t_L g1169 ( 
.A1(n_1064),
.A2(n_680),
.B1(n_779),
.B2(n_971),
.C1(n_1041),
.C2(n_1037),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_992),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1006),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1064),
.A2(n_971),
.B1(n_731),
.B2(n_1046),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1175)
);

AOI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1046),
.A2(n_894),
.B(n_731),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1006),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1078),
.A2(n_894),
.B(n_1026),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_989),
.A2(n_1025),
.B(n_977),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1121),
.B(n_1107),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1094),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1132),
.B(n_1115),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1101),
.A2(n_1160),
.B1(n_1092),
.B2(n_1100),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1101),
.A2(n_1092),
.B1(n_1100),
.B2(n_1156),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1091),
.B(n_1099),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1113),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1174),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1129),
.B(n_1126),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1125),
.B(n_1144),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1091),
.B(n_1099),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1156),
.A2(n_1166),
.B1(n_1159),
.B2(n_1173),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1159),
.A2(n_1166),
.B1(n_1173),
.B2(n_1106),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1126),
.B(n_1112),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1145),
.A2(n_1152),
.B1(n_1136),
.B2(n_1093),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1123),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1112),
.B(n_1108),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1125),
.B(n_1141),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1110),
.B(n_1122),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1120),
.B(n_1110),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1111),
.B(n_1162),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1096),
.A2(n_1157),
.B(n_1178),
.C(n_1098),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1169),
.A2(n_1176),
.B(n_1098),
.C(n_1178),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1104),
.B(n_1145),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1151),
.B(n_1169),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1127),
.A2(n_1122),
.B(n_1133),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1128),
.A2(n_1143),
.B(n_1157),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1127),
.B(n_1150),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1122),
.B(n_1148),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1147),
.Y(n_1209)
);

BUFx2_ASAP7_75t_SL g1210 ( 
.A(n_1095),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1147),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1128),
.A2(n_1143),
.B(n_1102),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1149),
.A2(n_1134),
.B1(n_1116),
.B2(n_1139),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1134),
.A2(n_1139),
.B1(n_1109),
.B2(n_1154),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1103),
.A2(n_1179),
.B(n_1175),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1146),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_1124),
.B(n_1161),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1131),
.B(n_1140),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1170),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1153),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1155),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1105),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1118),
.B(n_1171),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1164),
.B(n_1158),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1138),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1172),
.B(n_1119),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1138),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1114),
.B(n_1137),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1135),
.B(n_1119),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1172),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1130),
.B(n_1146),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1172),
.B(n_1177),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1117),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_SL g1234 ( 
.A(n_1168),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_L g1235 ( 
.A1(n_1114),
.A2(n_1142),
.B(n_1113),
.C(n_1165),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1113),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1177),
.B(n_1113),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1163),
.A2(n_1128),
.B(n_1143),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1100),
.A2(n_1101),
.B(n_971),
.C(n_928),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1101),
.A2(n_981),
.B1(n_779),
.B2(n_1045),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1121),
.B(n_1107),
.Y(n_1241)
);

AND2x6_ASAP7_75t_L g1242 ( 
.A(n_1109),
.B(n_963),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1101),
.A2(n_981),
.B1(n_779),
.B2(n_1045),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_981),
.B1(n_779),
.B2(n_1045),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1128),
.A2(n_1143),
.B(n_1157),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1121),
.B(n_1107),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1198),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1206),
.B(n_1245),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1238),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1206),
.B(n_1245),
.Y(n_1250)
);

OR2x2_ASAP7_75t_SL g1251 ( 
.A(n_1193),
.B(n_1204),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1188),
.B(n_1183),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1238),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_SL g1254 ( 
.A(n_1186),
.B(n_1202),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1227),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1186),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1184),
.A2(n_1244),
.B1(n_1243),
.B2(n_1240),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1238),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1225),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_1224),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1206),
.B(n_1245),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1211),
.B(n_1212),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1211),
.B(n_1212),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1199),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1239),
.A2(n_1205),
.B(n_1196),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1181),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1201),
.A2(n_1235),
.B(n_1239),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1219),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1219),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1198),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1220),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1215),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1229),
.B(n_1226),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1221),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1229),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1205),
.A2(n_1213),
.B(n_1192),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1214),
.B(n_1203),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1218),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1186),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1191),
.A2(n_1231),
.B(n_1194),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1231),
.A2(n_1208),
.B(n_1185),
.Y(n_1282)
);

OR2x6_ASAP7_75t_L g1283 ( 
.A(n_1190),
.B(n_1236),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1236),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1270),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1263),
.B(n_1200),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1248),
.B(n_1180),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1248),
.B(n_1246),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1248),
.B(n_1241),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1250),
.B(n_1242),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1263),
.B(n_1187),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1260),
.B(n_1242),
.Y(n_1292)
);

AND2x2_ASAP7_75t_SL g1293 ( 
.A(n_1257),
.B(n_1216),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1261),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1270),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1260),
.B(n_1242),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1276),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1265),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1280),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1265),
.B(n_1187),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1262),
.B(n_1207),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1252),
.B(n_1207),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1262),
.B(n_1182),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1264),
.B(n_1232),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_SL g1305 ( 
.A(n_1256),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1273),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1264),
.B(n_1230),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1269),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1257),
.A2(n_1189),
.B1(n_1216),
.B2(n_1197),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1255),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1261),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1293),
.B(n_1252),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1294),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1307),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1302),
.A2(n_1254),
.B1(n_1278),
.B2(n_1283),
.Y(n_1315)
);

OAI211xp5_ASAP7_75t_L g1316 ( 
.A1(n_1302),
.A2(n_1278),
.B(n_1268),
.C(n_1284),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1285),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1293),
.B(n_1254),
.C(n_1268),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_R g1319 ( 
.A(n_1300),
.B(n_1233),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1293),
.A2(n_1277),
.B1(n_1281),
.B2(n_1266),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1301),
.B(n_1282),
.Y(n_1321)
);

NOR4xp25_ASAP7_75t_SL g1322 ( 
.A(n_1293),
.B(n_1258),
.C(n_1253),
.D(n_1249),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1301),
.B(n_1287),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1299),
.B(n_1283),
.Y(n_1324)
);

AOI33xp33_ASAP7_75t_L g1325 ( 
.A1(n_1309),
.A2(n_1284),
.A3(n_1279),
.B1(n_1267),
.B2(n_1272),
.B3(n_1275),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1309),
.A2(n_1251),
.B1(n_1268),
.B2(n_1216),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1294),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1301),
.B(n_1282),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1311),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1299),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1298),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1311),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1298),
.Y(n_1333)
);

AOI31xp33_ASAP7_75t_L g1334 ( 
.A1(n_1292),
.A2(n_1251),
.A3(n_1233),
.B(n_1271),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1287),
.B(n_1282),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_R g1336 ( 
.A(n_1305),
.B(n_1222),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1297),
.B(n_1282),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1303),
.B(n_1286),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1295),
.A2(n_1258),
.B(n_1249),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1292),
.A2(n_1277),
.B1(n_1281),
.B2(n_1266),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1304),
.B(n_1286),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1310),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1296),
.A2(n_1251),
.B1(n_1217),
.B2(n_1271),
.Y(n_1343)
);

AOI22x1_ASAP7_75t_L g1344 ( 
.A1(n_1290),
.A2(n_1216),
.B1(n_1210),
.B2(n_1195),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1296),
.A2(n_1283),
.B1(n_1280),
.B2(n_1256),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1300),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1287),
.B(n_1282),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1305),
.A2(n_1271),
.B1(n_1247),
.B2(n_1283),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1288),
.B(n_1274),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1310),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1339),
.B(n_1317),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1339),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1342),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1324),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1341),
.B(n_1291),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1324),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1339),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1342),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1335),
.B(n_1249),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1318),
.A2(n_1277),
.B(n_1266),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1324),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1350),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_SL g1363 ( 
.A(n_1322),
.B(n_1223),
.C(n_1291),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1339),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1350),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1335),
.B(n_1308),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1313),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1327),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1327),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1330),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1320),
.A2(n_1306),
.B(n_1295),
.Y(n_1372)
);

BUFx8_ASAP7_75t_L g1373 ( 
.A(n_1316),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1329),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1329),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1332),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1346),
.B(n_1288),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1354),
.B(n_1361),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1353),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1351),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1351),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1371),
.B(n_1347),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1353),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1371),
.B(n_1321),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1353),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1371),
.B(n_1321),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1358),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1351),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1358),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1358),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1362),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1368),
.B(n_1332),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1371),
.B(n_1328),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1368),
.B(n_1331),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1362),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1362),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1367),
.B(n_1333),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1360),
.B(n_1336),
.Y(n_1399)
);

OAI33xp33_ASAP7_75t_L g1400 ( 
.A1(n_1367),
.A2(n_1312),
.A3(n_1326),
.B1(n_1315),
.B2(n_1343),
.B3(n_1259),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1351),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1354),
.B(n_1337),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1367),
.B(n_1314),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1337),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1361),
.B(n_1324),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1363),
.A2(n_1326),
.B(n_1340),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1365),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1356),
.B(n_1330),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1365),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1360),
.A2(n_1277),
.B(n_1322),
.Y(n_1410)
);

AOI33xp33_ASAP7_75t_L g1411 ( 
.A1(n_1369),
.A2(n_1345),
.A3(n_1314),
.B1(n_1337),
.B2(n_1279),
.B3(n_1288),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1356),
.B(n_1330),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1356),
.B(n_1323),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_R g1414 ( 
.A(n_1356),
.B(n_1319),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1356),
.B(n_1323),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1356),
.B(n_1349),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1355),
.B(n_1341),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1369),
.B(n_1289),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1355),
.B(n_1338),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1394),
.B(n_1355),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1411),
.B(n_1378),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1419),
.B(n_1377),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1399),
.B(n_1363),
.C(n_1334),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1380),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1378),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1378),
.B(n_1359),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1419),
.B(n_1377),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1400),
.A2(n_1406),
.B1(n_1277),
.B2(n_1373),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1379),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1396),
.B(n_1349),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1408),
.B(n_1359),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1396),
.B(n_1325),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1394),
.B(n_1369),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1414),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1405),
.B(n_1370),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_L g1436 ( 
.A(n_1406),
.B(n_1344),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1380),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1380),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1417),
.B(n_1370),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1384),
.B(n_1289),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1408),
.B(n_1359),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1379),
.Y(n_1442)
);

OAI32xp33_ASAP7_75t_L g1443 ( 
.A1(n_1400),
.A2(n_1352),
.A3(n_1364),
.B1(n_1357),
.B2(n_1373),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1412),
.B(n_1359),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1381),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1383),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1383),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1410),
.A2(n_1334),
.B1(n_1344),
.B2(n_1299),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1366),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1405),
.B(n_1410),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1417),
.B(n_1286),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1384),
.B(n_1289),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1398),
.B(n_1370),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1386),
.B(n_1303),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1425),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1423),
.A2(n_1373),
.B1(n_1405),
.B2(n_1281),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1386),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1429),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1420),
.B(n_1398),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1436),
.A2(n_1373),
.B1(n_1281),
.B2(n_1405),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1435),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1436),
.A2(n_1414),
.B(n_1372),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1442),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1421),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1428),
.A2(n_1373),
.B1(n_1281),
.B2(n_1266),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1393),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1450),
.B(n_1393),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1446),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1426),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1426),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1420),
.B(n_1392),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1432),
.B(n_1413),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1431),
.B(n_1413),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1448),
.B(n_1373),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.B(n_1382),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1447),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_1415),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1457),
.B(n_1441),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1465),
.A2(n_1450),
.B1(n_1430),
.B2(n_1422),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1457),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1464),
.A2(n_1443),
.B1(n_1433),
.B2(n_1453),
.C(n_1444),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1456),
.A2(n_1444),
.B(n_1382),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1477),
.B(n_1449),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1415),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1455),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

XNOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1462),
.B(n_1348),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1477),
.B(n_1416),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

AOI221x1_ASAP7_75t_SL g1493 ( 
.A1(n_1468),
.A2(n_1478),
.B1(n_1463),
.B2(n_1474),
.C(n_1470),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1460),
.A2(n_1454),
.B1(n_1440),
.B2(n_1452),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1467),
.A2(n_1439),
.B(n_1404),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1476),
.A2(n_1403),
.B(n_1433),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1466),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1467),
.A2(n_1451),
.B1(n_1416),
.B2(n_1439),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1483),
.A2(n_1469),
.B1(n_1470),
.B2(n_1471),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1469),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1480),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1486),
.B(n_1459),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1481),
.A2(n_1471),
.B1(n_1467),
.B2(n_1479),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1459),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1497),
.B(n_1461),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1485),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1487),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1493),
.B(n_1461),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1496),
.B(n_1473),
.Y(n_1510)
);

OAI21xp33_ASAP7_75t_L g1511 ( 
.A1(n_1503),
.A2(n_1490),
.B(n_1484),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1510),
.B(n_1495),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1509),
.A2(n_1493),
.B1(n_1498),
.B2(n_1489),
.C(n_1492),
.Y(n_1513)
);

AOI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1501),
.A2(n_1494),
.B(n_1478),
.C(n_1463),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1499),
.A2(n_1467),
.B1(n_1475),
.B2(n_1473),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1504),
.B(n_1453),
.Y(n_1516)
);

OAI211xp5_ASAP7_75t_L g1517 ( 
.A1(n_1505),
.A2(n_1445),
.B(n_1438),
.C(n_1437),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1507),
.A2(n_1445),
.B(n_1438),
.C(n_1437),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1506),
.A2(n_1404),
.B(n_1402),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1516),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1511),
.A2(n_1508),
.B1(n_1500),
.B2(n_1502),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1518),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1512),
.A2(n_1515),
.B1(n_1513),
.B2(n_1519),
.Y(n_1523)
);

OAI222xp33_ASAP7_75t_L g1524 ( 
.A1(n_1514),
.A2(n_1424),
.B1(n_1381),
.B2(n_1388),
.C1(n_1401),
.C2(n_1404),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1520),
.B(n_1424),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1523),
.B(n_1403),
.C(n_1392),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1521),
.B(n_1402),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1522),
.B(n_1418),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1524),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1528),
.A2(n_1402),
.B1(n_1409),
.B2(n_1407),
.Y(n_1531)
);

NOR2xp67_ASAP7_75t_L g1532 ( 
.A(n_1530),
.B(n_1381),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1525),
.A2(n_1388),
.B1(n_1401),
.B2(n_1364),
.C(n_1357),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1529),
.A2(n_1385),
.B1(n_1409),
.B2(n_1407),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1526),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1527),
.B(n_1401),
.C(n_1388),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1532),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1531),
.B(n_1385),
.Y(n_1538)
);

AND3x4_ASAP7_75t_L g1539 ( 
.A(n_1537),
.B(n_1533),
.C(n_1534),
.Y(n_1539)
);

AOI322xp5_ASAP7_75t_L g1540 ( 
.A1(n_1539),
.A2(n_1538),
.A3(n_1536),
.B1(n_1352),
.B2(n_1357),
.C1(n_1364),
.C2(n_1395),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_SL g1541 ( 
.A(n_1540),
.B(n_1357),
.C(n_1352),
.Y(n_1541)
);

CKINVDCx14_ASAP7_75t_R g1542 ( 
.A(n_1541),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1542),
.Y(n_1543)
);

AOI22x1_ASAP7_75t_L g1544 ( 
.A1(n_1543),
.A2(n_1390),
.B1(n_1387),
.B2(n_1397),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1543),
.A2(n_1387),
.B1(n_1397),
.B2(n_1395),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1545),
.A2(n_1389),
.B1(n_1390),
.B2(n_1391),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1544),
.A2(n_1389),
.B1(n_1391),
.B2(n_1352),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1547),
.B(n_1228),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1546),
.B(n_1374),
.Y(n_1549)
);

XNOR2xp5_ASAP7_75t_L g1550 ( 
.A(n_1549),
.B(n_1234),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1548),
.A2(n_1364),
.B1(n_1375),
.B2(n_1376),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1550),
.A2(n_1375),
.B1(n_1374),
.B2(n_1376),
.Y(n_1552)
);

AOI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1552),
.A2(n_1551),
.B(n_1237),
.C(n_1375),
.Y(n_1553)
);


endmodule