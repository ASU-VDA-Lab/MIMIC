module fake_jpeg_11394_n_613 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_554;
wire n_280;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_64),
.Y(n_123)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_70),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_15),
.C(n_14),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_46),
.C(n_29),
.Y(n_157)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_12),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_82),
.B(n_85),
.Y(n_160)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_15),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_100),
.Y(n_161)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_10),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_30),
.B(n_10),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_108),
.Y(n_167)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_35),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_112),
.Y(n_181)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_30),
.B(n_11),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_17),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_19),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_46),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_128),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_132),
.B(n_159),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_64),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_139),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_77),
.A2(n_42),
.B1(n_28),
.B2(n_38),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_190),
.B(n_198),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_23),
.B1(n_38),
.B2(n_27),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_145),
.A2(n_182),
.B1(n_200),
.B2(n_36),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_57),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_148),
.B(n_171),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_11),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_75),
.A2(n_47),
.B(n_29),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_66),
.B(n_41),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_62),
.A2(n_38),
.B1(n_23),
.B2(n_43),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_67),
.B(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_43),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_75),
.A2(n_38),
.B1(n_23),
.B2(n_35),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_70),
.B(n_49),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_76),
.A2(n_117),
.B1(n_116),
.B2(n_114),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_182),
.B1(n_172),
.B2(n_152),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_110),
.A2(n_33),
.B1(n_56),
.B2(n_55),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_79),
.B(n_33),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_84),
.A2(n_27),
.B1(n_49),
.B2(n_47),
.Y(n_200)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_203),
.Y(n_309)
);

AO22x2_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_109),
.B1(n_105),
.B2(n_104),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_204),
.B(n_274),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_213),
.Y(n_275)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

NAND2x1_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_103),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_209),
.A2(n_273),
.B(n_3),
.Y(n_310)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_123),
.A2(n_95),
.B1(n_89),
.B2(n_88),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_211),
.A2(n_212),
.B1(n_259),
.B2(n_260),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_87),
.B1(n_57),
.B2(n_56),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_55),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_214),
.B(n_215),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_53),
.Y(n_215)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_217),
.B(n_262),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_145),
.A2(n_53),
.B1(n_48),
.B2(n_19),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_221),
.A2(n_241),
.B1(n_263),
.B2(n_137),
.Y(n_289)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_223),
.B(n_228),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_48),
.B1(n_39),
.B2(n_37),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_225),
.A2(n_226),
.B1(n_246),
.B2(n_265),
.Y(n_288)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_39),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_126),
.Y(n_229)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_230),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_11),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_232),
.Y(n_292)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_0),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_235),
.Y(n_299)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_236),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_237),
.Y(n_305)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_243),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_131),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_40),
.B1(n_36),
.B2(n_26),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_245),
.B(n_249),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_190),
.A2(n_40),
.B1(n_36),
.B2(n_26),
.Y(n_246)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_149),
.Y(n_248)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_167),
.B(n_1),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_251),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_163),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_167),
.B(n_1),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_254),
.Y(n_316)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_125),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_256),
.Y(n_320)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_258),
.Y(n_324)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_127),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_181),
.A2(n_40),
.A3(n_36),
.B1(n_26),
.B2(n_6),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_26),
.B(n_3),
.C(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_130),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_200),
.A2(n_195),
.B1(n_147),
.B2(n_175),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_264),
.B(n_268),
.Y(n_325)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_272),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_155),
.A2(n_36),
.B1(n_26),
.B2(n_5),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_181),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_133),
.B(n_2),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_206),
.B(n_198),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_276),
.B(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_180),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_201),
.C(n_158),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_278),
.B(n_247),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_226),
.A2(n_183),
.B1(n_189),
.B2(n_177),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_279),
.A2(n_307),
.B1(n_321),
.B2(n_211),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_244),
.A2(n_137),
.B(n_143),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_285),
.A2(n_284),
.B(n_294),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_209),
.B(n_153),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_302),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_289),
.B(n_308),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_177),
.B1(n_140),
.B2(n_170),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_293),
.A2(n_295),
.B1(n_248),
.B2(n_260),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_241),
.A2(n_140),
.B1(n_170),
.B2(n_142),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_240),
.A2(n_174),
.B1(n_176),
.B2(n_142),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_176),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_221),
.B(n_2),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_303),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_220),
.B(n_2),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_306),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_226),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_2),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_310),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_224),
.B(n_6),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_328),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_230),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_319),
.A2(n_322),
.B1(n_205),
.B2(n_271),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_204),
.A2(n_8),
.B1(n_9),
.B2(n_263),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_238),
.A2(n_8),
.B1(n_210),
.B2(n_253),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_218),
.B(n_242),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_204),
.B(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_267),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_216),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_205),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_345),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_275),
.B(n_204),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_369),
.Y(n_380)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_357),
.B1(n_308),
.B2(n_295),
.Y(n_388)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_340),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_342),
.B(n_367),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_285),
.A2(n_272),
.B(n_212),
.C(n_247),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g406 ( 
.A1(n_343),
.A2(n_281),
.B1(n_317),
.B2(n_331),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_314),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_275),
.B(n_203),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_346),
.B(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_329),
.A2(n_266),
.B1(n_270),
.B2(n_229),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_349),
.A2(n_372),
.B1(n_288),
.B2(n_302),
.Y(n_400)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_351),
.Y(n_381)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_314),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_360),
.Y(n_412)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_356),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_287),
.A2(n_288),
.B1(n_307),
.B2(n_276),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_286),
.A2(n_264),
.B1(n_256),
.B2(n_227),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_281),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_324),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_278),
.C(n_323),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_277),
.B(n_219),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_311),
.B(n_239),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_365),
.B(n_366),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_259),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_290),
.B(n_236),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_370),
.B(n_374),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_324),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_373),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_289),
.A2(n_236),
.B1(n_287),
.B2(n_308),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_304),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_290),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_333),
.B(n_313),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_377),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_369),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_392),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_373),
.B(n_316),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_386),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_316),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_332),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_388),
.A2(n_410),
.B1(n_350),
.B2(n_346),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_353),
.B(n_371),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_405),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_349),
.Y(n_392)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_402),
.B1(n_355),
.B2(n_364),
.Y(n_426)
);

OAI22x1_ASAP7_75t_SL g402 ( 
.A1(n_372),
.A2(n_303),
.B1(n_306),
.B2(n_308),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_299),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_407),
.B(n_334),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_357),
.A2(n_293),
.B1(n_323),
.B2(n_303),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_299),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_339),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_428),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_359),
.B(n_332),
.Y(n_415)
);

AO21x1_ASAP7_75t_L g478 ( 
.A1(n_415),
.A2(n_426),
.B(n_330),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_388),
.A2(n_335),
.B1(n_342),
.B2(n_367),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_416),
.A2(n_432),
.B1(n_434),
.B2(n_384),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_418),
.A2(n_444),
.B(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_341),
.Y(n_420)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_361),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_422),
.C(n_437),
.Y(n_449)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_423),
.Y(n_477)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_338),
.B1(n_355),
.B2(n_364),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_427),
.A2(n_430),
.B1(n_433),
.B2(n_435),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_396),
.B(n_341),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_355),
.B1(n_350),
.B2(n_354),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_385),
.B(n_363),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_410),
.A2(n_334),
.B1(n_343),
.B2(n_363),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_409),
.A2(n_382),
.B1(n_402),
.B2(n_380),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_440),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_323),
.C(n_343),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_343),
.B1(n_359),
.B2(n_370),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_438),
.A2(n_407),
.B1(n_406),
.B2(n_408),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_327),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_439),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_389),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_292),
.Y(n_441)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_318),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_442),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_343),
.C(n_331),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_445),
.C(n_391),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_408),
.A2(n_351),
.B1(n_336),
.B2(n_315),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_292),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_394),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_379),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_448),
.A2(n_444),
.B(n_426),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_450),
.A2(n_458),
.B1(n_447),
.B2(n_413),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_412),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_460),
.Y(n_483)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_455),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_416),
.A2(n_392),
.B1(n_391),
.B2(n_406),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_418),
.A2(n_412),
.B(n_406),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_467),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_405),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_466),
.C(n_468),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_386),
.C(n_377),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_415),
.Y(n_485)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_401),
.C(n_398),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_305),
.C(n_381),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_383),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_476),
.C(n_325),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_381),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_472),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_434),
.A2(n_383),
.B1(n_390),
.B2(n_381),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_473),
.A2(n_479),
.B(n_436),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_427),
.A2(n_399),
.B1(n_390),
.B2(n_403),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_423),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_317),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_478),
.A2(n_440),
.B1(n_417),
.B2(n_425),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_435),
.B(n_430),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_481),
.A2(n_487),
.B(n_489),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_467),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_496),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_459),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_484),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_488),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_432),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_420),
.B(n_428),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_491),
.A2(n_495),
.B1(n_455),
.B2(n_464),
.Y(n_527)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_450),
.A2(n_419),
.B1(n_441),
.B2(n_414),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_448),
.A2(n_446),
.B(n_414),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_466),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_499),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_471),
.A2(n_429),
.B1(n_403),
.B2(n_395),
.Y(n_500)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_500),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_452),
.A2(n_395),
.B1(n_393),
.B2(n_399),
.Y(n_501)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_462),
.B(n_325),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_507),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_470),
.B(n_305),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_505),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_301),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_504),
.Y(n_529)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_457),
.Y(n_505)
);

OAI32xp33_ASAP7_75t_L g507 ( 
.A1(n_451),
.A2(n_393),
.A3(n_368),
.B1(n_340),
.B2(n_375),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_449),
.C(n_479),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_502),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_449),
.C(n_468),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_512),
.C(n_514),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_460),
.C(n_473),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_490),
.A2(n_458),
.B1(n_478),
.B2(n_461),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_513),
.A2(n_526),
.B1(n_522),
.B2(n_521),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_474),
.C(n_476),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_472),
.C(n_475),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_523),
.C(n_508),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_461),
.C(n_465),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_527),
.A2(n_505),
.B1(n_494),
.B2(n_480),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_489),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_531),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_490),
.A2(n_463),
.B(n_464),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_454),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_530),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_484),
.C(n_487),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_537),
.C(n_540),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_536),
.B(n_539),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_496),
.C(n_491),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_509),
.B(n_485),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_495),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_506),
.C(n_499),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_506),
.C(n_480),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_544),
.C(n_312),
.Y(n_566)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_515),
.Y(n_543)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_518),
.C(n_524),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_546),
.B1(n_547),
.B2(n_348),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_481),
.B1(n_493),
.B2(n_477),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_527),
.A2(n_493),
.B1(n_454),
.B2(n_507),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_515),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_548),
.Y(n_555)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

OAI321xp33_ASAP7_75t_L g556 ( 
.A1(n_549),
.A2(n_528),
.A3(n_521),
.B1(n_529),
.B2(n_525),
.C(n_522),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_550),
.B(n_551),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_517),
.B(n_352),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_552),
.A2(n_518),
.B1(n_520),
.B2(n_526),
.Y(n_554)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_556),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_558),
.B(n_566),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_544),
.A2(n_520),
.B1(n_513),
.B2(n_530),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_560),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_532),
.Y(n_560)
);

OAI321xp33_ASAP7_75t_L g563 ( 
.A1(n_541),
.A2(n_532),
.A3(n_516),
.B1(n_498),
.B2(n_456),
.C(n_397),
.Y(n_563)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_552),
.A2(n_516),
.B1(n_498),
.B2(n_397),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_564),
.A2(n_569),
.B1(n_550),
.B2(n_540),
.Y(n_572)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_565),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_542),
.A2(n_498),
.B1(n_297),
.B2(n_280),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_551),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_535),
.A2(n_326),
.B1(n_280),
.B2(n_312),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_572),
.B(n_557),
.Y(n_590)
);

MAJx2_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_534),
.C(n_533),
.Y(n_573)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_573),
.Y(n_586)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_574),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_554),
.A2(n_533),
.B1(n_280),
.B2(n_326),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_575),
.A2(n_555),
.B1(n_562),
.B2(n_561),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_326),
.C(n_301),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_569),
.C(n_564),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_309),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_579),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_559),
.A2(n_565),
.B(n_566),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_560),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_583),
.B(n_585),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_587),
.B(n_589),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_558),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_590),
.B(n_591),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_557),
.C(n_298),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_576),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_592),
.B(n_575),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_586),
.A2(n_585),
.B(n_570),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_593),
.B(n_597),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_595),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_590),
.B(n_582),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_588),
.B(n_582),
.C(n_580),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_598),
.B(n_581),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_600),
.A2(n_603),
.B(n_596),
.Y(n_604)
);

NOR2x1_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_591),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_604),
.A2(n_606),
.B1(n_571),
.B2(n_572),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_601),
.A2(n_596),
.B(n_599),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_605),
.A2(n_583),
.B(n_352),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_602),
.B(n_584),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_607),
.A2(n_608),
.B(n_352),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_282),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_282),
.B(n_300),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_611),
.A2(n_300),
.B1(n_325),
.B2(n_283),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_300),
.B(n_283),
.Y(n_613)
);


endmodule