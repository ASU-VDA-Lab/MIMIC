module fake_ariane_1309_n_1090 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_255, n_122, n_257, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1090);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_257;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1090;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_466;
wire n_756;
wire n_1016;
wire n_346;
wire n_940;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_851;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_193),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_170),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_90),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_221),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_159),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_91),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_172),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_146),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_252),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_111),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_104),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_188),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_101),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_14),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_72),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_131),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_11),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_125),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_99),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_129),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_43),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_145),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_183),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_5),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_45),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_216),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_179),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_238),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_107),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_41),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_71),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_178),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_32),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_21),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_79),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_244),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_92),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_86),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_66),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_140),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_55),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_255),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_134),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_248),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_284),
.Y(n_327)
);

BUFx2_ASAP7_75t_SL g328 ( 
.A(n_265),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_312),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_319),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_263),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_312),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_314),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_264),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_0),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_277),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_313),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_314),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_267),
.Y(n_345)
);

BUFx2_ASAP7_75t_SL g346 ( 
.A(n_265),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_277),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_272),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_273),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_274),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_321),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_265),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_313),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_313),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_321),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_326),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_266),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_276),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_281),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_329),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_285),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_345),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_R g377 ( 
.A(n_354),
.B(n_278),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_348),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_352),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_300),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_358),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_329),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_338),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_338),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_291),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_335),
.A2(n_287),
.B1(n_290),
.B2(n_297),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_342),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_359),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_347),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_347),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_268),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_360),
.B(n_268),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_360),
.B(n_292),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_362),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_306),
.Y(n_422)
);

AO21x2_ASAP7_75t_L g423 ( 
.A1(n_374),
.A2(n_322),
.B(n_318),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_302),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_362),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_280),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_398),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_302),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_375),
.B(n_302),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_282),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_0),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_375),
.B(n_310),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_310),
.B1(n_293),
.B2(n_295),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_286),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_383),
.B(n_299),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_304),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_305),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_307),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_308),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_391),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_376),
.B(n_311),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_417),
.B(n_416),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_407),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_371),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_407),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_418),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_402),
.B(n_1),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_386),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_408),
.B(n_381),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_381),
.B(n_315),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_372),
.Y(n_473)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_373),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_378),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_389),
.B(n_316),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_380),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_389),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_415),
.B1(n_411),
.B2(n_410),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_317),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_323),
.B(n_320),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

AND2x6_ASAP7_75t_SL g492 ( 
.A(n_469),
.B(n_339),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_443),
.B(n_324),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_464),
.A2(n_415),
.B1(n_411),
.B2(n_410),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_428),
.B(n_325),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_474),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_448),
.B(n_436),
.C(n_477),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_428),
.B(n_310),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_414),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_485),
.B(n_419),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_448),
.B(n_310),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_465),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_454),
.B(n_1),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_459),
.A2(n_344),
.B1(n_339),
.B2(n_371),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_438),
.B(n_2),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_2),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_430),
.A2(n_419),
.B1(n_344),
.B2(n_393),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_429),
.B(n_390),
.Y(n_513)
);

NAND2x1_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_49),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_483),
.A2(n_484),
.B1(n_461),
.B2(n_423),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_470),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_461),
.B(n_3),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_390),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_437),
.B(n_422),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_446),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_422),
.B(n_393),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_423),
.B(n_427),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_442),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_430),
.B(n_399),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_439),
.B(n_399),
.Y(n_527)
);

BUFx5_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_455),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_3),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_439),
.B(n_4),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_445),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_462),
.A2(n_436),
.B(n_433),
.C(n_426),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_471),
.B(n_423),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g536 ( 
.A(n_456),
.B(n_7),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_436),
.B(n_9),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_484),
.B(n_9),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_441),
.B(n_10),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_456),
.B(n_10),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_463),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_483),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_463),
.A2(n_480),
.B1(n_429),
.B2(n_457),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_440),
.B(n_15),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_479),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_425),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_457),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_440),
.B(n_452),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_440),
.B(n_15),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_429),
.B(n_16),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_452),
.B(n_16),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_481),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_424),
.B(n_17),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_452),
.B(n_17),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_424),
.B(n_18),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_467),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_544),
.A2(n_468),
.B1(n_476),
.B2(n_459),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_546),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_SL g563 ( 
.A(n_542),
.B(n_450),
.C(n_18),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_545),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_503),
.B(n_473),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_548),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_497),
.B(n_446),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_446),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_531),
.A2(n_421),
.B(n_435),
.C(n_431),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_519),
.A2(n_434),
.B1(n_420),
.B2(n_431),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_521),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_501),
.B(n_473),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_555),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_558),
.A2(n_476),
.B1(n_468),
.B2(n_421),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_549),
.B(n_524),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_435),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_SL g581 ( 
.A(n_542),
.B(n_19),
.C(n_20),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_532),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_495),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_525),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_SL g585 ( 
.A(n_505),
.B(n_19),
.C(n_20),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_488),
.B(n_498),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_513),
.B(n_449),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_517),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_546),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_558),
.A2(n_540),
.B1(n_527),
.B2(n_526),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_495),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_508),
.A2(n_453),
.B(n_449),
.C(n_473),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_513),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_513),
.B(n_453),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_420),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_534),
.B(n_420),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_509),
.B(n_420),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_520),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_522),
.B(n_475),
.Y(n_604)
);

AND3x1_ASAP7_75t_SL g605 ( 
.A(n_536),
.B(n_21),
.C(n_22),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_518),
.B(n_475),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_537),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_504),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_520),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_520),
.Y(n_611)
);

OR2x4_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_420),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_492),
.A2(n_475),
.B1(n_434),
.B2(n_482),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_525),
.B(n_434),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_511),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_486),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_489),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_494),
.B(n_434),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_541),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_516),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_434),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_570),
.A2(n_554),
.B(n_547),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_564),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_577),
.B(n_515),
.Y(n_625)
);

OAI21x1_ASAP7_75t_SL g626 ( 
.A1(n_588),
.A2(n_557),
.B(n_533),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_600),
.A2(n_596),
.B(n_514),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_603),
.B(n_543),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_593),
.A2(n_489),
.B1(n_496),
.B2(n_506),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_562),
.Y(n_631)
);

OA22x2_ASAP7_75t_L g632 ( 
.A1(n_616),
.A2(n_556),
.B1(n_552),
.B2(n_538),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_602),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_567),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_600),
.A2(n_535),
.B(n_523),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_621),
.A2(n_523),
.B(n_500),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_562),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_592),
.B(n_551),
.Y(n_638)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_563),
.A2(n_556),
.B(n_490),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_580),
.A2(n_528),
.B(n_482),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_567),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_570),
.A2(n_528),
.B(n_482),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_602),
.B(n_482),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_580),
.A2(n_528),
.B(n_482),
.Y(n_644)
);

O2A1O1Ixp5_ASAP7_75t_SL g645 ( 
.A1(n_608),
.A2(n_528),
.B(n_24),
.C(n_22),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_569),
.A2(n_528),
.B1(n_25),
.B2(n_23),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_569),
.A2(n_52),
.B(n_50),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_568),
.A2(n_54),
.B(n_53),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_616),
.B(n_23),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_24),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_25),
.Y(n_651)
);

NOR2x1_ASAP7_75t_L g652 ( 
.A(n_592),
.B(n_262),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_591),
.A2(n_26),
.B(n_27),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_594),
.B(n_56),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_568),
.B(n_26),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_579),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_611),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_589),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_604),
.B(n_28),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_614),
.A2(n_58),
.B(n_57),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_586),
.A2(n_60),
.B(n_59),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_586),
.A2(n_62),
.B(n_61),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

INVx3_ASAP7_75t_SL g665 ( 
.A(n_609),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

AO31x2_ASAP7_75t_L g667 ( 
.A1(n_587),
.A2(n_163),
.A3(n_258),
.B(n_257),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_593),
.A2(n_615),
.B(n_581),
.C(n_566),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_565),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_560),
.B(n_29),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_599),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_560),
.B(n_30),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_572),
.B(n_30),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_619),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_587),
.A2(n_64),
.B(n_63),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_571),
.A2(n_67),
.B(n_65),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

AOI211x1_ASAP7_75t_L g678 ( 
.A1(n_578),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_610),
.A2(n_69),
.B(n_68),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_590),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_629),
.B(n_573),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_597),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_670),
.A2(n_601),
.B1(n_618),
.B2(n_598),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_628),
.A2(n_610),
.B(n_575),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_677),
.B(n_613),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_624),
.B(n_594),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_624),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_640),
.A2(n_610),
.B(n_575),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_624),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_666),
.B(n_601),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_644),
.A2(n_584),
.B(n_561),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_622),
.A2(n_614),
.B(n_612),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_681),
.B(n_599),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_669),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_665),
.B(n_590),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_622),
.A2(n_618),
.B(n_559),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_671),
.Y(n_698)
);

OA21x2_ASAP7_75t_L g699 ( 
.A1(n_642),
.A2(n_576),
.B(n_559),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_642),
.A2(n_584),
.B(n_561),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_679),
.B(n_599),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_651),
.B(n_606),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_627),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_636),
.A2(n_576),
.B(n_583),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_623),
.Y(n_705)
);

AOI21xp33_ASAP7_75t_SL g706 ( 
.A1(n_674),
.A2(n_650),
.B(n_646),
.Y(n_706)
);

AO31x2_ASAP7_75t_L g707 ( 
.A1(n_630),
.A2(n_602),
.A3(n_612),
.B(n_620),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_634),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_641),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_668),
.B(n_607),
.Y(n_710)
);

AO31x2_ASAP7_75t_L g711 ( 
.A1(n_625),
.A2(n_620),
.A3(n_605),
.B(n_585),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_672),
.A2(n_598),
.B1(n_590),
.B2(n_614),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_657),
.B(n_598),
.Y(n_713)
);

AO21x2_ASAP7_75t_L g714 ( 
.A1(n_635),
.A2(n_595),
.B(n_611),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_646),
.A2(n_674),
.B1(n_653),
.B2(n_673),
.Y(n_715)
);

AO21x2_ASAP7_75t_L g716 ( 
.A1(n_626),
.A2(n_611),
.B(n_73),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_611),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_648),
.A2(n_34),
.A3(n_35),
.B(n_36),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_676),
.A2(n_74),
.B(n_70),
.Y(n_719)
);

OA21x2_ASAP7_75t_L g720 ( 
.A1(n_662),
.A2(n_76),
.B(n_75),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_675),
.A2(n_680),
.B(n_645),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_667),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_639),
.A2(n_78),
.B(n_77),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_671),
.B(n_35),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_660),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_631),
.B(n_36),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_631),
.B(n_37),
.Y(n_728)
);

AOI21x1_ASAP7_75t_L g729 ( 
.A1(n_632),
.A2(n_81),
.B(n_80),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_656),
.B(n_679),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_653),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_655),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_659),
.B(n_38),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_631),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_656),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_637),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_639),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_637),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_715),
.A2(n_637),
.B1(n_652),
.B2(n_656),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_682),
.B(n_658),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_690),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_715),
.A2(n_638),
.B1(n_633),
.B2(n_654),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_690),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_683),
.B(n_633),
.Y(n_744)
);

OAI222xp33_ASAP7_75t_L g745 ( 
.A1(n_731),
.A2(n_678),
.B1(n_661),
.B2(n_647),
.C1(n_667),
.C2(n_47),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_722),
.A2(n_643),
.B(n_667),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_733),
.A2(n_710),
.B1(n_697),
.B2(n_726),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_695),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_722),
.A2(n_643),
.B(n_678),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_703),
.Y(n_750)
);

AOI21xp33_ASAP7_75t_L g751 ( 
.A1(n_706),
.A2(n_42),
.B(n_44),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_733),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_730),
.B(n_46),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_R g754 ( 
.A(n_699),
.B(n_82),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_705),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_708),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_709),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_693),
.A2(n_47),
.B(n_48),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_736),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_SL g760 ( 
.A(n_710),
.B(n_48),
.C(n_83),
.Y(n_760)
);

AO21x2_ASAP7_75t_L g761 ( 
.A1(n_723),
.A2(n_84),
.B(n_85),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_730),
.B(n_87),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_697),
.A2(n_259),
.B1(n_89),
.B2(n_93),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_716),
.A2(n_88),
.B(n_94),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_702),
.B(n_95),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_707),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_732),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_737),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.C(n_106),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_736),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_703),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_690),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_730),
.Y(n_772)
);

AO21x2_ASAP7_75t_L g773 ( 
.A1(n_723),
.A2(n_108),
.B(n_112),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_699),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_698),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_725),
.B(n_116),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_721),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_687),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_684),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_696),
.B(n_256),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_727),
.B(n_120),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_734),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_721),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_688),
.B(n_121),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_716),
.A2(n_122),
.B(n_123),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_714),
.Y(n_786)
);

INVx4_ASAP7_75t_SL g787 ( 
.A(n_707),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_701),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_684),
.B(n_124),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_738),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_688),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_728),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_714),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_687),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_130),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_701),
.Y(n_796)
);

NAND4xp25_ASAP7_75t_L g797 ( 
.A(n_712),
.B(n_132),
.C(n_133),
.D(n_135),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_755),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_789),
.A2(n_691),
.B1(n_686),
.B2(n_712),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_756),
.Y(n_800)
);

INVx5_ASAP7_75t_L g801 ( 
.A(n_741),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_757),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_748),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_750),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_789),
.A2(n_691),
.B1(n_701),
.B2(n_694),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_744),
.B(n_717),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_752),
.B(n_717),
.C(n_698),
.Y(n_807)
);

BUFx5_ASAP7_75t_L g808 ( 
.A(n_791),
.Y(n_808)
);

OAI211xp5_ASAP7_75t_SL g809 ( 
.A1(n_752),
.A2(n_711),
.B(n_718),
.C(n_735),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_747),
.A2(n_691),
.B1(n_694),
.B2(n_729),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_797),
.A2(n_694),
.B1(n_699),
.B2(n_735),
.Y(n_811)
);

OAI211xp5_ASAP7_75t_L g812 ( 
.A1(n_751),
.A2(n_711),
.B(n_718),
.C(n_713),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_759),
.B(n_707),
.Y(n_813)
);

AOI21xp33_ASAP7_75t_L g814 ( 
.A1(n_754),
.A2(n_724),
.B(n_720),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_782),
.B(n_707),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_760),
.A2(n_724),
.B1(n_700),
.B2(n_720),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_775),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_750),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_SL g819 ( 
.A1(n_758),
.A2(n_711),
.B1(n_718),
.B2(n_700),
.C(n_685),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_753),
.B(n_711),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_747),
.A2(n_720),
.B1(n_718),
.B2(n_685),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_753),
.A2(n_692),
.B1(n_689),
.B2(n_719),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_760),
.A2(n_774),
.B1(n_776),
.B2(n_740),
.Y(n_824)
);

BUFx4f_ASAP7_75t_SL g825 ( 
.A(n_769),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_L g826 ( 
.A1(n_745),
.A2(n_719),
.B1(n_704),
.B2(n_139),
.C(n_141),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_739),
.A2(n_689),
.B1(n_692),
.B2(n_704),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_790),
.Y(n_828)
);

OA21x2_ASAP7_75t_L g829 ( 
.A1(n_746),
.A2(n_136),
.B(n_138),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_739),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_766),
.B(n_149),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_774),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_772),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_791),
.Y(n_834)
);

AOI221xp5_ASAP7_75t_L g835 ( 
.A1(n_745),
.A2(n_792),
.B1(n_765),
.B2(n_763),
.C(n_768),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_742),
.A2(n_153),
.B(n_154),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_770),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_770),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_766),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_792),
.A2(n_155),
.B(n_156),
.C(n_157),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_777),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_741),
.B(n_158),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_763),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_778),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_779),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_780),
.B(n_168),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_781),
.B(n_169),
.Y(n_847)
);

OAI221xp5_ASAP7_75t_L g848 ( 
.A1(n_784),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.C(n_175),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_787),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_798),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_813),
.B(n_787),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_806),
.B(n_787),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_828),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_815),
.B(n_777),
.Y(n_854)
);

INVx4_ASAP7_75t_R g855 ( 
.A(n_820),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_801),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_817),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_839),
.B(n_783),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_L g860 ( 
.A1(n_835),
.A2(n_824),
.B1(n_836),
.B2(n_809),
.C(n_840),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_802),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_803),
.B(n_783),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_804),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_825),
.B(n_743),
.Y(n_864)
);

OAI221xp5_ASAP7_75t_SL g865 ( 
.A1(n_812),
.A2(n_807),
.B1(n_826),
.B2(n_811),
.C(n_832),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_838),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_844),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_801),
.B(n_741),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_841),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_821),
.B(n_786),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_819),
.B(n_786),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_818),
.B(n_793),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_831),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_829),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_807),
.B(n_793),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_819),
.B(n_823),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_823),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_827),
.B(n_816),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_810),
.A2(n_761),
.B1(n_773),
.B2(n_795),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_834),
.B(n_743),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_808),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_833),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_808),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_808),
.Y(n_887)
);

NOR2x1_ASAP7_75t_L g888 ( 
.A(n_833),
.B(n_771),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_801),
.B(n_741),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_808),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_808),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_805),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_836),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_814),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_822),
.B(n_749),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_822),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_822),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_799),
.B(n_771),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_846),
.B(n_796),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_848),
.A2(n_785),
.B(n_764),
.C(n_762),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_842),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_830),
.B(n_788),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_830),
.B(n_788),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_845),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_843),
.B(n_761),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_828),
.B(n_778),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_867),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_853),
.B(n_773),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_880),
.B(n_878),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_880),
.B(n_762),
.Y(n_912)
);

AOI221xp5_ASAP7_75t_L g913 ( 
.A1(n_860),
.A2(n_767),
.B1(n_794),
.B2(n_754),
.C(n_185),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_857),
.Y(n_914)
);

OAI221xp5_ASAP7_75t_SL g915 ( 
.A1(n_878),
.A2(n_794),
.B1(n_182),
.B2(n_184),
.C(n_186),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_879),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_863),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_879),
.B(n_181),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_895),
.B(n_187),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_906),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_863),
.Y(n_921)
);

NOR4xp25_ASAP7_75t_SL g922 ( 
.A(n_865),
.B(n_192),
.C(n_194),
.D(n_195),
.Y(n_922)
);

OAI221xp5_ASAP7_75t_L g923 ( 
.A1(n_893),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.C(n_199),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_850),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_866),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_874),
.B(n_200),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_850),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_872),
.B(n_201),
.Y(n_928)
);

OAI33xp33_ASAP7_75t_L g929 ( 
.A1(n_894),
.A2(n_202),
.A3(n_203),
.B1(n_204),
.B2(n_205),
.B3(n_206),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_861),
.B(n_207),
.Y(n_930)
);

AOI33xp33_ASAP7_75t_L g931 ( 
.A1(n_893),
.A2(n_872),
.A3(n_861),
.B1(n_894),
.B2(n_881),
.B3(n_871),
.Y(n_931)
);

OAI211xp5_ASAP7_75t_L g932 ( 
.A1(n_905),
.A2(n_208),
.B(n_209),
.C(n_210),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_870),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_870),
.Y(n_934)
);

OAI321xp33_ASAP7_75t_L g935 ( 
.A1(n_907),
.A2(n_211),
.A3(n_213),
.B1(n_214),
.B2(n_215),
.C(n_217),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_882),
.A2(n_218),
.B(n_219),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_854),
.B(n_220),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_869),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_866),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_895),
.B(n_222),
.Y(n_940)
);

AOI221xp5_ASAP7_75t_L g941 ( 
.A1(n_871),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_906),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_867),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_916),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_910),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_911),
.B(n_885),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_933),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_934),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_911),
.B(n_908),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_914),
.B(n_858),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_938),
.B(n_869),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_909),
.B(n_864),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_927),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_910),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_938),
.B(n_884),
.Y(n_956)
);

AND2x4_ASAP7_75t_SL g957 ( 
.A(n_912),
.B(n_889),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_938),
.B(n_884),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_912),
.B(n_909),
.Y(n_959)
);

NOR2x1p5_ASAP7_75t_L g960 ( 
.A(n_943),
.B(n_903),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_931),
.Y(n_961)
);

NAND2x1_ASAP7_75t_L g962 ( 
.A(n_912),
.B(n_855),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_912),
.B(n_891),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_943),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_918),
.B(n_858),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_931),
.B(n_898),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_918),
.B(n_859),
.Y(n_967)
);

NAND2x1_ASAP7_75t_SL g968 ( 
.A(n_928),
.B(n_888),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_917),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_928),
.B(n_891),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_917),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_921),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_919),
.B(n_896),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_947),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_968),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_947),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_948),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_966),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_970),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_948),
.Y(n_980)
);

NOR3x1_ASAP7_75t_L g981 ( 
.A(n_961),
.B(n_896),
.C(n_926),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_957),
.B(n_919),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_954),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_961),
.A2(n_932),
.B(n_935),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_950),
.B(n_898),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_950),
.B(n_862),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_944),
.B(n_875),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_954),
.Y(n_988)
);

XNOR2x1_ASAP7_75t_L g989 ( 
.A(n_967),
.B(n_937),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_949),
.B(n_862),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_984),
.A2(n_962),
.B(n_959),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_978),
.A2(n_913),
.B1(n_929),
.B2(n_936),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_R g993 ( 
.A(n_982),
.B(n_964),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_989),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_984),
.A2(n_915),
.B(n_959),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_990),
.B(n_949),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_982),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_975),
.B(n_964),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_981),
.B(n_946),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_974),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_976),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_977),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_992),
.A2(n_936),
.B1(n_907),
.B2(n_941),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_994),
.B(n_995),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_993),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_993),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_997),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_946),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1000),
.B(n_980),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_1004),
.A2(n_998),
.B(n_991),
.Y(n_1011)
);

NAND2x1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.B(n_1001),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1007),
.Y(n_1014)
);

OAI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_1003),
.A2(n_992),
.B1(n_955),
.B2(n_945),
.C(n_967),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_1003),
.A2(n_1002),
.B(n_902),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1014),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_1011),
.B(n_1005),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_1008),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_1012),
.Y(n_1020)
);

AOI211xp5_ASAP7_75t_L g1021 ( 
.A1(n_1016),
.A2(n_1009),
.B(n_923),
.C(n_901),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_1018),
.B(n_1015),
.C(n_922),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_940),
.C(n_919),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_1020),
.B(n_940),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_1021),
.B(n_952),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_1017),
.B(n_987),
.Y(n_1026)
);

AND2x4_ASAP7_75t_SL g1027 ( 
.A(n_1019),
.B(n_951),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1020),
.A2(n_987),
.B(n_988),
.Y(n_1028)
);

OAI22xp33_ASAP7_75t_SL g1029 ( 
.A1(n_1024),
.A2(n_945),
.B1(n_955),
.B2(n_965),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_1022),
.Y(n_1030)
);

AOI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_1026),
.A2(n_882),
.B1(n_983),
.B2(n_876),
.C(n_936),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_1028),
.A2(n_876),
.B1(n_930),
.B2(n_902),
.C(n_953),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1027),
.B(n_979),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1025),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1030),
.A2(n_1023),
.B1(n_920),
.B2(n_942),
.C(n_940),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_1033),
.B(n_951),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1031),
.A2(n_960),
.B1(n_970),
.B2(n_937),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1029),
.Y(n_1039)
);

AOI221xp5_ASAP7_75t_L g1040 ( 
.A1(n_1032),
.A2(n_900),
.B1(n_965),
.B2(n_899),
.C(n_972),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1034),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_1041),
.B(n_883),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_1039),
.B(n_886),
.C(n_887),
.Y(n_1044)
);

AND4x1_ASAP7_75t_L g1045 ( 
.A(n_1036),
.B(n_973),
.C(n_963),
.D(n_888),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1037),
.B(n_973),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1038),
.B(n_986),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

AOI221xp5_ASAP7_75t_L g1049 ( 
.A1(n_1039),
.A2(n_971),
.B1(n_969),
.B2(n_985),
.C(n_963),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1035),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1042),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_1048),
.A2(n_957),
.B1(n_897),
.B2(n_856),
.Y(n_1052)
);

NAND4xp75_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_956),
.C(n_958),
.D(n_887),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1046),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_1044),
.A2(n_971),
.B1(n_969),
.B2(n_956),
.C(n_958),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1049),
.A2(n_892),
.B1(n_897),
.B2(n_875),
.Y(n_1056)
);

NAND4xp25_ASAP7_75t_L g1057 ( 
.A(n_1047),
.B(n_1043),
.C(n_1045),
.D(n_886),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_1042),
.B(n_962),
.C(n_904),
.Y(n_1058)
);

NOR4xp25_ASAP7_75t_L g1059 ( 
.A(n_1042),
.B(n_904),
.C(n_890),
.D(n_968),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1042),
.B(n_892),
.C(n_877),
.Y(n_1060)
);

OAI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1044),
.A2(n_890),
.B1(n_877),
.B2(n_856),
.C(n_939),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_1042),
.B(n_852),
.C(n_851),
.Y(n_1062)
);

OAI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1042),
.A2(n_856),
.B(n_852),
.C(n_851),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_1051),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1054),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1062),
.Y(n_1066)
);

XNOR2xp5_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_889),
.Y(n_1067)
);

CKINVDCx12_ASAP7_75t_R g1068 ( 
.A(n_1052),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_1063),
.B(n_856),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1053),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1059),
.Y(n_1071)
);

AO22x2_ASAP7_75t_L g1072 ( 
.A1(n_1065),
.A2(n_1060),
.B1(n_1058),
.B2(n_1056),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1066),
.Y(n_1073)
);

OA21x2_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_1055),
.B(n_868),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1066),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_SL g1076 ( 
.A1(n_1073),
.A2(n_1068),
.B1(n_1067),
.B2(n_1069),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1075),
.A2(n_856),
.B1(n_889),
.B2(n_868),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1071),
.A2(n_939),
.B(n_925),
.Y(n_1078)
);

OAI22x1_ASAP7_75t_L g1079 ( 
.A1(n_1074),
.A2(n_1072),
.B1(n_889),
.B2(n_868),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_925),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_854),
.Y(n_1081)
);

AOI222xp33_ASAP7_75t_L g1082 ( 
.A1(n_1081),
.A2(n_1076),
.B1(n_1077),
.B2(n_921),
.C1(n_233),
.C2(n_234),
.Y(n_1082)
);

XNOR2xp5_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_230),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1081),
.A2(n_231),
.B(n_232),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_235),
.B(n_236),
.Y(n_1085)
);

AOI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1083),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.C1(n_241),
.C2(n_242),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1086),
.A2(n_1082),
.B1(n_873),
.B2(n_855),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1085),
.Y(n_1088)
);

OAI221xp5_ASAP7_75t_R g1089 ( 
.A1(n_1087),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.C(n_247),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_1088),
.B(n_249),
.C(n_251),
.Y(n_1090)
);


endmodule