module real_jpeg_6521_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_1),
.Y(n_177)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_2),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_3),
.A2(n_72),
.B1(n_132),
.B2(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_3),
.A2(n_132),
.B1(n_280),
.B2(n_315),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_3),
.A2(n_132),
.B1(n_384),
.B2(n_386),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_56),
.B1(n_59),
.B2(n_61),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_61),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_4),
.A2(n_61),
.B1(n_288),
.B2(n_355),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_5),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_5),
.A2(n_66),
.B1(n_90),
.B2(n_229),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_6),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_10),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_10),
.A2(n_205),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_10),
.B(n_270),
.C(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_10),
.B(n_110),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_10),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_10),
.B(n_63),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_10),
.B(n_124),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_12),
.A2(n_130),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_12),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_120),
.B1(n_157),
.B2(n_220),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_12),
.A2(n_157),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_12),
.A2(n_157),
.B1(n_266),
.B2(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_77),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_15),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_15),
.A2(n_69),
.B1(n_75),
.B2(n_180),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_15),
.A2(n_69),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_16),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_16),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_16),
.A2(n_118),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_16),
.A2(n_41),
.B1(n_67),
.B2(n_118),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_16),
.A2(n_118),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_245),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_244),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_223),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_21),
.B(n_223),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_163),
.C(n_181),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_22),
.A2(n_23),
.B1(n_163),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_94),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_24),
.B(n_95),
.C(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_73),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_25),
.B(n_73),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_55),
.B1(n_62),
.B2(n_64),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_26),
.A2(n_254),
.B(n_261),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_26),
.A2(n_62),
.B1(n_294),
.B2(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_26),
.A2(n_261),
.B(n_340),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_63),
.B1(n_65),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_27),
.A2(n_63),
.B1(n_165),
.B2(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_27),
.B(n_262),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_44),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_30),
.Y(n_166)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_32),
.Y(n_168)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_32),
.Y(n_231)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_33),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_33),
.Y(n_341)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_45),
.B1(n_49),
.B2(n_52),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_44),
.A2(n_294),
.B(n_298),
.Y(n_293)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_47),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_47),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_51),
.Y(n_356)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_54),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_55),
.A2(n_62),
.B(n_298),
.Y(n_411)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_68),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_63),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_80),
.B1(n_87),
.B2(n_92),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_74),
.Y(n_216)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_76),
.Y(n_290)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_78),
.Y(n_278)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_80),
.B(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_80),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_80),
.A2(n_172),
.B1(n_213),
.B2(n_354),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_85),
.Y(n_288)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_86),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_86),
.Y(n_317)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_88),
.A2(n_170),
.B1(n_171),
.B2(n_176),
.Y(n_169)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_128),
.B1(n_161),
.B2(n_162),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_95),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_110),
.B1(n_114),
.B2(n_122),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_96),
.A2(n_218),
.B(n_221),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_96),
.A2(n_221),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_96),
.B(n_114),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_97),
.A2(n_123),
.B1(n_222),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_97),
.A2(n_219),
.B1(n_222),
.B2(n_383),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_109),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_103),
.Y(n_365)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_103),
.Y(n_372)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_107),
.Y(n_240)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_108),
.Y(n_348)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_108),
.Y(n_388)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_115),
.B(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_136),
.B1(n_156),
.B2(n_159),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_159),
.B(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_136),
.A2(n_156),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_137),
.A2(n_407),
.B(n_408),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_141),
.Y(n_198)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_152),
.B2(n_154),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_159),
.B(n_205),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_163),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_169),
.Y(n_235)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_212),
.B1(n_214),
.B2(n_216),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_170),
.A2(n_173),
.B(n_176),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_170),
.A2(n_276),
.B(n_283),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_170),
.A2(n_205),
.B(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_175),
.Y(n_329)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_181),
.B(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.C(n_217),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_182),
.A2(n_183),
.B1(n_217),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_SL g407 ( 
.A1(n_186),
.A2(n_204),
.B(n_205),
.Y(n_407)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_189),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_210),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_190),
.A2(n_210),
.B1(n_211),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_190),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_193),
.A3(n_197),
.B1(n_199),
.B2(n_204),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_205),
.A2(n_345),
.B(n_349),
.Y(n_344)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_217),
.Y(n_421)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI32xp33_ASAP7_75t_L g359 ( 
.A1(n_220),
.A2(n_350),
.A3(n_360),
.B1(n_362),
.B2(n_366),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_222),
.A2(n_383),
.B(n_389),
.Y(n_382)
);

BUFx24_ASAP7_75t_SL g437 ( 
.A(n_223),
.Y(n_437)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.CI(n_234),
.CON(n_223),
.SN(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_243),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_414),
.B(n_433),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_395),
.B(n_413),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_374),
.B(n_394),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_334),
.B(n_373),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_301),
.B(n_333),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_274),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_274),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_253),
.A2(n_263),
.B1(n_264),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_260),
.Y(n_361)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_260),
.Y(n_369)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_291),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_292),
.C(n_300),
.Y(n_335)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_299),
.B2(n_300),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_324),
.B(n_332),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_312),
.B(n_323),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_311),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_322),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_318),
.B(n_321),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_353),
.B(n_357),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_330),
.Y(n_332)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_336),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_351),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_342),
.C(n_351),
.Y(n_375)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_359),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_375),
.B(n_376),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_393),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_380),
.C(n_393),
.Y(n_396)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_390),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_391),
.C(n_392),
.Y(n_401)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_397),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_398)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_401),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_402),
.C(n_404),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_409),
.B2(n_412),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_410),
.C(n_411),
.Y(n_424)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_409),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_428),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_417),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_425),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.C(n_424),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_422),
.A2(n_423),
.B1(n_424),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_430),
.Y(n_434)
);


endmodule