module fake_jpeg_27780_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_34),
.B1(n_27),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_24),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_64),
.B1(n_65),
.B2(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_34),
.B1(n_21),
.B2(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_17),
.B1(n_22),
.B2(n_29),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_66),
.B(n_67),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_70),
.B1(n_97),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_32),
.B1(n_20),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_79),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_84),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_33),
.B1(n_19),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_58),
.B1(n_50),
.B2(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_98),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_16),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_0),
.Y(n_132)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_35),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_65),
.B1(n_63),
.B2(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_103),
.Y(n_120)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_58),
.B1(n_50),
.B2(n_59),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_48),
.B1(n_36),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_121),
.B1(n_102),
.B2(n_103),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_36),
.B1(n_33),
.B2(n_19),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_81),
.B1(n_80),
.B2(n_86),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_33),
.B1(n_19),
.B2(n_36),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_30),
.C(n_33),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_69),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_76),
.B(n_82),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_147),
.B1(n_126),
.B2(n_127),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_157),
.B1(n_159),
.B2(n_165),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_93),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_140),
.B(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_137),
.B(n_138),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_67),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_87),
.B(n_79),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_71),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_144),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_151),
.Y(n_199)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_115),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_92),
.B(n_95),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_70),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_111),
.B1(n_106),
.B2(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_160),
.B1(n_131),
.B2(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_100),
.B(n_104),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_26),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_90),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_125),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_185),
.B1(n_187),
.B2(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_107),
.C(n_128),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_173),
.C(n_184),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_177),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_117),
.C(n_129),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_117),
.B(n_129),
.C(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_176),
.B(n_178),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_2),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_131),
.C(n_119),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_135),
.A2(n_114),
.B1(n_85),
.B2(n_83),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_114),
.B1(n_85),
.B2(n_83),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_73),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_198),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_133),
.B1(n_84),
.B2(n_89),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_150),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_72),
.B1(n_68),
.B2(n_31),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_68),
.B1(n_31),
.B2(n_16),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_139),
.B(n_16),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_204),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_136),
.C(n_148),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_207),
.C(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_198),
.B1(n_151),
.B2(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_208),
.B(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_154),
.C(n_165),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_177),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_68),
.C(n_31),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_68),
.C(n_15),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_220),
.C(n_196),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_223),
.B(n_176),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_14),
.C(n_13),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_221),
.B1(n_214),
.B2(n_195),
.Y(n_233)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_14),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_231),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_200),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_182),
.B(n_175),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_225),
.C(n_203),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_243),
.C(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_166),
.B1(n_185),
.B2(n_193),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_242),
.B1(n_219),
.B2(n_213),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_201),
.B1(n_204),
.B2(n_212),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_189),
.C(n_182),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_167),
.B1(n_191),
.B2(n_168),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_169),
.C(n_171),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_250),
.C(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_181),
.C(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_261),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_263),
.C(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_217),
.C(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_218),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_216),
.C(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_239),
.B1(n_235),
.B2(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_247),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_229),
.C(n_249),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_282),
.C(n_266),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_268),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_254),
.C(n_229),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_243),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_287),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_271),
.B1(n_261),
.B2(n_257),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_288),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_246),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_254),
.B(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

OAI221xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_265),
.B1(n_252),
.B2(n_232),
.C(n_260),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_298),
.B(n_5),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_282),
.C(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_267),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_247),
.B(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_302),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_3),
.B(n_4),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_5),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_305),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_286),
.B(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_312),
.C(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_310),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_283),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_288),
.C(n_289),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_298),
.C(n_7),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_6),
.C(n_7),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_6),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_311),
.B(n_306),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_314),
.B(n_315),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.C(n_8),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_9),
.B(n_6),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_6),
.B(n_8),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_8),
.Y(n_330)
);


endmodule