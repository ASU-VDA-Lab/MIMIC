module fake_jpeg_30503_n_527 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_6),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_61),
.B(n_85),
.Y(n_138)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_29),
.B(n_6),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_6),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_99),
.B(n_104),
.Y(n_166)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_12),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_15),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_106),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_41),
.B1(n_27),
.B2(n_46),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_111),
.A2(n_112),
.B1(n_133),
.B2(n_136),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_41),
.B1(n_27),
.B2(n_46),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_61),
.A2(n_37),
.B1(n_29),
.B2(n_44),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_114),
.B(n_164),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_30),
.B1(n_53),
.B2(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_118),
.A2(n_132),
.B1(n_158),
.B2(n_53),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_53),
.B1(n_32),
.B2(n_36),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_37),
.B1(n_25),
.B2(n_36),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_65),
.A2(n_25),
.B1(n_36),
.B2(n_32),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_69),
.A2(n_25),
.B1(n_36),
.B2(n_32),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_107),
.B1(n_84),
.B2(n_78),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_96),
.A2(n_53),
.B1(n_25),
.B2(n_32),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_98),
.A2(n_24),
.B(n_52),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_100),
.B(n_24),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_48),
.Y(n_177)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_177),
.Y(n_225)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_119),
.Y(n_174)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_178),
.A2(n_201),
.B1(n_202),
.B2(n_215),
.Y(n_235)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_90),
.B1(n_91),
.B2(n_76),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_182),
.A2(n_197),
.B1(n_209),
.B2(n_223),
.Y(n_251)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_196),
.B1(n_158),
.B2(n_132),
.Y(n_245)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_193),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_138),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_194),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_136),
.B1(n_138),
.B2(n_117),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_67),
.B1(n_66),
.B2(n_57),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_18),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_203),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_131),
.A2(n_50),
.B1(n_52),
.B2(n_45),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_146),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_150),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_152),
.B(n_49),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_206),
.B(n_207),
.Y(n_263)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

NAND2x1_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_214),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_139),
.A2(n_54),
.B1(n_35),
.B2(n_47),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_18),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_224),
.C(n_33),
.Y(n_231)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_48),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_148),
.A2(n_47),
.B1(n_35),
.B2(n_40),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_222),
.B1(n_161),
.B2(n_135),
.Y(n_255)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_126),
.A2(n_47),
.B1(n_35),
.B2(n_40),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_18),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_49),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_243),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_44),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_230),
.B(n_240),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_18),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_194),
.B(n_153),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_200),
.B(n_159),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_261),
.B1(n_210),
.B2(n_224),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_126),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_129),
.Y(n_247)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_196),
.B(n_156),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_192),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_180),
.A2(n_189),
.B1(n_208),
.B2(n_210),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_180),
.A2(n_156),
.B1(n_160),
.B2(n_170),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_143),
.B1(n_174),
.B2(n_144),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_265),
.A2(n_274),
.B1(n_294),
.B2(n_228),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_268),
.A2(n_272),
.B1(n_290),
.B2(n_238),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_204),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_271),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_224),
.B1(n_185),
.B2(n_183),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_170),
.B1(n_144),
.B2(n_145),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_236),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_243),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_277),
.C(n_291),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_175),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_222),
.B(n_207),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_281),
.B(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_228),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_283),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_188),
.B(n_212),
.Y(n_281)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_235),
.A2(n_199),
.B1(n_145),
.B2(n_160),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_285),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_239),
.A2(n_124),
.B1(n_219),
.B2(n_218),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_240),
.A2(n_176),
.B1(n_191),
.B2(n_184),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_190),
.C(n_154),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_226),
.A2(n_186),
.B(n_179),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_181),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_297),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_247),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_15),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_296),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_251),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_293),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_298),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_231),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_303),
.C(n_278),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_246),
.C(n_230),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_228),
.Y(n_305)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_292),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_307),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_312),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_266),
.B(n_225),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_229),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_321),
.B(n_322),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

FAx1_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_263),
.CI(n_236),
.CON(n_323),
.SN(n_323)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_275),
.B(n_296),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_274),
.B1(n_287),
.B2(n_297),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_229),
.Y(n_325)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_326),
.B(n_328),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_263),
.B(n_241),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_328),
.A2(n_285),
.B(n_265),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_330),
.A2(n_339),
.B1(n_306),
.B2(n_348),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_323),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_291),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_303),
.Y(n_359)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_287),
.B1(n_266),
.B2(n_282),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_358),
.B1(n_317),
.B2(n_324),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_351),
.C(n_354),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_280),
.B(n_273),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_340),
.A2(n_341),
.B(n_342),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_318),
.A2(n_284),
.B(n_253),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_282),
.B(n_294),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_299),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_311),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_348),
.A2(n_356),
.B(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_244),
.Y(n_351)
);

OAI32xp33_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_256),
.A3(n_253),
.B1(n_264),
.B2(n_271),
.Y(n_352)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_244),
.C(n_258),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_258),
.C(n_232),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_300),
.C(n_323),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_305),
.A2(n_328),
.B(n_307),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_305),
.A2(n_232),
.B(n_288),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_256),
.B1(n_283),
.B2(n_289),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_387),
.C(n_351),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_325),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_361),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_325),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_338),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_366),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_368),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_308),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_303),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_349),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_301),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_375),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_335),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_313),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_377),
.B(n_381),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_324),
.B1(n_298),
.B2(n_323),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_379),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_301),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_339),
.A2(n_309),
.B1(n_300),
.B2(n_305),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_380),
.A2(n_323),
.B(n_311),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_335),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_385),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_344),
.B(n_321),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_386),
.A2(n_329),
.B1(n_358),
.B2(n_346),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_389),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_349),
.B(n_327),
.Y(n_389)
);

BUFx12_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_392),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_379),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_394),
.B(n_370),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_383),
.A2(n_356),
.B(n_347),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_396),
.B(n_397),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_398),
.A2(n_410),
.B1(n_396),
.B2(n_415),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_354),
.C(n_340),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_374),
.C(n_377),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_405),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_381),
.B(n_341),
.CI(n_344),
.CON(n_404),
.SN(n_404)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_346),
.B(n_345),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_406),
.A2(n_378),
.B1(n_365),
.B2(n_387),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_364),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_408),
.A2(n_414),
.B1(n_416),
.B2(n_319),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_383),
.A2(n_331),
.B(n_329),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_412),
.B(n_418),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_331),
.B(n_345),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_369),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_342),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_314),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_369),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_372),
.B1(n_360),
.B2(n_380),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_376),
.A2(n_357),
.B(n_331),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_361),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_420),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_421),
.A2(n_398),
.B1(n_403),
.B2(n_399),
.Y(n_450)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_429),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_435),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_439),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_SL g428 ( 
.A1(n_411),
.A2(n_372),
.B(n_330),
.C(n_315),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_412),
.B(n_400),
.C(n_395),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_384),
.C(n_314),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_410),
.A2(n_384),
.B1(n_353),
.B2(n_311),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_418),
.B1(n_416),
.B2(n_414),
.Y(n_444)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_440),
.Y(n_458)
);

XNOR2x1_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_401),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_327),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_397),
.A2(n_362),
.B(n_319),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_437),
.B(n_413),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_400),
.A2(n_319),
.B1(n_304),
.B2(n_286),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_408),
.B1(n_391),
.B2(n_402),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_446),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_444),
.A2(n_436),
.B1(n_428),
.B2(n_432),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_409),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_447),
.A2(n_310),
.B(n_259),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_455),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_452),
.B1(n_457),
.B2(n_459),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_409),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_453),
.C(n_426),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_395),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_423),
.A2(n_407),
.B1(n_404),
.B2(n_304),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g456 ( 
.A(n_424),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_259),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_422),
.A2(n_404),
.B1(n_392),
.B2(n_286),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_438),
.A2(n_392),
.B1(n_233),
.B2(n_237),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_467),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_430),
.B(n_439),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_464),
.A2(n_473),
.B(n_476),
.Y(n_478)
);

AO21x1_ASAP7_75t_L g465 ( 
.A1(n_458),
.A2(n_430),
.B(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_460),
.B(n_443),
.C(n_450),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_234),
.B(n_249),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_442),
.A2(n_432),
.B1(n_428),
.B2(n_427),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_442),
.A2(n_431),
.B1(n_429),
.B2(n_420),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_392),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_472),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_447),
.B(n_237),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_254),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_259),
.C(n_234),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_453),
.A2(n_451),
.B1(n_448),
.B2(n_446),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_242),
.B1(n_227),
.B2(n_234),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_249),
.B1(n_242),
.B2(n_310),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_479),
.A2(n_478),
.B1(n_482),
.B2(n_480),
.Y(n_504)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_310),
.CI(n_227),
.CON(n_481),
.SN(n_481)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_310),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_485),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_242),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_488),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_471),
.A2(n_227),
.B(n_252),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_487),
.A2(n_473),
.B1(n_254),
.B2(n_465),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_462),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_254),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_485),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_494),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_490),
.B(n_484),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_499),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_491),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_467),
.B1(n_475),
.B2(n_463),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_479),
.C(n_15),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_475),
.B1(n_7),
.B2(n_8),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_504),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_481),
.A2(n_7),
.B(n_12),
.C(n_10),
.Y(n_503)
);

NOR2x1p5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_7),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_499),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_498),
.Y(n_513)
);

OAI321xp33_ASAP7_75t_L g514 ( 
.A1(n_507),
.A2(n_503),
.A3(n_505),
.B1(n_509),
.B2(n_500),
.C(n_512),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_498),
.B(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_508),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_497),
.C(n_501),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_514),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_496),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_516),
.A2(n_507),
.B(n_15),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_7),
.C(n_8),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_519),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_520),
.A2(n_515),
.B(n_2),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

A2O1A1O1Ixp25_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_521),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_0),
.B(n_3),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_5),
.B1(n_507),
.B2(n_523),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_5),
.Y(n_527)
);


endmodule