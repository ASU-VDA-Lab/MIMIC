module real_jpeg_12563_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_2),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_14),
.C(n_30),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_5),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_12)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_17),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_34),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_26),
.B(n_33),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_24),
.Y(n_8)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_12),
.B(n_18),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_10),
.A2(n_12),
.B1(n_20),
.B2(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_14),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_21),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_39),
.B(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_46),
.Y(n_45)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_51),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);


endmodule