module fake_jpeg_10330_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_2),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_2),
.B1(n_3),
.B2(n_1),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_18),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_4),
.C(n_5),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_22),
.C(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx9p33_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_13),
.B1(n_9),
.B2(n_8),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_9),
.B1(n_13),
.B2(n_8),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_8),
.B1(n_28),
.B2(n_24),
.Y(n_35)
);

XOR2x1_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_12),
.Y(n_28)
);

XOR2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_20),
.B(n_16),
.Y(n_32)
);

BUFx24_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_9),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI31xp67_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_24),
.A3(n_34),
.B(n_39),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.C(n_37),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_24),
.Y(n_42)
);


endmodule