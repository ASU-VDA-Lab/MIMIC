module fake_jpeg_31144_n_156 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_156);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_26),
.B1(n_18),
.B2(n_22),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_26),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_48),
.B1(n_30),
.B2(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_60),
.Y(n_77)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_29),
.Y(n_87)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

XOR2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_46),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_74),
.C(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_80),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_43),
.B1(n_37),
.B2(n_23),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_50),
.B(n_51),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_14),
.C(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_29),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_55),
.B1(n_64),
.B2(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_30),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_91),
.B(n_101),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_21),
.B(n_23),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_53),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_91),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_23),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_74),
.C(n_77),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_102),
.B1(n_81),
.B2(n_75),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_21),
.B1(n_59),
.B2(n_4),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_71),
.B1(n_78),
.B2(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_101),
.C(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_92),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_84),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_69),
.B1(n_71),
.B2(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_101),
.B(n_106),
.Y(n_121)
);

AOI21x1_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_119),
.B(n_113),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_99),
.A3(n_93),
.B1(n_97),
.B2(n_11),
.C1(n_9),
.C2(n_10),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_10),
.C(n_119),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_126),
.C(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_95),
.C(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_104),
.B1(n_102),
.B2(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_133),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_115),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_121),
.B(n_127),
.C(n_120),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_107),
.C(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_75),
.B1(n_125),
.B2(n_129),
.Y(n_143)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_124),
.Y(n_140)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_136),
.B(n_92),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_142),
.B(n_138),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_120),
.A3(n_122),
.B1(n_129),
.B2(n_125),
.C1(n_108),
.C2(n_111),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_5),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_146),
.B(n_140),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_135),
.B(n_144),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_141),
.B(n_59),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_151),
.B(n_141),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_153),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_59),
.Y(n_156)
);


endmodule