module real_jpeg_15510_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_0),
.A2(n_6),
.B1(n_41),
.B2(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_0),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_0),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_0),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_0),
.B(n_141),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_0),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_0),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_0),
.B(n_104),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_1),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_1),
.B(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_2),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_2),
.B(n_122),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_5),
.Y(n_98)
);

AND2x4_ASAP7_75t_SL g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_6),
.B(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_6),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_7),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_7),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_7),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_7),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_7),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_7),
.B(n_353),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

NAND2x1_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_10),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_36),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_11),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_11),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_11),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_11),
.B(n_402),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_12),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_12),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_12),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_12),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_12),
.B(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_13),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_13),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_391),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_215),
.B(n_390),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_172),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_20),
.B(n_172),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_21),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_61),
.C(n_83),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_23),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.C(n_49),
.Y(n_23)
);

XNOR2x2_ASAP7_75t_L g269 ( 
.A(n_24),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_32),
.C(n_35),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_27),
.B(n_163),
.Y(n_426)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_39),
.A2(n_40),
.B1(n_49),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_40),
.A2(n_237),
.B(n_243),
.Y(n_236)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_44),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_48),
.Y(n_165)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_49),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_58),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_51),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_50),
.A2(n_51),
.B1(n_58),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g427 ( 
.A(n_51),
.B(n_97),
.C(n_103),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_55),
.B(n_186),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_57),
.Y(n_421)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_61),
.A2(n_83),
.B1(n_84),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.C(n_79),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.C(n_70),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_63),
.B(n_67),
.C(n_70),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_63),
.B(n_70),
.Y(n_249)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_63),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_66),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_67),
.B(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_73),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_81),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_82),
.Y(n_406)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_85),
.B(n_87),
.C(n_91),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_87),
.A2(n_88),
.B1(n_230),
.B2(n_231),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_88),
.B(n_223),
.C(n_230),
.Y(n_222)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_130),
.B1(n_170),
.B2(n_171),
.Y(n_92)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_93),
.B(n_171),
.C(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_94),
.B(n_108),
.C(n_116),
.Y(n_431)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_97),
.A2(n_106),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_98),
.B(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_100),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_103),
.B1(n_113),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_109),
.C(n_113),
.Y(n_108)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_114),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_117),
.B(n_121),
.C(n_125),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_119),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_128),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_158),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_131),
.B(n_159),
.C(n_160),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_147),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_135),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.C(n_143),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_136),
.A2(n_143),
.B1(n_144),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_143),
.B(n_258),
.C(n_261),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_143),
.A2(n_144),
.B1(n_258),
.B2(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_153),
.C(n_155),
.Y(n_169)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_169),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_162),
.B(n_167),
.C(n_169),
.Y(n_430)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.C(n_181),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_182),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_208),
.C(n_212),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_183),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_198),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_185),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_198),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_194),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_196),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_199),
.A2(n_202),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_202),
.A2(n_255),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_202),
.B(n_330),
.C(n_336),
.Y(n_363)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_203),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_212),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_386),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_274),
.C(n_279),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_266),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_SL g389 ( 
.A(n_220),
.B(n_266),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_250),
.C(n_264),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_221),
.B(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_235),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_236),
.C(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_223),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_224),
.B(n_227),
.Y(n_320)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_224),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_224),
.A2(n_339),
.B1(n_340),
.B2(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_248),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_251),
.B(n_264),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.C(n_262),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_252),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_257),
.B(n_263),
.Y(n_370)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_269),
.C(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_275),
.Y(n_388)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_276),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_381),
.B(n_385),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_366),
.B(n_380),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_324),
.B(n_365),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_311),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_283),
.B(n_311),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_298),
.C(n_305),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_285),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_289),
.C(n_293),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_298),
.A2(n_299),
.B1(n_305),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_300),
.B(n_302),
.Y(n_337)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

AO22x1_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_308),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_352),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_317),
.C(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_320),
.C(n_321),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_359),
.B(n_364),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_341),
.B(n_358),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_338),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_338),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_336),
.B2(n_337),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_340),
.Y(n_350)
);

AOI21x1_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_351),
.B(n_357),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_349),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_349),
.Y(n_357)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_363),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_378),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_378),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_371),
.B2(n_372),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_373),
.C(n_377),
.Y(n_382)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_382),
.B(n_383),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.C(n_389),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_432),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_396),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_423),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_411),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_407),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_418),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_431),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_427),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);


endmodule