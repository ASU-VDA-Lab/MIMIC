module fake_jpeg_12812_n_45 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_2),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_25),
.Y(n_33)
);

NOR4xp25_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_26),
.C(n_22),
.D(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_17),
.B1(n_5),
.B2(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_37),
.B(n_30),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_10),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_3),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.C(n_38),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_31),
.B(n_8),
.C(n_12),
.D(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_11),
.Y(n_45)
);


endmodule