module fake_jpeg_27750_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_27),
.C(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_41),
.B1(n_16),
.B2(n_17),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_28),
.B1(n_31),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_41),
.B1(n_58),
.B2(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_28),
.B1(n_31),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_21),
.B1(n_23),
.B2(n_16),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_69),
.B1(n_32),
.B2(n_44),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_65),
.B1(n_48),
.B2(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_38),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_83),
.B1(n_89),
.B2(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_37),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_54),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_40),
.CON(n_93),
.SN(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_33),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_37),
.B1(n_42),
.B2(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_89),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_112),
.B1(n_55),
.B2(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_97),
.Y(n_124)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_65),
.B1(n_44),
.B2(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_113),
.Y(n_140)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_48),
.B1(n_55),
.B2(n_62),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_90),
.B(n_51),
.C(n_78),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_81),
.B1(n_71),
.B2(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_42),
.B1(n_77),
.B2(n_55),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_99),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_136),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_80),
.B(n_79),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_131),
.B(n_24),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_87),
.B1(n_88),
.B2(n_84),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_70),
.B1(n_76),
.B2(n_91),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_76),
.B(n_60),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_34),
.C(n_90),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_141),
.C(n_34),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_95),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_143),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_63),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_131),
.B1(n_135),
.B2(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_153),
.B(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_163),
.B1(n_117),
.B2(n_136),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_168),
.B1(n_169),
.B2(n_134),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_96),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_90),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_115),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_127),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_77),
.B1(n_116),
.B2(n_42),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_128),
.B(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_51),
.B1(n_46),
.B2(n_34),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_180),
.B1(n_186),
.B2(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_118),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_191),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_163),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_117),
.C(n_125),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_184),
.C(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_166),
.B1(n_157),
.B2(n_130),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_185),
.B1(n_188),
.B2(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_133),
.B1(n_126),
.B2(n_134),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_133),
.C(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_133),
.B1(n_42),
.B2(n_106),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_22),
.B1(n_17),
.B2(n_18),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_25),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_146),
.A2(n_106),
.B1(n_24),
.B2(n_22),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_25),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_15),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_159),
.B1(n_170),
.B2(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_184),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_174),
.B1(n_148),
.B2(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_221),
.B1(n_14),
.B2(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_217),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_164),
.C(n_150),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_211),
.C(n_214),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_169),
.B1(n_168),
.B2(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_177),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_160),
.C(n_46),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_160),
.B1(n_24),
.B2(n_22),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_15),
.C(n_19),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_19),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_15),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_221)
);

AOI221xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_182),
.B1(n_175),
.B2(n_188),
.C(n_178),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_173),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_237),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

AO221x1_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_208),
.B1(n_206),
.B2(n_202),
.C(n_214),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_12),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_11),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_243),
.B(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_210),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_256),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_203),
.B1(n_205),
.B2(n_201),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_205),
.B(n_213),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_2),
.B(n_3),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_222),
.B1(n_241),
.B2(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_210),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_207),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_11),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_229),
.C(n_233),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_228),
.B1(n_222),
.B2(n_224),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_271),
.B1(n_249),
.B2(n_251),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.C(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_230),
.C(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_264),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_227),
.B(n_207),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_275),
.B(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_216),
.C(n_1),
.Y(n_267)
);

OAI21x1_ASAP7_75t_SL g270 ( 
.A1(n_254),
.A2(n_0),
.B(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_246),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_3),
.B(n_4),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_255),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_268),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_244),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_289),
.B(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_285),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_256),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_267),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_266),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_296),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_297),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_6),
.B(n_7),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_279),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_287),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_286),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_295),
.B(n_281),
.C(n_8),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_303),
.B(n_300),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_311),
.B(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_314),
.B1(n_306),
.B2(n_9),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_7),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_8),
.Y(n_318)
);


endmodule