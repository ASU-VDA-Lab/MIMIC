module fake_jpeg_1726_n_494 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_50),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_60),
.Y(n_96)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_91),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_66),
.B(n_84),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_47),
.B1(n_30),
.B2(n_34),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_72),
.B(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_0),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_88),
.Y(n_101)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_20),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_85),
.B(n_86),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_15),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_3),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_97),
.A2(n_149),
.B1(n_93),
.B2(n_36),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_110),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_114),
.A2(n_41),
.B1(n_46),
.B2(n_42),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_122),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_30),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_146),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_39),
.B1(n_37),
.B2(n_44),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_131),
.B1(n_136),
.B2(n_23),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_135),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_63),
.A2(n_39),
.B1(n_37),
.B2(n_44),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_48),
.B(n_51),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_71),
.A2(n_81),
.B1(n_90),
.B2(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_37),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_138),
.B(n_139),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_80),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_47),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_142),
.B(n_145),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_70),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_67),
.B(n_29),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_52),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_47),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_83),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_157),
.B(n_164),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_101),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_117),
.Y(n_165)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_127),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_169),
.B(n_172),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_107),
.A2(n_70),
.B(n_31),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_170),
.A2(n_177),
.B(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_55),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_173),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_174),
.B(n_180),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_29),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_209),
.C(n_124),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_23),
.B(n_18),
.Y(n_177)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_121),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_99),
.A2(n_23),
.B1(n_31),
.B2(n_38),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_182),
.A2(n_185),
.B1(n_189),
.B2(n_5),
.Y(n_253)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_99),
.A2(n_42),
.B1(n_18),
.B2(n_40),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_94),
.B(n_18),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_114),
.A2(n_78),
.B1(n_77),
.B2(n_41),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_194),
.B1(n_198),
.B2(n_118),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_104),
.A2(n_42),
.B1(n_31),
.B2(n_40),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_121),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_200),
.Y(n_213)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_100),
.A2(n_33),
.B(n_50),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_109),
.A2(n_57),
.B1(n_53),
.B2(n_49),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_105),
.A2(n_57),
.B1(n_53),
.B2(n_22),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_208),
.B1(n_210),
.B2(n_143),
.Y(n_223)
);

AOI22x1_ASAP7_75t_L g198 ( 
.A1(n_140),
.A2(n_143),
.B1(n_120),
.B2(n_113),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_137),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_105),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_104),
.B(n_3),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_125),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_210)
);

AO21x2_ASAP7_75t_L g295 ( 
.A1(n_212),
.A2(n_240),
.B(n_242),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_238),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_239),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_154),
.A2(n_125),
.B1(n_102),
.B2(n_140),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_254),
.B1(n_210),
.B2(n_208),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_227),
.B(n_206),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_100),
.C(n_94),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_228),
.B(n_258),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_181),
.A2(n_148),
.B1(n_120),
.B2(n_102),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_186),
.B1(n_156),
.B2(n_167),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_96),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_172),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_154),
.A2(n_98),
.B1(n_103),
.B2(n_148),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_212),
.B1(n_223),
.B2(n_198),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_162),
.A2(n_134),
.A3(n_109),
.B1(n_126),
.B2(n_115),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_188),
.A2(n_103),
.B1(n_98),
.B2(n_134),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_174),
.A2(n_126),
.B1(n_115),
.B2(n_137),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_112),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_243),
.B(n_244),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_161),
.B(n_4),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_253),
.A2(n_254),
.B1(n_211),
.B2(n_159),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_170),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_179),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_6),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_179),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_164),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_6),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_262),
.A2(n_263),
.B1(n_270),
.B2(n_272),
.Y(n_346)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_215),
.B(n_211),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_308),
.B(n_261),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_214),
.A2(n_219),
.B1(n_251),
.B2(n_236),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_278),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_206),
.B1(n_196),
.B2(n_173),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_193),
.B(n_177),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_273),
.A2(n_275),
.B(n_276),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_194),
.B1(n_198),
.B2(n_207),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_215),
.B(n_251),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_173),
.B(n_163),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_214),
.A2(n_201),
.B1(n_167),
.B2(n_168),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_277),
.A2(n_298),
.B1(n_302),
.B2(n_305),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_161),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_281),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_156),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_282),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_217),
.A2(n_184),
.A3(n_195),
.B1(n_199),
.B2(n_209),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_180),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_219),
.B(n_167),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_205),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_217),
.B(n_200),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_291),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_191),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_250),
.A2(n_203),
.B1(n_192),
.B2(n_169),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_220),
.B(n_157),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_224),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_228),
.B(n_203),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_165),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_242),
.A2(n_190),
.B1(n_165),
.B2(n_175),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_178),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_245),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_250),
.A2(n_183),
.B(n_7),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_268),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_321),
.C(n_322),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_SL g315 ( 
.A(n_269),
.B(n_296),
.C(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_334),
.C(n_297),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_316),
.Y(n_358)
);

AO21x2_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_239),
.B(n_226),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_319),
.A2(n_338),
.B(n_283),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_216),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_216),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_268),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_328),
.B(n_331),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_273),
.B(n_308),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_245),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_224),
.C(n_257),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_307),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_295),
.A2(n_257),
.B1(n_225),
.B2(n_230),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_337),
.B1(n_342),
.B2(n_345),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_295),
.A2(n_230),
.B1(n_225),
.B2(n_241),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_R g338 ( 
.A(n_290),
.B(n_241),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_295),
.A2(n_241),
.B1(n_249),
.B2(n_256),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_249),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_347),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_281),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_295),
.A2(n_218),
.B1(n_222),
.B2(n_237),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_291),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_363),
.B(n_371),
.Y(n_386)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_366),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_341),
.A2(n_288),
.B1(n_300),
.B2(n_270),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_372),
.B(n_374),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_271),
.C(n_301),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_364),
.C(n_369),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_295),
.B1(n_266),
.B2(n_288),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_287),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_275),
.B(n_294),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_324),
.B(n_303),
.C(n_276),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_326),
.A2(n_295),
.B1(n_266),
.B2(n_263),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_280),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_330),
.B(n_341),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_317),
.A2(n_282),
.B(n_272),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_298),
.B(n_285),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_284),
.C(n_237),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_342),
.C(n_314),
.Y(n_394)
);

A2O1A1O1Ixp25_ASAP7_75t_L g377 ( 
.A1(n_317),
.A2(n_262),
.B(n_293),
.C(n_265),
.D(n_229),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_380),
.B(n_336),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_299),
.Y(n_378)
);

AOI221xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_310),
.B1(n_346),
.B2(n_344),
.C(n_338),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_337),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_310),
.A2(n_293),
.B(n_265),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_385),
.B1(n_396),
.B2(n_381),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_356),
.A2(n_319),
.B1(n_332),
.B2(n_343),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_406),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_378),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_408),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_380),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_355),
.A2(n_319),
.B1(n_345),
.B2(n_332),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_319),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_407),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_333),
.C(n_323),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_401),
.C(n_409),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_340),
.C(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_318),
.Y(n_403)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_371),
.A2(n_313),
.B(n_339),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_327),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_363),
.A2(n_339),
.B(n_327),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_329),
.C(n_292),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_372),
.C(n_367),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_420),
.C(n_428),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_413),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_404),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_415),
.B(n_425),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_419),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_402),
.A2(n_358),
.B1(n_351),
.B2(n_381),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_421),
.B1(n_386),
.B2(n_400),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_349),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_374),
.C(n_351),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_396),
.A2(n_357),
.B1(n_377),
.B2(n_373),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_353),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_424),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_375),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_368),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_360),
.B1(n_350),
.B2(n_329),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_429),
.B1(n_388),
.B2(n_403),
.Y(n_433)
);

OA22x2_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_360),
.B1(n_292),
.B2(n_299),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_394),
.B(n_382),
.C(n_398),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_407),
.C(n_409),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_229),
.C(n_222),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_352),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g450 ( 
.A(n_430),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_385),
.B1(n_383),
.B2(n_393),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_434),
.A2(n_439),
.B1(n_444),
.B2(n_448),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_389),
.B1(n_400),
.B2(n_398),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_389),
.B1(n_393),
.B2(n_383),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_440),
.Y(n_453)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_429),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_438),
.B(n_441),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_431),
.A2(n_406),
.B1(n_391),
.B2(n_408),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_442),
.B(n_445),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_411),
.A2(n_386),
.B1(n_382),
.B2(n_352),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_420),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_410),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_417),
.A2(n_9),
.B(n_11),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_451),
.A2(n_427),
.B(n_424),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_457),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_410),
.C(n_425),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_434),
.A2(n_423),
.B1(n_430),
.B2(n_412),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_458),
.A2(n_13),
.B1(n_14),
.B2(n_453),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_446),
.B(n_440),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_440),
.B1(n_435),
.B2(n_448),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_440),
.B1(n_446),
.B2(n_451),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_428),
.C(n_416),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_11),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_416),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_463),
.B(n_464),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_457),
.B(n_450),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_469),
.B(n_471),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_473),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_452),
.C(n_455),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_9),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_475),
.B(n_454),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_13),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_474),
.Y(n_482)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_466),
.A2(n_462),
.B1(n_475),
.B2(n_471),
.C(n_460),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_478),
.B1(n_470),
.B2(n_465),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_469),
.A2(n_453),
.B(n_458),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_480),
.A2(n_481),
.B(n_13),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_467),
.A2(n_464),
.B(n_463),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_483),
.B(n_484),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_465),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_485),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_13),
.C(n_482),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_486),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_487),
.A2(n_484),
.B(n_486),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_489),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_492),
.B(n_491),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_488),
.Y(n_494)
);


endmodule