module fake_jpeg_3214_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_7),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_43),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_23),
.B1(n_18),
.B2(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_57),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_30),
.B1(n_40),
.B2(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_61),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_22),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_9),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_41),
.B1(n_25),
.B2(n_17),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_83),
.B1(n_69),
.B2(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_17),
.B(n_25),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_69),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_25),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_49),
.B1(n_62),
.B2(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_92),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_50),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_98),
.C(n_100),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_99),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_69),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_52),
.B1(n_46),
.B2(n_67),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_78),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_79),
.C(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_82),
.B(n_77),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_90),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_100),
.C(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_76),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_109),
.B(n_82),
.C(n_77),
.Y(n_111)
);

NOR4xp25_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_110),
.C(n_106),
.D(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_106),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_105),
.B(n_109),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_119),
.B(n_121),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_110),
.B(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_113),
.C(n_102),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_117),
.C(n_81),
.Y(n_126)
);

OAI31xp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_63),
.A3(n_28),
.B(n_84),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_114),
.B(n_87),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_63),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_62),
.B(n_65),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule