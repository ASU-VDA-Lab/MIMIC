module fake_jpeg_17975_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_30),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_64),
.Y(n_76)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_41),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_34),
.B1(n_24),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_60),
.B1(n_36),
.B2(n_40),
.Y(n_74)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_68),
.B1(n_26),
.B2(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_43),
.B(n_33),
.C(n_31),
.Y(n_69)
);

AOI211xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_83),
.B(n_93),
.C(n_76),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_43),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_91),
.C(n_54),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_85),
.B1(n_27),
.B2(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_84),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_44),
.B1(n_20),
.B2(n_21),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_102)
);

NOR2x1_ASAP7_75t_R g103 ( 
.A(n_80),
.B(n_19),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_33),
.A3(n_44),
.B1(n_21),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_30),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_32),
.C(n_17),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_66),
.B1(n_48),
.B2(n_50),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_99),
.B1(n_106),
.B2(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_49),
.B1(n_58),
.B2(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_105),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_0),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_113),
.B(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_67),
.B1(n_61),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_61),
.B1(n_56),
.B2(n_46),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_54),
.B(n_1),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_46),
.B1(n_21),
.B2(n_32),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_89),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_80),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_80),
.B1(n_91),
.B2(n_88),
.Y(n_131)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_127),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_121),
.C(n_132),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_73),
.B1(n_90),
.B2(n_70),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_95),
.B(n_90),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_73),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_109),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_99),
.B(n_116),
.C(n_97),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_124),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_79),
.B1(n_75),
.B2(n_82),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_120),
.B1(n_110),
.B2(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_81),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_70),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_131),
.C(n_149),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_159),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_99),
.B1(n_102),
.B2(n_111),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_155),
.A2(n_158),
.B1(n_160),
.B2(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_166),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_111),
.B1(n_117),
.B2(n_97),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_103),
.B1(n_75),
.B2(n_77),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_95),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_71),
.B1(n_77),
.B2(n_46),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_179),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_132),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_163),
.B(n_154),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_187),
.C(n_188),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_195),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_134),
.C(n_142),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_134),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_142),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.C(n_161),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_154),
.B1(n_152),
.B2(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_175),
.B1(n_122),
.B2(n_126),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_203),
.B(n_206),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_152),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_150),
.B(n_153),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_159),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_160),
.C(n_165),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_125),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_125),
.C(n_130),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_157),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_151),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_153),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_122),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_193),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_178),
.B1(n_200),
.B2(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_234),
.B1(n_215),
.B2(n_199),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_204),
.C(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_224),
.C(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_188),
.C(n_172),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_190),
.C(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_190),
.C(n_173),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_17),
.C(n_23),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_175),
.B(n_130),
.C(n_156),
.D(n_126),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_137),
.B(n_32),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_244),
.C(n_246),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_205),
.CI(n_216),
.CON(n_240),
.SN(n_240)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_9),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_235),
.B(n_198),
.C(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_245),
.B1(n_247),
.B2(n_230),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_9),
.B1(n_15),
.B2(n_3),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_17),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_234),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_23),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.C(n_9),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_227),
.C(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_257),
.B(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_259),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_256),
.Y(n_268)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_229),
.A3(n_231),
.B1(n_233),
.B2(n_232),
.C(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_262),
.B1(n_12),
.B2(n_4),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_246),
.C(n_249),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_8),
.B(n_4),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_272),
.Y(n_278)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_238),
.B(n_244),
.Y(n_265)
);

AOI31xp33_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_269),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_271),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_241),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_252),
.C(n_1),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_5),
.C(n_6),
.Y(n_275)
);

AOI31xp67_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_7),
.A3(n_8),
.B(n_10),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_8),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_15),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_271),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_285),
.B(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_276),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_15),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_275),
.CI(n_16),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_292),
.B(n_291),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_287),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_16),
.Y(n_295)
);


endmodule