module fake_jpeg_15241_n_123 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_17),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_22),
.B1(n_14),
.B2(n_34),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_57),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_24),
.B(n_13),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_13),
.A3(n_16),
.B1(n_15),
.B2(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_34),
.B1(n_26),
.B2(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_62),
.B1(n_58),
.B2(n_49),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_21),
.B1(n_25),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_65),
.B1(n_51),
.B2(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_50),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_74),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_88),
.B1(n_68),
.B2(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_45),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_88),
.C(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_97),
.C(n_70),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_96),
.B1(n_64),
.B2(n_78),
.C(n_75),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_63),
.B(n_75),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_81),
.B(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_102),
.B1(n_105),
.B2(n_97),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.C(n_104),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_44),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_27),
.B(n_32),
.C(n_28),
.D(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_15),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_23),
.B(n_46),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_94),
.C(n_93),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_23),
.C(n_28),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_57),
.B1(n_10),
.B2(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_8),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_110),
.B(n_9),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_0),
.Y(n_120)
);

NAND4xp25_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_46),
.C(n_1),
.D(n_2),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_116),
.B1(n_4),
.B2(n_3),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_3),
.Y(n_123)
);


endmodule