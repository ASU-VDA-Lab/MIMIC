module fake_ariane_2807_n_2148 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2148);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2148;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_60),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_126),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_28),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_69),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_56),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_100),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_31),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_34),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_111),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_88),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_110),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_162),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_130),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_78),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_71),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_128),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_71),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_202),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_149),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_96),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_83),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_187),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_143),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_6),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_142),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_112),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_207),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_163),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_118),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_72),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_132),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_92),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_97),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_214),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_57),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_82),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_22),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_32),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_131),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_116),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_178),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_105),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_180),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_108),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_10),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_98),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_114),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_146),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_17),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_10),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_22),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_79),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_134),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_34),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_56),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_127),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_63),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_52),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_217),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_195),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_137),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_99),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_53),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_125),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_12),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_120),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_51),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_66),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_213),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_70),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_72),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_33),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_117),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_29),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_47),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_91),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_67),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_8),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_26),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_159),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_170),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_157),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_138),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_7),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_155),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_156),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_145),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_37),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_216),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_172),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_194),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_135),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_218),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_103),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_208),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_57),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_67),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_2),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_21),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_150),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_198),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_190),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_52),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_12),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_165),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_53),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_167),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_37),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_8),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_203),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_31),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_48),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_41),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_61),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_129),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_19),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_40),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_1),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_101),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_154),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_66),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_36),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_148),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_13),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_173),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_42),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_136),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_89),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_54),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_133),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_123),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_29),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_65),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_32),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_61),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_139),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_54),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_188),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_43),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_35),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_48),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_59),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_169),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_161),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_75),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_46),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_160),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_141),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_25),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_209),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_25),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_39),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_5),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_49),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_55),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_94),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_204),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_181),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_21),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_39),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_17),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_93),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_192),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_24),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_85),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_182),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_14),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_58),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_44),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_60),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_76),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_23),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_64),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_229),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_239),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_241),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_235),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_279),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_394),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_295),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_328),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_313),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_313),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_246),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_313),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_313),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_228),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_252),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_347),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_386),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_221),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_224),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_331),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_412),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_331),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_227),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_331),
.Y(n_473)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_231),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_331),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_331),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_224),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_334),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_274),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_425),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_256),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_334),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_234),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_284),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_234),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_274),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_278),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_402),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_256),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_357),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_320),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_320),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_340),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_287),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_407),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_290),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_340),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_292),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_303),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_308),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_248),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_248),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_251),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_251),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_263),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_326),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_333),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_254),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_254),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_255),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_253),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_255),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_266),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_359),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_266),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_283),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_283),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_267),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_338),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_332),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_332),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_244),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_391),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_280),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_359),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_291),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_373),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_373),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_361),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_363),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_411),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_297),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_301),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_305),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_364),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_309),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_317),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_312),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_439),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_365),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_316),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_317),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_319),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_366),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_330),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_369),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_236),
.Y(n_555)
);

CKINVDCx14_ASAP7_75t_R g556 ( 
.A(n_393),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_337),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_393),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_393),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_341),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_342),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_366),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_351),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_433),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_470),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_457),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_481),
.B(n_325),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_489),
.B(n_222),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_457),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_220),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_230),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_480),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_458),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_446),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_449),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_449),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_460),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_448),
.Y(n_584)
);

AND3x2_ASAP7_75t_L g585 ( 
.A(n_463),
.B(n_379),
.C(n_353),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_451),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_451),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_442),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_321),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_464),
.B(n_226),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_452),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_452),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_492),
.B(n_321),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_453),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_486),
.A2(n_369),
.B1(n_375),
.B2(n_370),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_453),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_456),
.B(n_270),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_462),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_469),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_469),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_450),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_479),
.B(n_232),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_233),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_488),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_488),
.B(n_240),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_445),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_496),
.B(n_441),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_471),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_473),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_496),
.B(n_243),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_459),
.A2(n_440),
.B1(n_375),
.B2(n_378),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_476),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_506),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_519),
.B(n_530),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_558),
.B(n_270),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_506),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_507),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_477),
.B(n_249),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_507),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_508),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_467),
.B(n_348),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_508),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_447),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_490),
.A2(n_370),
.B1(n_382),
.B2(n_378),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_362),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_497),
.B(n_499),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_513),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_564),
.A2(n_440),
.B1(n_438),
.B2(n_409),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_487),
.B(n_250),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_514),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_516),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_519),
.B(n_264),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_530),
.B(n_268),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_515),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_515),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_517),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_454),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_455),
.Y(n_653)
);

CKINVDCx6p67_ASAP7_75t_R g654 ( 
.A(n_555),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_517),
.Y(n_655)
);

OA21x2_ASAP7_75t_L g656 ( 
.A1(n_518),
.A2(n_521),
.B(n_520),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_474),
.B(n_372),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_521),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_656),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_602),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_575),
.B(n_502),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_503),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_625),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_572),
.B(n_504),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_625),
.B(n_511),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_625),
.B(n_512),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_565),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_656),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_572),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_568),
.B(n_589),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_656),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_656),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_623),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_602),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_601),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_568),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_624),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_631),
.B(n_557),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_624),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_643),
.B(n_524),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_535),
.C(n_534),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_572),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_624),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_576),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_601),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_602),
.Y(n_688)
);

AND3x1_ASAP7_75t_L g689 ( 
.A(n_621),
.B(n_381),
.C(n_376),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_637),
.B(n_541),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_631),
.B(n_635),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_602),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_638),
.B(n_548),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_624),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_605),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_571),
.B(n_554),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_635),
.B(n_510),
.Y(n_698)
);

AO21x2_ASAP7_75t_L g699 ( 
.A1(n_566),
.A2(n_273),
.B(n_272),
.Y(n_699)
);

AND3x2_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_484),
.C(n_468),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_621),
.A2(n_382),
.B1(n_397),
.B2(n_392),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_658),
.B(n_466),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_566),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_658),
.B(n_563),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_574),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_623),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_642),
.A2(n_392),
.B1(n_401),
.B2(n_397),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_642),
.A2(n_529),
.B1(n_531),
.B2(n_523),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_574),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_589),
.B(n_562),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_578),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_584),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_589),
.B(n_270),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_590),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_588),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_578),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_579),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_606),
.A2(n_401),
.B1(n_409),
.B2(n_408),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_600),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_580),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_589),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_580),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_600),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_606),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_627),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_623),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_623),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_581),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_594),
.B(n_545),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_581),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_594),
.B(n_609),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_594),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_605),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_613),
.B(n_544),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_600),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_610),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_594),
.B(n_550),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_610),
.Y(n_740)
);

CKINVDCx6p67_ASAP7_75t_R g741 ( 
.A(n_654),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_614),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_612),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_609),
.B(n_552),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_582),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_613),
.A2(n_552),
.B1(n_553),
.B2(n_546),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_633),
.B(n_527),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_623),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_627),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_614),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_615),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_609),
.B(n_410),
.C(n_408),
.Y(n_752)
);

AO21x2_ASAP7_75t_L g753 ( 
.A1(n_582),
.A2(n_285),
.B(n_282),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_586),
.B(n_528),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_617),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_587),
.Y(n_758)
);

BUFx6f_ASAP7_75t_SL g759 ( 
.A(n_646),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_617),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_652),
.B(n_222),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_619),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_623),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_270),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_640),
.Y(n_765)
);

INVxp33_ASAP7_75t_SL g766 ( 
.A(n_653),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_592),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_592),
.B(n_270),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_600),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_593),
.B(n_522),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_653),
.B(n_223),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_640),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_593),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_596),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_600),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_619),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_613),
.A2(n_385),
.B1(n_389),
.B2(n_384),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_632),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_640),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_596),
.B(n_522),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_598),
.B(n_525),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_654),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_646),
.B(n_223),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_598),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_599),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_599),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_570),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_590),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_640),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_640),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_640),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_607),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_570),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_573),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_573),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_567),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_597),
.B(n_491),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_567),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_583),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_567),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_608),
.B(n_536),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_629),
.B(n_525),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_583),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_646),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_613),
.B(n_493),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_591),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_600),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_585),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_646),
.B(n_225),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_591),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_595),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_567),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_634),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_629),
.B(n_225),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_629),
.B(n_660),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_595),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_629),
.B(n_660),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_632),
.A2(n_335),
.B1(n_417),
.B2(n_410),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_660),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_660),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_664),
.A2(n_641),
.B(n_644),
.C(n_636),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_792),
.B(n_697),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_782),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_SL g825 ( 
.A(n_759),
.B(n_465),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_680),
.B(n_788),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_678),
.B(n_672),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_678),
.B(n_616),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_819),
.B(n_647),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_672),
.B(n_648),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_672),
.B(n_663),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_671),
.B(n_237),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_759),
.B(n_559),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_712),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_680),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_756),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_712),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_788),
.B(n_498),
.Y(n_838)
);

HB1xp67_ASAP7_75t_SL g839 ( 
.A(n_669),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_671),
.B(n_237),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_667),
.B(n_636),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_703),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_668),
.B(n_641),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_773),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_714),
.B(n_494),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_773),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_671),
.B(n_238),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_725),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_644),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_684),
.B(n_820),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_672),
.B(n_649),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_672),
.B(n_649),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_669),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_693),
.B(n_651),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_691),
.B(n_651),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_684),
.B(n_238),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_684),
.B(n_820),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_SL g858 ( 
.A(n_759),
.B(n_417),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_725),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_728),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_705),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_677),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_821),
.B(n_242),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_672),
.B(n_657),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_722),
.B(n_657),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_728),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_691),
.B(n_495),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_722),
.B(n_626),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_734),
.B(n_626),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_783),
.B(n_538),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_698),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_709),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_734),
.B(n_630),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_687),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_687),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_698),
.B(n_639),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_711),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_695),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_694),
.B(n_639),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_683),
.B(n_645),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_755),
.B(n_539),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_694),
.B(n_645),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_696),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_711),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_801),
.B(n_650),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_736),
.B(n_540),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_736),
.B(n_650),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_805),
.B(n_809),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_716),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_655),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_675),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_670),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_661),
.A2(n_659),
.B1(n_655),
.B2(n_547),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_735),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_686),
.B(n_549),
.Y(n_895)
);

OAI221xp5_ASAP7_75t_L g896 ( 
.A1(n_777),
.A2(n_428),
.B1(n_390),
.B2(n_400),
.C(n_405),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_695),
.B(n_245),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_704),
.B(n_715),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_715),
.B(n_549),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_738),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_666),
.B(n_659),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_739),
.B(n_420),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_784),
.B(n_245),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_784),
.B(n_675),
.Y(n_904)
);

OAI22xp33_ASAP7_75t_L g905 ( 
.A1(n_813),
.A2(n_432),
.B1(n_414),
.B2(n_436),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_716),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_666),
.B(n_526),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_670),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_665),
.B(n_420),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_675),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_679),
.B(n_532),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_681),
.B(n_532),
.Y(n_912)
);

INVxp33_ASAP7_75t_L g913 ( 
.A(n_747),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_743),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_805),
.B(n_551),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_685),
.B(n_533),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_675),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_717),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_717),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_740),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_718),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_675),
.B(n_247),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_706),
.B(n_247),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_702),
.B(n_422),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_804),
.B(n_422),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_743),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_706),
.B(n_257),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_726),
.B(n_533),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_740),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_710),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_706),
.B(n_257),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_718),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_742),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_749),
.A2(n_778),
.B(n_750),
.C(n_751),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_706),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_661),
.A2(n_537),
.B1(n_542),
.B2(n_543),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_L g937 ( 
.A(n_721),
.B(n_600),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_733),
.B(n_542),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_814),
.B(n_423),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_721),
.A2(n_730),
.B1(n_732),
.B2(n_723),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_815),
.B(n_543),
.Y(n_941)
);

INVx6_ASAP7_75t_L g942 ( 
.A(n_808),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_706),
.B(n_727),
.Y(n_943)
);

INVxp33_ASAP7_75t_L g944 ( 
.A(n_719),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_665),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_817),
.B(n_744),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_690),
.B(n_429),
.C(n_421),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_746),
.B(n_547),
.Y(n_948)
);

INVx8_ASAP7_75t_L g949 ( 
.A(n_665),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_732),
.A2(n_423),
.B1(n_427),
.B2(n_435),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_750),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_751),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_752),
.B(n_427),
.Y(n_953)
);

AO22x2_ASAP7_75t_L g954 ( 
.A1(n_707),
.A2(n_560),
.B1(n_551),
.B2(n_561),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_745),
.B(n_258),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_745),
.B(n_258),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_758),
.A2(n_437),
.B(n_560),
.C(n_561),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_758),
.B(n_767),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_767),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_727),
.B(n_259),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_774),
.Y(n_961)
);

NAND2xp33_ASAP7_75t_L g962 ( 
.A(n_774),
.B(n_259),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_754),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_701),
.B(n_478),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_797),
.B(n_478),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_785),
.B(n_260),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_727),
.B(n_260),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_741),
.B(n_482),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_700),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_766),
.Y(n_970)
);

AND2x6_ASAP7_75t_SL g971 ( 
.A(n_797),
.B(n_482),
.Y(n_971)
);

INVx8_ASAP7_75t_L g972 ( 
.A(n_713),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_785),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_754),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_808),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_786),
.B(n_261),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_761),
.B(n_435),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_786),
.B(n_261),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_808),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_771),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_802),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_727),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_854),
.B(n_766),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_918),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_942),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_823),
.B(n_708),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_854),
.A2(n_676),
.B(n_688),
.C(n_662),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_853),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_871),
.B(n_797),
.Y(n_989)
);

NOR2x1p5_ASAP7_75t_L g990 ( 
.A(n_824),
.B(n_741),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_862),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_945),
.B(n_797),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_885),
.B(n_670),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_SL g994 ( 
.A(n_944),
.B(n_813),
.Y(n_994)
);

AND2x6_ASAP7_75t_SL g995 ( 
.A(n_895),
.B(n_689),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_891),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_918),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_878),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_831),
.B(n_727),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_874),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_860),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_875),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_878),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_883),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_930),
.B(n_748),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_837),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_945),
.B(n_720),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_839),
.B(n_673),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_842),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_965),
.A2(n_829),
.B1(n_888),
.B2(n_881),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_934),
.A2(n_780),
.B(n_781),
.C(n_770),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_826),
.B(n_818),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_829),
.B(n_835),
.Y(n_1013)
);

NOR2x2_ASAP7_75t_L g1014 ( 
.A(n_870),
.B(n_662),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_SL g1015 ( 
.A(n_970),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_891),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_942),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_838),
.B(n_845),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_855),
.B(n_673),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_855),
.B(n_876),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_834),
.A2(n_848),
.B1(n_866),
.B2(n_859),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_925),
.B(n_729),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_954),
.A2(n_753),
.B1(n_699),
.B2(n_674),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_888),
.B(n_915),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_977),
.A2(n_438),
.B(n_757),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_899),
.B(n_827),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_851),
.B(n_729),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_828),
.B(n_713),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_891),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_841),
.A2(n_688),
.B(n_692),
.C(n_676),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_894),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_900),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_942),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_968),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_954),
.A2(n_753),
.B1(n_699),
.B2(n_674),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_886),
.B(n_713),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_965),
.A2(n_713),
.B1(n_776),
.B2(n_762),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_920),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_929),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_933),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_886),
.B(n_713),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_915),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_972),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_951),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_914),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_926),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_861),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_980),
.B(n_748),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_981),
.B(n_748),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_849),
.B(n_757),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_952),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_954),
.A2(n_753),
.B1(n_699),
.B2(n_811),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_822),
.A2(n_776),
.B(n_762),
.C(n_760),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_841),
.A2(n_692),
.B(n_760),
.C(n_791),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_872),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_963),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_975),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_892),
.A2(n_790),
.B(n_789),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_887),
.B(n_793),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_979),
.B(n_720),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_971),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_867),
.B(n_794),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_974),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_911),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_852),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_898),
.B(n_763),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_972),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_891),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_949),
.B(n_720),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_946),
.A2(n_790),
.B(n_789),
.Y(n_1070)
);

AND3x2_ASAP7_75t_SL g1071 ( 
.A(n_825),
.B(n_795),
.C(n_787),
.Y(n_1071)
);

AND2x6_ASAP7_75t_SL g1072 ( 
.A(n_977),
.B(n_483),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_972),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_908),
.A2(n_791),
.B(n_765),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_879),
.B(n_794),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_905),
.A2(n_896),
.B1(n_964),
.B2(n_884),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_879),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_872),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_882),
.B(n_806),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_949),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_949),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_884),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_909),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_961),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_953),
.B(n_765),
.C(n_763),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_969),
.B(n_737),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_882),
.B(n_806),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_912),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_864),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_870),
.Y(n_1091)
);

INVx5_ASAP7_75t_L g1092 ( 
.A(n_917),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_916),
.Y(n_1093)
);

AND2x6_ASAP7_75t_L g1094 ( 
.A(n_830),
.B(n_729),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_917),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_890),
.B(n_811),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_836),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_843),
.A2(n_765),
.B(n_772),
.C(n_779),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_844),
.B(n_772),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_961),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_846),
.Y(n_1101)
);

OR2x2_ASAP7_75t_SL g1102 ( 
.A(n_833),
.B(n_905),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_890),
.B(n_843),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_902),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_902),
.B(n_483),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_917),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_832),
.B(n_265),
.C(n_262),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_953),
.B(n_787),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_973),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_924),
.B(n_485),
.Y(n_1110)
);

BUFx4f_ASAP7_75t_L g1111 ( 
.A(n_917),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_924),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_865),
.B(n_948),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_913),
.B(n_485),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_897),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_939),
.A2(n_779),
.B(n_772),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_903),
.B(n_779),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_877),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_SL g1119 ( 
.A1(n_939),
.A2(n_398),
.B1(n_277),
.B2(n_276),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_889),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_982),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_906),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_910),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_903),
.B(n_795),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_936),
.B(n_816),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_935),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_919),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_863),
.B(n_798),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_893),
.A2(n_810),
.B1(n_803),
.B2(n_799),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_936),
.B(n_799),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_SL g1131 ( 
.A(n_832),
.B(n_265),
.C(n_262),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_921),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_938),
.B(n_803),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_935),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_934),
.B(n_810),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_R g1136 ( 
.A(n_858),
.B(n_937),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_907),
.B(n_798),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_932),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_868),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_893),
.A2(n_769),
.B1(n_807),
.B2(n_737),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_897),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_959),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_928),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_982),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_869),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_950),
.B(n_501),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_982),
.Y(n_1148)
);

INVx4_ASAP7_75t_L g1149 ( 
.A(n_982),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_880),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_822),
.A2(n_800),
.B1(n_798),
.B2(n_807),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_SL g1152 ( 
.A(n_840),
.B(n_271),
.C(n_269),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_957),
.B(n_769),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_955),
.B(n_501),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_873),
.Y(n_1155)
);

AND3x4_ASAP7_75t_L g1156 ( 
.A(n_988),
.B(n_947),
.C(n_618),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1020),
.A2(n_941),
.B1(n_940),
.B2(n_901),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1001),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1019),
.A2(n_904),
.B(n_943),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_983),
.B(n_956),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1067),
.B(n_724),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_1081),
.B(n_856),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1013),
.B(n_966),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1008),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_1053),
.A2(n_904),
.B(n_943),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1070),
.A2(n_857),
.B(n_850),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1033),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1104),
.B(n_856),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_991),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1081),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1045),
.B(n_962),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_989),
.A2(n_978),
.B1(n_976),
.B2(n_374),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_993),
.A2(n_857),
.B(n_850),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1103),
.A2(n_840),
.B1(n_847),
.B2(n_931),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_999),
.A2(n_923),
.B(n_922),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1009),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_994),
.A2(n_967),
.B1(n_960),
.B2(n_931),
.Y(n_1177)
);

CKINVDCx16_ASAP7_75t_R g1178 ( 
.A(n_1015),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_989),
.A2(n_275),
.B1(n_271),
.B2(n_269),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_1007),
.B(n_796),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1015),
.B(n_275),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_L g1182 ( 
.A(n_990),
.B(n_922),
.Y(n_1182)
);

BUFx4f_ASAP7_75t_L g1183 ( 
.A(n_992),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1013),
.B(n_847),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1010),
.B(n_923),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1104),
.B(n_927),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1001),
.B(n_927),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1077),
.B(n_796),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1112),
.B(n_796),
.Y(n_1189)
);

BUFx2_ASAP7_75t_SL g1190 ( 
.A(n_1081),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1081),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1006),
.B(n_796),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_327),
.B(n_367),
.C(n_380),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1018),
.B(n_505),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_1080),
.B(n_276),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1021),
.B(n_1072),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1034),
.B(n_1024),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1053),
.A2(n_620),
.B(n_603),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1047),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1024),
.B(n_812),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1111),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1000),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1002),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1067),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1055),
.Y(n_1205)
);

AND2x6_ASAP7_75t_L g1206 ( 
.A(n_1007),
.B(n_812),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1050),
.A2(n_300),
.B(n_304),
.C(n_293),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1077),
.B(n_812),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1046),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1069),
.B(n_1086),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1026),
.A2(n_356),
.B(n_354),
.C(n_349),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1078),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1073),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1004),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1066),
.A2(n_358),
.B(n_310),
.C(n_314),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_985),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1111),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1012),
.B(n_277),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1073),
.B(n_724),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1074),
.A2(n_775),
.B(n_724),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1082),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1084),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1073),
.B(n_315),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1058),
.A2(n_1079),
.B(n_1075),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1119),
.A2(n_1042),
.B1(n_992),
.B2(n_1091),
.Y(n_1225)
);

OAI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_1107),
.A2(n_318),
.B(n_315),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1076),
.B(n_505),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1042),
.Y(n_1228)
);

INVx5_ASAP7_75t_L g1229 ( 
.A(n_1069),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1144),
.B(n_603),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1102),
.A2(n_418),
.B1(n_430),
.B2(n_416),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1146),
.B(n_622),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1100),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_986),
.A2(n_426),
.B(n_344),
.C(n_324),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1061),
.B(n_431),
.C(n_318),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1076),
.A2(n_430),
.B1(n_371),
.B2(n_374),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1114),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1109),
.Y(n_1238)
);

OR2x6_ASAP7_75t_SL g1239 ( 
.A(n_1110),
.B(n_371),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_996),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_R g1241 ( 
.A(n_1017),
.B(n_377),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1073),
.B(n_377),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1069),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1155),
.B(n_724),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1014),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1060),
.B(n_383),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1105),
.B(n_567),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_987),
.A2(n_388),
.B(n_413),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1064),
.B(n_1088),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1066),
.A2(n_322),
.B(n_368),
.C(n_399),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_995),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1062),
.A2(n_404),
.B(n_406),
.C(n_434),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1060),
.B(n_1092),
.Y(n_1253)
);

CKINVDCx8_ASAP7_75t_R g1254 ( 
.A(n_1083),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_996),
.Y(n_1255)
);

CKINVDCx8_ASAP7_75t_R g1256 ( 
.A(n_1092),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1093),
.B(n_775),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1154),
.B(n_567),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1087),
.A2(n_775),
.B(n_345),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1120),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1092),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_996),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_R g1263 ( 
.A(n_1057),
.B(n_383),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_L g1264 ( 
.A(n_1150),
.B(n_387),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1059),
.A2(n_343),
.B(n_286),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1113),
.B(n_577),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1115),
.B(n_387),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1092),
.B(n_395),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1031),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1043),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_996),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1118),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1115),
.A2(n_395),
.B(n_396),
.C(n_398),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1054),
.A2(n_336),
.B(n_288),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1143),
.B(n_577),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1095),
.B(n_396),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1095),
.B(n_415),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1030),
.A2(n_339),
.B(n_289),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1133),
.A2(n_346),
.B(n_294),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1135),
.A2(n_350),
.B(n_296),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1098),
.A2(n_352),
.B(n_298),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1097),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1137),
.A2(n_355),
.B(n_299),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1101),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1097),
.B(n_577),
.Y(n_1285)
);

CKINVDCx14_ASAP7_75t_R g1286 ( 
.A(n_1136),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1122),
.Y(n_1287)
);

NOR3xp33_ASAP7_75t_SL g1288 ( 
.A(n_1032),
.B(n_431),
.C(n_418),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1011),
.A2(n_1151),
.B(n_1096),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1095),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1036),
.A2(n_1041),
.B1(n_1141),
.B2(n_1048),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1095),
.B(n_577),
.Y(n_1292)
);

NOR2x1_ASAP7_75t_L g1293 ( 
.A(n_1126),
.B(n_577),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_SL g1294 ( 
.A(n_1145),
.B(n_415),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1086),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1136),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1117),
.A2(n_1128),
.B(n_1011),
.C(n_1005),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1038),
.A2(n_416),
.B1(n_604),
.B2(n_577),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1147),
.B(n_604),
.Y(n_1299)
);

NOR3xp33_ASAP7_75t_SL g1300 ( 
.A(n_1039),
.B(n_281),
.C(n_302),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1005),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_SL g1302 ( 
.A(n_1040),
.B(n_307),
.C(n_311),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1145),
.B(n_323),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1044),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1051),
.B(n_604),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1139),
.B(n_329),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1166),
.A2(n_1027),
.B(n_1052),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1289),
.A2(n_1224),
.B(n_1157),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1169),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1175),
.A2(n_1108),
.B(n_1022),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1297),
.A2(n_1145),
.B(n_1029),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1237),
.B(n_1056),
.Y(n_1312)
);

NOR4xp25_ASAP7_75t_L g1313 ( 
.A(n_1282),
.B(n_1124),
.C(n_1023),
.D(n_1035),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1167),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1237),
.B(n_1063),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_L g1316 ( 
.A(n_1158),
.B(n_1150),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1174),
.A2(n_1029),
.B(n_1068),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1209),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1272),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1173),
.A2(n_1035),
.B(n_1023),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1236),
.A2(n_1107),
.B1(n_1131),
.B2(n_1152),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1287),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1174),
.A2(n_1106),
.B(n_1121),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_1181),
.Y(n_1324)
);

OAI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1168),
.A2(n_1131),
.B(n_1152),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1178),
.B(n_1139),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1249),
.B(n_1127),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1228),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1207),
.A2(n_1128),
.B(n_1049),
.C(n_1037),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1202),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1203),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1249),
.B(n_1132),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1214),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_SL g1334 ( 
.A(n_1196),
.B(n_1149),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1210),
.B(n_1164),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1163),
.B(n_1138),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1194),
.B(n_1142),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1195),
.Y(n_1338)
);

AOI31xp67_ASAP7_75t_L g1339 ( 
.A1(n_1266),
.A2(n_1184),
.A3(n_1148),
.B(n_1188),
.Y(n_1339)
);

CKINVDCx14_ASAP7_75t_R g1340 ( 
.A(n_1263),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1160),
.A2(n_1085),
.B(n_1116),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1256),
.Y(n_1342)
);

BUFx2_ASAP7_75t_R g1343 ( 
.A(n_1239),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1251),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1198),
.A2(n_1129),
.B(n_1125),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1201),
.Y(n_1346)
);

AO32x2_ASAP7_75t_L g1347 ( 
.A1(n_1231),
.A2(n_1071),
.A3(n_1149),
.B1(n_1085),
.B2(n_1065),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1301),
.B(n_1065),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1193),
.A2(n_1185),
.A3(n_1280),
.B(n_1298),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1156),
.A2(n_1049),
.B1(n_1089),
.B2(n_1153),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1252),
.A2(n_1099),
.B1(n_984),
.B2(n_997),
.C(n_1028),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1284),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1186),
.A2(n_1130),
.B1(n_1153),
.B2(n_1099),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_1153),
.B1(n_1089),
.B2(n_1140),
.Y(n_1354)
);

BUFx4_ASAP7_75t_SL g1355 ( 
.A(n_1216),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1188),
.A2(n_1068),
.B(n_1029),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1197),
.B(n_1296),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1248),
.A2(n_1094),
.B(n_998),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1306),
.B(n_1003),
.Y(n_1359)
);

AOI221xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1226),
.A2(n_1134),
.B1(n_1090),
.B2(n_1123),
.C(n_1106),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1165),
.A2(n_1248),
.B(n_1220),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1208),
.A2(n_1121),
.B(n_1016),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1269),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1208),
.A2(n_1106),
.B(n_1016),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1298),
.A2(n_1071),
.A3(n_1094),
.B(n_1150),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1165),
.A2(n_1090),
.B(n_1134),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1259),
.A2(n_1121),
.B(n_1016),
.Y(n_1367)
);

OA22x2_ASAP7_75t_L g1368 ( 
.A1(n_1225),
.A2(n_1123),
.B1(n_1043),
.B2(n_360),
.Y(n_1368)
);

AND3x1_ASAP7_75t_L g1369 ( 
.A(n_1235),
.B(n_0),
.C(n_3),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1286),
.B(n_1150),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1183),
.B(n_4),
.Y(n_1371)
);

NAND3x1_ASAP7_75t_L g1372 ( 
.A(n_1182),
.B(n_7),
.C(n_9),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1210),
.B(n_1068),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1267),
.B(n_1068),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1229),
.B(n_1243),
.Y(n_1375)
);

O2A1O1Ixp5_ASAP7_75t_SL g1376 ( 
.A1(n_1218),
.A2(n_604),
.B(n_764),
.C(n_768),
.Y(n_1376)
);

AOI31xp67_ASAP7_75t_L g1377 ( 
.A1(n_1291),
.A2(n_768),
.A3(n_764),
.B(n_604),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1179),
.A2(n_9),
.B(n_11),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1275),
.A2(n_768),
.B(n_764),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1303),
.A2(n_11),
.B(n_15),
.C(n_16),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1183),
.B(n_15),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1305),
.A2(n_306),
.B(n_84),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1234),
.A2(n_306),
.B(n_19),
.C(n_20),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1305),
.A2(n_86),
.B(n_219),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1230),
.A2(n_77),
.B(n_206),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1230),
.A2(n_151),
.B(n_193),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1192),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1254),
.B(n_18),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1215),
.A2(n_18),
.B(n_20),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1189),
.A2(n_306),
.B(n_191),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1250),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1391)
);

OAI22x1_ASAP7_75t_L g1392 ( 
.A1(n_1245),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1176),
.A2(n_90),
.A3(n_177),
.B(n_176),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1304),
.B(n_35),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1161),
.A2(n_87),
.B(n_174),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1245),
.B(n_36),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1293),
.A2(n_1232),
.B(n_1292),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1232),
.A2(n_189),
.B(n_166),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1261),
.A2(n_38),
.B(n_41),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1290),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1247),
.A2(n_38),
.B(n_44),
.Y(n_1401)
);

AO22x2_ASAP7_75t_L g1402 ( 
.A1(n_1295),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1260),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1240),
.A2(n_104),
.B(n_152),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1190),
.B(n_50),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1201),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1180),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1229),
.B(n_147),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1281),
.A2(n_1278),
.B(n_1274),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1171),
.B(n_50),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_SL g1411 ( 
.A1(n_1246),
.A2(n_51),
.B(n_55),
.C(n_58),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1187),
.B(n_59),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1227),
.A2(n_1244),
.B(n_1257),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1199),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1200),
.B(n_62),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1205),
.A2(n_124),
.A3(n_122),
.B(n_115),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1212),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1300),
.A2(n_1302),
.B(n_1288),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1253),
.A2(n_62),
.B(n_63),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1241),
.B(n_64),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1172),
.B(n_65),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1221),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1257),
.A2(n_68),
.B(n_69),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1201),
.Y(n_1424)
);

BUFx4_ASAP7_75t_SL g1425 ( 
.A(n_1285),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1217),
.B(n_1273),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1299),
.B(n_68),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1217),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1211),
.A2(n_1162),
.B(n_1265),
.C(n_1279),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1295),
.B(n_70),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1222),
.B(n_73),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1283),
.A2(n_73),
.B(n_1258),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1244),
.A2(n_1270),
.B(n_1277),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1233),
.B(n_1238),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1255),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1264),
.B(n_1276),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1437)
);

AOI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_1223),
.B(n_1242),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1170),
.B(n_1191),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1170),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1170),
.A2(n_1191),
.B(n_1271),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1262),
.A2(n_1243),
.B(n_1229),
.Y(n_1442)
);

NAND2x1_ASAP7_75t_L g1443 ( 
.A(n_1204),
.B(n_1213),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1180),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1191),
.B(n_1180),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1204),
.B(n_1213),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1219),
.A2(n_1180),
.B(n_1206),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1206),
.B(n_1020),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1166),
.A2(n_1289),
.B(n_1159),
.Y(n_1449)
);

INVxp67_ASAP7_75t_SL g1450 ( 
.A(n_1158),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1168),
.A2(n_854),
.B(n_1104),
.C(n_823),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1237),
.B(n_983),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1239),
.A2(n_983),
.B1(n_944),
.B2(n_1104),
.Y(n_1453)
);

OAI21xp33_ASAP7_75t_L g1454 ( 
.A1(n_1168),
.A2(n_983),
.B(n_664),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1166),
.A2(n_1289),
.B(n_1159),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1167),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1282),
.A2(n_1174),
.B1(n_983),
.B2(n_1236),
.C(n_1289),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1169),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1166),
.A2(n_1289),
.B(n_1159),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1169),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1237),
.B(n_983),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1358),
.A2(n_1409),
.B(n_1320),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1454),
.A2(n_1451),
.B(n_1389),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1454),
.A2(n_1389),
.B(n_1457),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1307),
.Y(n_1466)
);

AO222x2_ASAP7_75t_L g1467 ( 
.A1(n_1420),
.A2(n_1343),
.B1(n_1453),
.B2(n_1396),
.C1(n_1392),
.C2(n_1412),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1335),
.B(n_1447),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1348),
.B(n_1336),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1378),
.A2(n_1325),
.B1(n_1457),
.B2(n_1321),
.C(n_1421),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1450),
.B(n_1371),
.Y(n_1471)
);

INVx8_ASAP7_75t_L g1472 ( 
.A(n_1407),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1312),
.B(n_1315),
.Y(n_1473)
);

OAI211xp5_ASAP7_75t_L g1474 ( 
.A1(n_1378),
.A2(n_1325),
.B(n_1401),
.C(n_1391),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1381),
.B(n_1402),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1448),
.A2(n_1329),
.B(n_1383),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1327),
.B(n_1332),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1402),
.A2(n_1321),
.B1(n_1401),
.B2(n_1368),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1361),
.A2(n_1366),
.B(n_1310),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1369),
.B(n_1419),
.C(n_1432),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1344),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1317),
.A2(n_1323),
.B(n_1345),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1428),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1357),
.B(n_1334),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1367),
.A2(n_1409),
.B(n_1311),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1309),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1385),
.A2(n_1386),
.B(n_1398),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1407),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1355),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1407),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1326),
.B(n_1388),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1335),
.B(n_1408),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1328),
.B(n_1330),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1405),
.A2(n_1334),
.B1(n_1350),
.B2(n_1354),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1331),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1333),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1413),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1337),
.B(n_1387),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1384),
.A2(n_1397),
.B(n_1364),
.Y(n_1500)
);

CKINVDCx14_ASAP7_75t_R g1501 ( 
.A(n_1340),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1427),
.B(n_1318),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1352),
.B(n_1363),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1405),
.B(n_1369),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_SL g1505 ( 
.A1(n_1448),
.A2(n_1429),
.B(n_1432),
.C(n_1374),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1350),
.A2(n_1415),
.B1(n_1405),
.B2(n_1359),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1353),
.A2(n_1358),
.B(n_1362),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1353),
.A2(n_1341),
.B(n_1360),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1458),
.B(n_1460),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1342),
.B(n_1319),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1408),
.B(n_1313),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1341),
.A2(n_1423),
.B(n_1354),
.C(n_1426),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1360),
.B(n_1313),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1433),
.A2(n_1411),
.B(n_1356),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1373),
.Y(n_1515)
);

BUFx4_ASAP7_75t_SL g1516 ( 
.A(n_1338),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1322),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1424),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1342),
.B(n_1370),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1382),
.A2(n_1390),
.B(n_1413),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1406),
.B(n_1314),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_1324),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1403),
.A2(n_1417),
.B1(n_1422),
.B2(n_1414),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1394),
.A2(n_1410),
.B1(n_1436),
.B2(n_1372),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1335),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1430),
.A2(n_1437),
.B1(n_1444),
.B2(n_1431),
.Y(n_1526)
);

OAI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1380),
.A2(n_1431),
.B(n_1438),
.C(n_1351),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1440),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1376),
.A2(n_1404),
.B(n_1395),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1440),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1434),
.Y(n_1532)
);

AO21x1_ASAP7_75t_L g1533 ( 
.A1(n_1445),
.A2(n_1439),
.B(n_1435),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1379),
.A2(n_1443),
.B(n_1442),
.Y(n_1534)
);

NOR2xp67_ASAP7_75t_L g1535 ( 
.A(n_1456),
.B(n_1316),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1393),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1446),
.B(n_1400),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1347),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1347),
.A2(n_1349),
.B(n_1365),
.C(n_1400),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1440),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1346),
.B(n_1441),
.Y(n_1541)
);

OR2x4_ASAP7_75t_L g1542 ( 
.A(n_1346),
.B(n_1418),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1379),
.A2(n_1399),
.B(n_1377),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1393),
.A2(n_1416),
.B(n_1349),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1346),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1425),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1365),
.A2(n_1349),
.B1(n_1393),
.B2(n_1416),
.Y(n_1547)
);

AOI21xp33_ASAP7_75t_L g1548 ( 
.A1(n_1365),
.A2(n_1207),
.B(n_1234),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1416),
.A2(n_1236),
.B1(n_954),
.B2(n_1454),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1318),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1428),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1407),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1309),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1309),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1454),
.A2(n_1236),
.B1(n_954),
.B2(n_1402),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1307),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1412),
.B(n_1196),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1309),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1407),
.Y(n_1561)
);

NAND2x1p5_ASAP7_75t_L g1562 ( 
.A(n_1407),
.B(n_1229),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1454),
.A2(n_854),
.B(n_1451),
.C(n_1378),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_SL g1564 ( 
.A1(n_1451),
.A2(n_1297),
.B(n_1454),
.C(n_1448),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1224),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1454),
.A2(n_1236),
.B1(n_954),
.B2(n_1402),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1407),
.Y(n_1569)
);

INVx11_ASAP7_75t_L g1570 ( 
.A(n_1355),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1355),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1318),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1309),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1224),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1454),
.A2(n_983),
.B1(n_1451),
.B2(n_1104),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1576)
);

BUFx2_ASAP7_75t_SL g1577 ( 
.A(n_1428),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1339),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1454),
.B(n_983),
.C(n_664),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1448),
.B(n_1454),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1358),
.A2(n_1409),
.B(n_1320),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1454),
.B(n_664),
.C(n_628),
.D(n_643),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1585)
);

CKINVDCx11_ASAP7_75t_R g1586 ( 
.A(n_1338),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1309),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1407),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1308),
.A2(n_1455),
.B(n_1449),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1309),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1308),
.A2(n_1455),
.B(n_1449),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1224),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1318),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1412),
.B(n_1196),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1309),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1402),
.A2(n_1236),
.B1(n_954),
.B2(n_646),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1307),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1454),
.A2(n_983),
.B1(n_1451),
.B2(n_1104),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1339),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1454),
.A2(n_983),
.B1(n_1451),
.B2(n_1104),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1454),
.A2(n_983),
.B(n_1451),
.C(n_1104),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1453),
.A2(n_905),
.B1(n_944),
.B2(n_689),
.C(n_1104),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1454),
.A2(n_983),
.B(n_664),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1454),
.A2(n_983),
.B1(n_1451),
.B2(n_1104),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1309),
.Y(n_1612)
);

BUFx8_ASAP7_75t_L g1613 ( 
.A(n_1318),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1454),
.A2(n_1236),
.B1(n_954),
.B2(n_1402),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1407),
.B(n_1229),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1454),
.A2(n_1236),
.B1(n_954),
.B2(n_1402),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1428),
.Y(n_1617)
);

CKINVDCx8_ASAP7_75t_R g1618 ( 
.A(n_1324),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1335),
.B(n_1210),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1454),
.A2(n_983),
.B(n_664),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1355),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1309),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1454),
.A2(n_983),
.B1(n_1451),
.B2(n_1104),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1224),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1455),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1454),
.A2(n_854),
.B(n_1451),
.C(n_1378),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1308),
.A2(n_1455),
.B(n_1449),
.Y(n_1630)
);

AOI221x1_ASAP7_75t_SL g1631 ( 
.A1(n_1584),
.A2(n_1580),
.B1(n_1605),
.B2(n_1610),
.C(n_1603),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1585),
.B(n_1625),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1563),
.A2(n_1629),
.B1(n_1470),
.B2(n_1621),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1494),
.B(n_1503),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1607),
.C(n_1463),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1558),
.B(n_1598),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1477),
.B(n_1465),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1609),
.A2(n_1600),
.B1(n_1616),
.B2(n_1614),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1568),
.B(n_1582),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1487),
.Y(n_1642)
);

CKINVDCx6p67_ASAP7_75t_R g1643 ( 
.A(n_1586),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1474),
.A2(n_1512),
.B(n_1478),
.C(n_1464),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1474),
.A2(n_1512),
.B(n_1478),
.C(n_1600),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1556),
.A2(n_1614),
.B1(n_1616),
.B2(n_1567),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1485),
.B(n_1492),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_SL g1648 ( 
.A1(n_1504),
.A2(n_1521),
.B(n_1466),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1466),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1572),
.B(n_1596),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1589),
.B(n_1608),
.Y(n_1652)
);

CKINVDCx6p67_ASAP7_75t_R g1653 ( 
.A(n_1586),
.Y(n_1653)
);

BUFx2_ASAP7_75t_R g1654 ( 
.A(n_1490),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1511),
.B(n_1550),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1501),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1657)
);

AOI21x1_ASAP7_75t_SL g1658 ( 
.A1(n_1557),
.A2(n_1602),
.B(n_1498),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1556),
.A2(n_1567),
.B1(n_1480),
.B2(n_1626),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1513),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1575),
.A2(n_1495),
.B1(n_1606),
.B2(n_1506),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1606),
.A2(n_1564),
.B(n_1505),
.C(n_1495),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1542),
.A2(n_1546),
.B1(n_1549),
.B2(n_1476),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1565),
.A2(n_1595),
.B(n_1574),
.Y(n_1665)
);

OAI22x1_ASAP7_75t_L g1666 ( 
.A1(n_1467),
.A2(n_1555),
.B1(n_1599),
.B2(n_1624),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1613),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1509),
.B(n_1473),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1493),
.A2(n_1524),
.B(n_1526),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1493),
.A2(n_1527),
.B(n_1569),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1554),
.B(n_1560),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_SL g1672 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1544),
.A2(n_1520),
.B(n_1486),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1573),
.B(n_1587),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1565),
.A2(n_1574),
.B(n_1595),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1527),
.A2(n_1569),
.B(n_1508),
.Y(n_1676)
);

AOI21x1_ASAP7_75t_SL g1677 ( 
.A1(n_1541),
.A2(n_1542),
.B(n_1510),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_SL g1678 ( 
.A(n_1619),
.B(n_1561),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1564),
.A2(n_1505),
.B(n_1513),
.C(n_1581),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1592),
.B(n_1612),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1532),
.B(n_1581),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1549),
.A2(n_1507),
.B(n_1548),
.C(n_1539),
.Y(n_1683)
);

AOI31xp33_ASAP7_75t_L g1684 ( 
.A1(n_1501),
.A2(n_1571),
.A3(n_1622),
.B(n_1467),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1528),
.B(n_1551),
.Y(n_1685)
);

OA22x2_ASAP7_75t_L g1686 ( 
.A1(n_1538),
.A2(n_1588),
.B1(n_1481),
.B2(n_1540),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1484),
.A2(n_1577),
.B1(n_1522),
.B2(n_1518),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1551),
.B(n_1617),
.Y(n_1688)
);

O2A1O1Ixp5_ASAP7_75t_L g1689 ( 
.A1(n_1627),
.A2(n_1507),
.B(n_1520),
.C(n_1530),
.Y(n_1689)
);

AND2x2_ASAP7_75t_SL g1690 ( 
.A(n_1489),
.B(n_1536),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1537),
.B(n_1517),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1613),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1472),
.B(n_1491),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_R g1695 ( 
.A(n_1482),
.B(n_1618),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1531),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1552),
.A2(n_1579),
.B(n_1559),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1515),
.B(n_1545),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1514),
.A2(n_1547),
.B1(n_1583),
.B2(n_1462),
.C(n_1523),
.Y(n_1699)
);

O2A1O1Ixp5_ASAP7_75t_L g1700 ( 
.A1(n_1578),
.A2(n_1604),
.B(n_1533),
.C(n_1553),
.Y(n_1700)
);

AOI21x1_ASAP7_75t_SL g1701 ( 
.A1(n_1516),
.A2(n_1488),
.B(n_1570),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1561),
.A2(n_1535),
.B1(n_1491),
.B2(n_1590),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1553),
.B(n_1590),
.Y(n_1703)
);

O2A1O1Ixp5_ASAP7_75t_L g1704 ( 
.A1(n_1578),
.A2(n_1604),
.B(n_1536),
.C(n_1543),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1491),
.A2(n_1615),
.B1(n_1562),
.B2(n_1489),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1516),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1472),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1489),
.B(n_1534),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1500),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1591),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1591),
.B(n_1630),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1483),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1593),
.A2(n_1630),
.B(n_1597),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1593),
.B(n_1479),
.Y(n_1714)
);

AOI21x1_ASAP7_75t_SL g1715 ( 
.A1(n_1566),
.A2(n_1601),
.B(n_1623),
.Y(n_1715)
);

AOI21x1_ASAP7_75t_SL g1716 ( 
.A1(n_1576),
.A2(n_1594),
.B(n_1611),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1620),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1628),
.B(n_1471),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1584),
.C(n_1621),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1565),
.A2(n_1595),
.B(n_1574),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1565),
.A2(n_1595),
.B(n_1574),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1584),
.C(n_1621),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1585),
.B(n_1625),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1629),
.B2(n_1470),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1726)
);

CKINVDCx11_ASAP7_75t_R g1727 ( 
.A(n_1618),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1584),
.C(n_1621),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1494),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1730)
);

AOI21x1_ASAP7_75t_SL g1731 ( 
.A1(n_1504),
.A2(n_983),
.B(n_1186),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1629),
.B2(n_1470),
.Y(n_1732)
);

AND2x6_ASAP7_75t_L g1733 ( 
.A(n_1489),
.B(n_1553),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1494),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1494),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1494),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1522),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1584),
.C(n_1621),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1565),
.A2(n_1595),
.B(n_1574),
.Y(n_1741)
);

INVxp33_ASAP7_75t_SL g1742 ( 
.A(n_1516),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1466),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1522),
.A2(n_1196),
.B1(n_1501),
.B2(n_1470),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1544),
.A2(n_1520),
.B(n_1486),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1512),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1512),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1629),
.B2(n_1470),
.Y(n_1751)
);

O2A1O1Ixp33_ASAP7_75t_L g1752 ( 
.A1(n_1563),
.A2(n_1629),
.B(n_1584),
.C(n_1621),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1629),
.B2(n_1470),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1466),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1629),
.B2(n_1470),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1758)
);

AOI21x1_ASAP7_75t_SL g1759 ( 
.A1(n_1504),
.A2(n_983),
.B(n_1186),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1613),
.Y(n_1760)
);

O2A1O1Ixp5_ASAP7_75t_L g1761 ( 
.A1(n_1463),
.A2(n_1464),
.B(n_1629),
.C(n_1563),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1466),
.Y(n_1762)
);

O2A1O1Ixp5_ASAP7_75t_L g1763 ( 
.A1(n_1463),
.A2(n_1464),
.B(n_1629),
.C(n_1563),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1544),
.A2(n_1520),
.B(n_1486),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1471),
.B(n_1502),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1708),
.B(n_1672),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1632),
.B(n_1724),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1714),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1637),
.A2(n_1645),
.B(n_1644),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1689),
.A2(n_1675),
.B(n_1665),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1642),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1649),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1746),
.B(n_1748),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1636),
.B(n_1729),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1660),
.B(n_1635),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1683),
.A2(n_1713),
.B(n_1675),
.Y(n_1777)
);

AOI21x1_ASAP7_75t_L g1778 ( 
.A1(n_1713),
.A2(n_1712),
.B(n_1725),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1734),
.B(n_1735),
.Y(n_1779)
);

OAI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1640),
.A2(n_1646),
.B1(n_1659),
.B2(n_1662),
.C1(n_1664),
.C2(n_1634),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1718),
.B(n_1711),
.Y(n_1781)
);

NOR2x1_ASAP7_75t_L g1782 ( 
.A(n_1669),
.B(n_1676),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1649),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1671),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1710),
.B(n_1689),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1674),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1665),
.B(n_1721),
.Y(n_1789)
);

BUFx12f_ASAP7_75t_L g1790 ( 
.A(n_1727),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1722),
.B(n_1741),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1681),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1754),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1733),
.Y(n_1794)
);

OAI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1761),
.A2(n_1763),
.B(n_1739),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1682),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1691),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1762),
.B(n_1673),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1704),
.A2(n_1700),
.B(n_1763),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1720),
.A2(n_1752),
.B(n_1739),
.C(n_1728),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1673),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1660),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1745),
.Y(n_1804)
);

AO21x2_ASAP7_75t_L g1805 ( 
.A1(n_1732),
.A2(n_1751),
.B(n_1753),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1690),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1745),
.Y(n_1807)
);

AO21x2_ASAP7_75t_L g1808 ( 
.A1(n_1757),
.A2(n_1663),
.B(n_1720),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1765),
.B(n_1657),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1699),
.A2(n_1717),
.B(n_1709),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

AO21x2_ASAP7_75t_L g1812 ( 
.A1(n_1663),
.A2(n_1728),
.B(n_1723),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1690),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_L g1814 ( 
.A(n_1733),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1686),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1686),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1730),
.B(n_1740),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1661),
.B(n_1633),
.Y(n_1818)
);

AO21x2_ASAP7_75t_L g1819 ( 
.A1(n_1723),
.A2(n_1752),
.B(n_1680),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1668),
.Y(n_1820)
);

OA21x2_ASAP7_75t_L g1821 ( 
.A1(n_1699),
.A2(n_1755),
.B(n_1756),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1680),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1697),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1697),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1719),
.B(n_1726),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1747),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1758),
.Y(n_1827)
);

AO21x2_ASAP7_75t_L g1828 ( 
.A1(n_1639),
.A2(n_1652),
.B(n_1641),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1737),
.B(n_1766),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1703),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1733),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1749),
.B(n_1764),
.Y(n_1833)
);

AO21x2_ASAP7_75t_L g1834 ( 
.A1(n_1655),
.A2(n_1670),
.B(n_1685),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1750),
.B(n_1651),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1733),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1638),
.B(n_1692),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1781),
.B(n_1688),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1828),
.B(n_1631),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1768),
.B(n_1666),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1803),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1773),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1793),
.B(n_1684),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1828),
.B(n_1698),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1828),
.B(n_1696),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1793),
.B(n_1775),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1803),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1775),
.B(n_1687),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1786),
.Y(n_1851)
);

INVx4_ASAP7_75t_L g1852 ( 
.A(n_1814),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1787),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1772),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1809),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1776),
.B(n_1826),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1790),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1772),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1679),
.Y(n_1859)
);

OAI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1778),
.A2(n_1716),
.B(n_1715),
.Y(n_1860)
);

INVxp67_ASAP7_75t_SL g1861 ( 
.A(n_1783),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1767),
.B(n_1678),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1832),
.B(n_1667),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1818),
.B(n_1693),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1832),
.B(n_1643),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1818),
.B(n_1760),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1653),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1826),
.B(n_1733),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1774),
.A2(n_1744),
.B1(n_1656),
.B2(n_1694),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1797),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1827),
.B(n_1742),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1827),
.B(n_1796),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1790),
.B(n_1706),
.Y(n_1873)
);

NOR2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1790),
.B(n_1707),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1778),
.A2(n_1716),
.B(n_1715),
.Y(n_1875)
);

AOI222xp33_ASAP7_75t_L g1876 ( 
.A1(n_1780),
.A2(n_1702),
.B1(n_1759),
.B2(n_1731),
.C1(n_1705),
.C2(n_1648),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1796),
.B(n_1695),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1837),
.B(n_1658),
.Y(n_1878)
);

OAI322xp33_ASAP7_75t_L g1879 ( 
.A1(n_1770),
.A2(n_1759),
.A3(n_1731),
.B1(n_1648),
.B2(n_1677),
.C1(n_1701),
.C2(n_1658),
.Y(n_1879)
);

OAI31xp33_ASAP7_75t_L g1880 ( 
.A1(n_1845),
.A2(n_1780),
.A3(n_1801),
.B(n_1822),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1854),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1841),
.A2(n_1774),
.B1(n_1805),
.B2(n_1812),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1843),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1876),
.A2(n_1808),
.B1(n_1805),
.B2(n_1812),
.Y(n_1884)
);

OAI31xp33_ASAP7_75t_L g1885 ( 
.A1(n_1845),
.A2(n_1801),
.A3(n_1822),
.B(n_1816),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1857),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1854),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1849),
.Y(n_1888)
);

A2O1A1Ixp33_ASAP7_75t_L g1889 ( 
.A1(n_1840),
.A2(n_1782),
.B(n_1795),
.C(n_1814),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1858),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1855),
.B(n_1825),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1862),
.B(n_1794),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1861),
.Y(n_1893)
);

OAI33xp33_ASAP7_75t_L g1894 ( 
.A1(n_1856),
.A2(n_1817),
.A3(n_1779),
.B1(n_1820),
.B2(n_1788),
.B3(n_1784),
.Y(n_1894)
);

NAND4xp25_ASAP7_75t_L g1895 ( 
.A(n_1871),
.B(n_1789),
.C(n_1791),
.D(n_1878),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1878),
.B(n_1829),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1841),
.A2(n_1808),
.B1(n_1805),
.B2(n_1812),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1848),
.B(n_1835),
.Y(n_1898)
);

OA21x2_ASAP7_75t_L g1899 ( 
.A1(n_1860),
.A2(n_1824),
.B(n_1802),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1852),
.A2(n_1819),
.B(n_1808),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1872),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_SL g1902 ( 
.A(n_1869),
.B(n_1785),
.C(n_1791),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_SL g1903 ( 
.A(n_1874),
.B(n_1829),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1859),
.B(n_1829),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1844),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1857),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1852),
.A2(n_1782),
.B1(n_1814),
.B2(n_1821),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1846),
.A2(n_1819),
.B1(n_1821),
.B2(n_1816),
.Y(n_1908)
);

AOI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1847),
.A2(n_1819),
.B1(n_1785),
.B2(n_1788),
.C(n_1784),
.Y(n_1909)
);

OAI211xp5_ASAP7_75t_L g1910 ( 
.A1(n_1850),
.A2(n_1789),
.B(n_1791),
.C(n_1771),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1852),
.A2(n_1819),
.B1(n_1815),
.B2(n_1834),
.Y(n_1911)
);

OAI221xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1850),
.A2(n_1789),
.B1(n_1785),
.B2(n_1835),
.C(n_1815),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1833),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1873),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1868),
.A2(n_1792),
.B1(n_1817),
.B2(n_1810),
.C(n_1779),
.Y(n_1915)
);

AO21x2_ASAP7_75t_L g1916 ( 
.A1(n_1875),
.A2(n_1823),
.B(n_1811),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1877),
.A2(n_1834),
.B1(n_1813),
.B2(n_1806),
.Y(n_1917)
);

OAI211xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1863),
.A2(n_1769),
.B(n_1830),
.C(n_1783),
.Y(n_1918)
);

INVx3_ASAP7_75t_SL g1919 ( 
.A(n_1839),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1870),
.A2(n_1792),
.B1(n_1777),
.B2(n_1820),
.C(n_1798),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1867),
.B(n_1654),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1859),
.B(n_1833),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1881),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1889),
.A2(n_1879),
.B(n_1836),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1883),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1884),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1887),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1897),
.A2(n_1867),
.B(n_1866),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1888),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1890),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1903),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1888),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1896),
.B(n_1891),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1909),
.A2(n_1807),
.B(n_1804),
.Y(n_1934)
);

OA21x2_ASAP7_75t_L g1935 ( 
.A1(n_1910),
.A2(n_1807),
.B(n_1804),
.Y(n_1935)
);

OA21x2_ASAP7_75t_L g1936 ( 
.A1(n_1920),
.A2(n_1811),
.B(n_1823),
.Y(n_1936)
);

NOR2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1914),
.B(n_1865),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1896),
.B(n_1838),
.Y(n_1938)
);

OR2x6_ASAP7_75t_L g1939 ( 
.A(n_1900),
.B(n_1831),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1919),
.B(n_1886),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1903),
.B(n_1862),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1898),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1916),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1898),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1891),
.B(n_1904),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1905),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1905),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1919),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1901),
.B(n_1842),
.Y(n_1949)
);

OR2x2_ASAP7_75t_SL g1950 ( 
.A(n_1902),
.B(n_1863),
.Y(n_1950)
);

INVxp67_ASAP7_75t_SL g1951 ( 
.A(n_1899),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1916),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1908),
.A2(n_1798),
.B(n_1853),
.Y(n_1953)
);

OR2x6_ASAP7_75t_L g1954 ( 
.A(n_1892),
.B(n_1831),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1931),
.B(n_1892),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1948),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1926),
.A2(n_1882),
.B1(n_1885),
.B2(n_1880),
.C(n_1911),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1935),
.Y(n_1958)
);

AOI211xp5_ASAP7_75t_L g1959 ( 
.A1(n_1924),
.A2(n_1889),
.B(n_1907),
.C(n_1912),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1926),
.A2(n_1894),
.B1(n_1915),
.B2(n_1917),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1931),
.B(n_1904),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1935),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1923),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1935),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1935),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1923),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1927),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1940),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1945),
.B(n_1922),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_L g1970 ( 
.A(n_1928),
.B(n_1895),
.C(n_1918),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1942),
.B(n_1913),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1935),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1936),
.B(n_1771),
.C(n_1800),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1942),
.B(n_1848),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1935),
.Y(n_1975)
);

NOR2x1p5_ASAP7_75t_L g1976 ( 
.A(n_1944),
.B(n_1914),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1950),
.Y(n_1977)
);

AND2x2_ASAP7_75t_SL g1978 ( 
.A(n_1953),
.B(n_1893),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1933),
.B(n_1938),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1954),
.B(n_1892),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1954),
.B(n_1886),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1952),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1950),
.B(n_1851),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1930),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1930),
.Y(n_1985)
);

INVx1_ASAP7_75t_SL g1986 ( 
.A(n_1940),
.Y(n_1986)
);

AND4x1_ASAP7_75t_L g1987 ( 
.A(n_1950),
.B(n_1921),
.C(n_1866),
.D(n_1864),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1925),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1953),
.A2(n_1777),
.B1(n_1834),
.B2(n_1810),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1952),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1952),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1943),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1943),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1929),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1963),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1956),
.B(n_1929),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1979),
.B(n_1938),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1979),
.B(n_1937),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1978),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1977),
.A2(n_1928),
.B(n_1953),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1961),
.B(n_1937),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1956),
.B(n_1932),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1974),
.B(n_1949),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1966),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1977),
.B(n_1974),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1988),
.B(n_1932),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1966),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1967),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1986),
.Y(n_2010)
);

NAND4xp25_ASAP7_75t_L g2011 ( 
.A(n_1968),
.B(n_1906),
.C(n_1941),
.D(n_1946),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1994),
.B(n_1946),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1967),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1994),
.B(n_1947),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1978),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1986),
.B(n_1947),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_1959),
.B(n_1953),
.C(n_1936),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1957),
.A2(n_1953),
.B1(n_1936),
.B2(n_1934),
.Y(n_2018)
);

NAND3xp33_ASAP7_75t_L g2019 ( 
.A(n_1959),
.B(n_1953),
.C(n_1936),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1978),
.B(n_1941),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1972),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1960),
.A2(n_1936),
.B1(n_1934),
.B2(n_1951),
.C(n_1939),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1972),
.Y(n_2023)
);

NAND2x2_ASAP7_75t_L g2024 ( 
.A(n_1968),
.B(n_1906),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_2017),
.A2(n_1970),
.B1(n_1960),
.B2(n_1936),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1995),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_2006),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_2010),
.Y(n_2028)
);

INVx1_ASAP7_75t_SL g2029 ( 
.A(n_2006),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_2019),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1996),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2021),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1997),
.B(n_1987),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1998),
.B(n_1955),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_2024),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2002),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2005),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2008),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2021),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_2003),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1998),
.B(n_1955),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_2020),
.B(n_1991),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1999),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2000),
.B(n_1984),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2009),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2023),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1997),
.B(n_1985),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_2016),
.Y(n_2048)
);

INVx4_ASAP7_75t_L g2049 ( 
.A(n_1999),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2020),
.B(n_1987),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2004),
.B(n_1971),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2001),
.B(n_1980),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2013),
.B(n_1985),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2001),
.B(n_1980),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2028),
.B(n_1968),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2027),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2027),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2028),
.B(n_1969),
.Y(n_2058)
);

O2A1O1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_2030),
.A2(n_2022),
.B(n_2015),
.C(n_1972),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_L g2060 ( 
.A(n_2025),
.B(n_2018),
.C(n_1973),
.Y(n_2060)
);

NAND3xp33_ASAP7_75t_SL g2061 ( 
.A(n_2050),
.B(n_2015),
.C(n_1989),
.Y(n_2061)
);

INVxp67_ASAP7_75t_SL g2062 ( 
.A(n_2030),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_2034),
.Y(n_2063)
);

AOI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2050),
.A2(n_1973),
.B(n_2011),
.C(n_1983),
.Y(n_2064)
);

AOI31xp33_ASAP7_75t_L g2065 ( 
.A1(n_2029),
.A2(n_2007),
.A3(n_2014),
.B(n_2012),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2030),
.A2(n_1989),
.B1(n_1972),
.B2(n_1962),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2034),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2043),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2043),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2049),
.B(n_1976),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_SL g2071 ( 
.A(n_2029),
.B(n_1981),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_2031),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2048),
.B(n_2031),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2048),
.B(n_1969),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2026),
.Y(n_2075)
);

OR3x2_ASAP7_75t_L g2076 ( 
.A(n_2051),
.B(n_1983),
.C(n_2024),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2026),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2063),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2068),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2067),
.B(n_2034),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_2062),
.B(n_2040),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2063),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2072),
.B(n_2040),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_2065),
.B(n_2034),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2069),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2058),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_2070),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2056),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_2071),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2057),
.Y(n_2090)
);

AOI222xp33_ASAP7_75t_L g2091 ( 
.A1(n_2061),
.A2(n_2044),
.B1(n_2050),
.B2(n_1964),
.C1(n_1962),
.C2(n_1975),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2072),
.B(n_2049),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2074),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2081),
.B(n_2055),
.Y(n_2094)
);

OAI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_2091),
.A2(n_2060),
.B1(n_2059),
.B2(n_2064),
.C(n_2044),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2080),
.B(n_2041),
.Y(n_2096)
);

AOI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_2081),
.A2(n_2076),
.B1(n_2073),
.B2(n_2066),
.C(n_2049),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2082),
.Y(n_2098)
);

NAND2x1_ASAP7_75t_L g2099 ( 
.A(n_2078),
.B(n_2042),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_L g2100 ( 
.A1(n_2084),
.A2(n_2071),
.B(n_2042),
.C(n_2035),
.Y(n_2100)
);

AOI221xp5_ASAP7_75t_SL g2101 ( 
.A1(n_2089),
.A2(n_2033),
.B1(n_2077),
.B2(n_2075),
.C(n_2037),
.Y(n_2101)
);

A2O1A1Ixp33_ASAP7_75t_L g2102 ( 
.A1(n_2084),
.A2(n_2042),
.B(n_2033),
.C(n_1965),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2078),
.B(n_2033),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2083),
.B(n_2049),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2092),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_L g2106 ( 
.A(n_2088),
.B(n_2042),
.C(n_2039),
.Y(n_2106)
);

OAI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2095),
.A2(n_1962),
.B1(n_1965),
.B2(n_1964),
.Y(n_2107)
);

INVxp67_ASAP7_75t_L g2108 ( 
.A(n_2094),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_2100),
.B(n_2042),
.Y(n_2109)
);

OA33x2_ASAP7_75t_L g2110 ( 
.A1(n_2103),
.A2(n_2047),
.A3(n_2086),
.B1(n_2090),
.B2(n_2093),
.B3(n_2085),
.Y(n_2110)
);

OAI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_2102),
.A2(n_2087),
.B(n_2079),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2097),
.A2(n_2035),
.B1(n_2041),
.B2(n_2032),
.Y(n_2112)
);

O2A1O1Ixp33_ASAP7_75t_SL g2113 ( 
.A1(n_2099),
.A2(n_2087),
.B(n_2035),
.C(n_2037),
.Y(n_2113)
);

AOI21xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2098),
.A2(n_2041),
.B(n_2038),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_2108),
.B(n_2096),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2111),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2114),
.B(n_2101),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_2110),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2109),
.B(n_2041),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_2112),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2113),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2107),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_2116),
.B(n_2105),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2118),
.A2(n_2106),
.B1(n_2104),
.B2(n_2032),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2118),
.B(n_2052),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2121),
.A2(n_2051),
.B1(n_2047),
.B2(n_2039),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2119),
.B(n_2052),
.Y(n_2127)
);

NAND4xp25_ASAP7_75t_L g2128 ( 
.A(n_2115),
.B(n_2054),
.C(n_2052),
.D(n_2032),
.Y(n_2128)
);

NOR2x1_ASAP7_75t_L g2129 ( 
.A(n_2125),
.B(n_2128),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2127),
.B(n_2054),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2124),
.B(n_2054),
.Y(n_2131)
);

NOR2x1_ASAP7_75t_L g2132 ( 
.A(n_2126),
.B(n_2117),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2130),
.Y(n_2133)
);

NOR3xp33_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_2120),
.C(n_2122),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2134),
.A2(n_2131),
.B1(n_2129),
.B2(n_2046),
.Y(n_2135)
);

AOI322xp5_ASAP7_75t_L g2136 ( 
.A1(n_2133),
.A2(n_2046),
.A3(n_2039),
.B1(n_1965),
.B2(n_1975),
.C1(n_1964),
.C2(n_1958),
.Y(n_2136)
);

CKINVDCx20_ASAP7_75t_R g2137 ( 
.A(n_2135),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2136),
.Y(n_2138)
);

NOR3xp33_ASAP7_75t_L g2139 ( 
.A(n_2138),
.B(n_2123),
.C(n_2046),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_SL g2140 ( 
.A1(n_2137),
.A2(n_2038),
.B(n_2036),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_2140),
.Y(n_2141)
);

AOI22x1_ASAP7_75t_L g2142 ( 
.A1(n_2139),
.A2(n_2045),
.B1(n_2036),
.B2(n_2023),
.Y(n_2142)
);

OAI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2141),
.A2(n_2045),
.B1(n_1991),
.B2(n_2053),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2143),
.B(n_2142),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2144),
.A2(n_1990),
.B(n_1982),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_1991),
.B1(n_2053),
.B2(n_1982),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2146),
.A2(n_1990),
.B1(n_1982),
.B2(n_1992),
.Y(n_2147)
);

AOI211xp5_ASAP7_75t_L g2148 ( 
.A1(n_2147),
.A2(n_1990),
.B(n_1992),
.C(n_1993),
.Y(n_2148)
);


endmodule