module real_aes_8744_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_841;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_532;
wire n_316;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_649;
wire n_293;
wire n_358;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_0), .A2(n_159), .B1(n_781), .B2(n_783), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_1), .A2(n_79), .B1(n_446), .B2(n_613), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_2), .A2(n_49), .B1(n_354), .B2(n_604), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_3), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_4), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_5), .A2(n_264), .B1(n_549), .B2(n_550), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_6), .A2(n_107), .B1(n_397), .B2(n_718), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_7), .A2(n_858), .B1(n_859), .B2(n_876), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_7), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_8), .A2(n_128), .B1(n_604), .B2(n_678), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_9), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_10), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_11), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_12), .A2(n_46), .B1(n_443), .B2(n_445), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_13), .A2(n_618), .B1(n_648), .B2(n_649), .Y(n_617) );
INVx1_ASAP7_75t_L g648 ( .A(n_13), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_14), .Y(n_726) );
INVx1_ASAP7_75t_L g732 ( .A(n_15), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_16), .A2(n_101), .B1(n_453), .B2(n_515), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_17), .A2(n_37), .B1(n_351), .B2(n_354), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_18), .A2(n_223), .B1(n_577), .B2(n_613), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_19), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_20), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_21), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_22), .A2(n_146), .B1(n_410), .B2(n_413), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_23), .A2(n_134), .B1(n_322), .B2(n_327), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_24), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_25), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_26), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_27), .A2(n_209), .B1(n_440), .B2(n_490), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_28), .A2(n_130), .B1(n_449), .B2(n_676), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_29), .A2(n_262), .B1(n_334), .B2(n_609), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_30), .Y(n_491) );
AO22x2_ASAP7_75t_L g295 ( .A1(n_31), .A2(n_94), .B1(n_296), .B2(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g854 ( .A(n_31), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_32), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_33), .A2(n_71), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_34), .A2(n_238), .B1(n_354), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_35), .A2(n_178), .B1(n_443), .B2(n_638), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_36), .A2(n_256), .B1(n_698), .B2(n_718), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_38), .A2(n_151), .B1(n_366), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_39), .A2(n_136), .B1(n_443), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_40), .A2(n_50), .B1(n_345), .B2(n_392), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_41), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_42), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_43), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g722 ( .A(n_44), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_45), .Y(n_730) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_47), .A2(n_95), .B1(n_296), .B2(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g855 ( .A(n_47), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_48), .A2(n_201), .B1(n_646), .B2(n_647), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_51), .A2(n_160), .B1(n_352), .B2(n_673), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_52), .Y(n_408) );
INVx1_ASAP7_75t_L g456 ( .A(n_53), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_54), .A2(n_243), .B1(n_518), .B2(n_519), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_55), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_56), .A2(n_197), .B1(n_440), .B2(n_613), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_57), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_58), .B(n_535), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_59), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_60), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_61), .A2(n_208), .B1(n_516), .B2(n_552), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_62), .A2(n_93), .B1(n_373), .B2(n_440), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_63), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_64), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_65), .A2(n_111), .B1(n_388), .B2(n_546), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_66), .A2(n_227), .B1(n_471), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_67), .A2(n_230), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_68), .A2(n_170), .B1(n_438), .B2(n_717), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_69), .A2(n_180), .B1(n_412), .B2(n_609), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_70), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_72), .A2(n_82), .B1(n_777), .B2(n_779), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_73), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_74), .B(n_728), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_75), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_76), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_77), .A2(n_138), .B1(n_322), .B2(n_466), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_78), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_80), .A2(n_220), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_81), .A2(n_129), .B1(n_373), .B2(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_83), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_84), .A2(n_190), .B1(n_577), .B2(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_85), .A2(n_106), .B1(n_391), .B2(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_86), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g614 ( .A1(n_87), .A2(n_158), .B1(n_167), .B2(n_532), .C1(n_563), .C2(n_615), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_88), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_89), .A2(n_90), .B1(n_440), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_91), .A2(n_192), .B1(n_613), .B2(n_678), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_92), .A2(n_150), .B1(n_419), .B2(n_423), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_96), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_97), .B(n_764), .Y(n_763) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_98), .A2(n_272), .B(n_281), .C(n_856), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_99), .A2(n_169), .B1(n_351), .B2(n_582), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_100), .Y(n_628) );
INVx1_ASAP7_75t_L g279 ( .A(n_102), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_103), .A2(n_194), .B1(n_391), .B2(n_393), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_104), .A2(n_251), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g633 ( .A(n_105), .Y(n_633) );
INVx1_ASAP7_75t_L g277 ( .A(n_108), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_109), .A2(n_171), .B1(n_371), .B2(n_440), .Y(n_611) );
INVx1_ASAP7_75t_L g631 ( .A(n_110), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_112), .A2(n_135), .B1(n_323), .B2(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_113), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_114), .A2(n_191), .B1(n_387), .B2(n_389), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_115), .A2(n_240), .B1(n_425), .B2(n_428), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_116), .A2(n_261), .B1(n_323), .B2(n_327), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_117), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_118), .A2(n_233), .B1(n_510), .B2(n_676), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_119), .Y(n_809) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_120), .A2(n_125), .B1(n_327), .B2(n_609), .Y(n_668) );
OA22x2_ASAP7_75t_L g655 ( .A1(n_121), .A2(n_656), .B1(n_657), .B2(n_679), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_121), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_122), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_123), .A2(n_222), .B1(n_584), .B2(n_587), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_124), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_126), .A2(n_218), .B1(n_449), .B2(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_127), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_131), .A2(n_133), .B1(n_600), .B2(n_601), .Y(n_599) );
OA22x2_ASAP7_75t_L g680 ( .A1(n_132), .A2(n_681), .B1(n_682), .B2(n_702), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_132), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_137), .A2(n_139), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_140), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_141), .B(n_765), .Y(n_866) );
XNOR2x2_ASAP7_75t_L g382 ( .A(n_142), .B(n_383), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_143), .Y(n_725) );
INVx2_ASAP7_75t_L g280 ( .A(n_144), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_145), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_147), .B(n_413), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_148), .A2(n_709), .B1(n_733), .B2(n_734), .Y(n_708) );
INVx1_ASAP7_75t_L g733 ( .A(n_148), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_149), .B(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_152), .A2(n_210), .B1(n_391), .B2(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_153), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_154), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_155), .Y(n_769) );
AND2x6_ASAP7_75t_L g276 ( .A(n_156), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_156), .Y(n_848) );
AO22x2_ASAP7_75t_L g305 ( .A1(n_157), .A2(n_221), .B1(n_296), .B2(n_300), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_161), .A2(n_185), .B1(n_438), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_162), .A2(n_234), .B1(n_417), .B2(n_421), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_163), .B(n_428), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_164), .A2(n_249), .B1(n_516), .B2(n_613), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_165), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_166), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_168), .A2(n_206), .B1(n_567), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_172), .A2(n_253), .B1(n_352), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_173), .A2(n_187), .B1(n_419), .B2(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_174), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_175), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_176), .B(n_421), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_177), .A2(n_204), .B1(n_345), .B2(n_346), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_179), .A2(n_245), .B1(n_642), .B2(n_676), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_181), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_182), .A2(n_270), .B1(n_543), .B2(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g559 ( .A(n_183), .Y(n_559) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_184), .A2(n_242), .B1(n_296), .B2(n_297), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_186), .A2(n_214), .B1(n_421), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_188), .A2(n_266), .B1(n_646), .B2(n_817), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_189), .A2(n_434), .B1(n_482), .B2(n_483), .Y(n_433) );
INVx1_ASAP7_75t_L g482 ( .A(n_189), .Y(n_482) );
AOI22xp5_ASAP7_75t_SL g554 ( .A1(n_193), .A2(n_555), .B1(n_589), .B2(n_590), .Y(n_554) );
INVx1_ASAP7_75t_L g590 ( .A(n_193), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_195), .A2(n_798), .B1(n_819), .B2(n_820), .Y(n_797) );
INVx1_ASAP7_75t_L g819 ( .A(n_195), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_196), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_198), .A2(n_225), .B1(n_392), .B2(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_199), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_200), .A2(n_244), .B1(n_322), .B2(n_539), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_202), .A2(n_226), .B1(n_322), .B2(n_327), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_203), .Y(n_623) );
INVx1_ASAP7_75t_L g568 ( .A(n_205), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_207), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_211), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_212), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_213), .A2(n_232), .B1(n_579), .B2(n_601), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_215), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_216), .Y(n_375) );
INVx1_ASAP7_75t_L g558 ( .A(n_217), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_219), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_221), .B(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_224), .B(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_228), .A2(n_260), .B1(n_453), .B2(n_601), .Y(n_639) );
INVx1_ASAP7_75t_L g823 ( .A(n_229), .Y(n_823) );
INVx1_ASAP7_75t_L g754 ( .A(n_231), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_235), .Y(n_553) );
INVx1_ASAP7_75t_L g565 ( .A(n_236), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_237), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_239), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_241), .B(n_471), .Y(n_629) );
INVx1_ASAP7_75t_L g851 ( .A(n_242), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_246), .A2(n_250), .B1(n_577), .B2(n_604), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g759 ( .A1(n_247), .A2(n_316), .B(n_760), .C(n_768), .Y(n_759) );
INVx1_ASAP7_75t_L g571 ( .A(n_248), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_252), .Y(n_360) );
INVx1_ASAP7_75t_L g296 ( .A(n_254), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_254), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_255), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_257), .Y(n_808) );
INVx1_ASAP7_75t_L g572 ( .A(n_258), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_259), .Y(n_338) );
OA22x2_ASAP7_75t_L g284 ( .A1(n_263), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_265), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_267), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_268), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_269), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_277), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_278), .A2(n_846), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_653), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_281) );
INVx1_ASAP7_75t_L g842 ( .A(n_282), .Y(n_842) );
XOR2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_380), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_342), .Y(n_287) );
NOR3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_313), .C(n_331), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_306), .B1(n_307), .B2(n_312), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_290), .A2(n_558), .B1(n_559), .B2(n_560), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_290), .A2(n_307), .B1(n_801), .B2(n_802), .Y(n_800) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g457 ( .A(n_291), .Y(n_457) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_292), .Y(n_499) );
BUFx3_ASAP7_75t_L g622 ( .A(n_292), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_292), .A2(n_309), .B1(n_832), .B2(n_833), .C(n_834), .Y(n_831) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
INVx2_ASAP7_75t_L g374 ( .A(n_293), .Y(n_374) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_294), .B(n_299), .Y(n_311) );
AND2x2_ASAP7_75t_L g353 ( .A(n_294), .B(n_337), .Y(n_353) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g318 ( .A(n_295), .B(n_299), .Y(n_318) );
AND2x2_ASAP7_75t_L g326 ( .A(n_295), .B(n_305), .Y(n_326) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_298), .Y(n_300) );
INVx2_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
INVx1_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_302), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g352 ( .A(n_302), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g427 ( .A(n_302), .B(n_374), .Y(n_427) );
AND2x6_ASAP7_75t_L g429 ( .A(n_302), .B(n_311), .Y(n_429) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
INVx1_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_303), .B(n_305), .Y(n_358) );
AND2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g349 ( .A(n_305), .B(n_330), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_307), .A2(n_496), .B1(n_497), .B2(n_500), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_307), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_309), .A2(n_499), .B1(n_722), .B2(n_723), .Y(n_721) );
BUFx3_ASAP7_75t_L g762 ( .A(n_309), .Y(n_762) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g460 ( .A(n_310), .Y(n_460) );
AND2x4_ASAP7_75t_L g345 ( .A(n_311), .B(n_319), .Y(n_345) );
AND2x2_ASAP7_75t_L g348 ( .A(n_311), .B(n_349), .Y(n_348) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_321), .Y(n_313) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_315), .A2(n_660), .B(n_661), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g835 ( .A1(n_315), .A2(n_836), .B(n_837), .Y(n_835) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g407 ( .A(n_317), .Y(n_407) );
INVx2_ASAP7_75t_SL g462 ( .A(n_317), .Y(n_462) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_317), .Y(n_490) );
INVx4_ASAP7_75t_L g564 ( .A(n_317), .Y(n_564) );
INVx2_ASAP7_75t_L g625 ( .A(n_317), .Y(n_625) );
AND2x6_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g480 ( .A(n_318), .Y(n_480) );
AND2x2_ASAP7_75t_L g363 ( .A(n_319), .B(n_353), .Y(n_363) );
AND2x6_ASAP7_75t_L g373 ( .A(n_319), .B(n_374), .Y(n_373) );
BUFx4f_ASAP7_75t_SL g615 ( .A(n_322), .Y(n_615) );
INVx2_ASAP7_75t_L g773 ( .A(n_322), .Y(n_773) );
BUFx12f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_323), .Y(n_414) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_323), .Y(n_471) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g336 ( .A(n_325), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g335 ( .A(n_326), .B(n_336), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_326), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g419 ( .A(n_326), .B(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_328), .Y(n_423) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_328), .Y(n_532) );
INVx1_ASAP7_75t_L g481 ( .A(n_329), .Y(n_481) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_338), .B2(n_339), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g803 ( .A1(n_333), .A2(n_562), .B1(n_804), .B2(n_805), .C(n_806), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_335), .Y(n_412) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_335), .Y(n_466) );
BUFx4f_ASAP7_75t_SL g539 ( .A(n_335), .Y(n_539) );
BUFx2_ASAP7_75t_L g567 ( .A(n_335), .Y(n_567) );
INVx1_ASAP7_75t_L g341 ( .A(n_337), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_339), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx4_ASAP7_75t_L g475 ( .A(n_340), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_340), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_570) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_340), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_340), .A2(n_627), .B1(n_745), .B2(n_746), .Y(n_744) );
AND2x2_ASAP7_75t_L g552 ( .A(n_341), .B(n_368), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_359), .C(n_369), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_350), .Y(n_343) );
INVx6_ASAP7_75t_L g403 ( .A(n_345), .Y(n_403) );
BUFx3_ASAP7_75t_L g438 ( .A(n_345), .Y(n_438) );
BUFx3_ASAP7_75t_L g586 ( .A(n_345), .Y(n_586) );
BUFx3_ASAP7_75t_L g698 ( .A(n_345), .Y(n_698) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx4_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
INVx5_ASAP7_75t_L g516 ( .A(n_347), .Y(n_516) );
INVx3_ASAP7_75t_L g550 ( .A(n_347), .Y(n_550) );
BUFx3_ASAP7_75t_L g602 ( .A(n_347), .Y(n_602) );
INVx8_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_349), .B(n_353), .Y(n_379) );
AND2x2_ASAP7_75t_L g441 ( .A(n_349), .B(n_353), .Y(n_441) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
INVx2_ASAP7_75t_L g444 ( .A(n_352), .Y(n_444) );
BUFx3_ASAP7_75t_L g518 ( .A(n_352), .Y(n_518) );
BUFx3_ASAP7_75t_L g604 ( .A(n_352), .Y(n_604) );
AND2x4_ASAP7_75t_L g367 ( .A(n_353), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
BUFx4f_ASAP7_75t_SL g453 ( .A(n_355), .Y(n_453) );
BUFx2_ASAP7_75t_L g519 ( .A(n_355), .Y(n_519) );
BUFx2_ASAP7_75t_L g579 ( .A(n_355), .Y(n_579) );
INVx6_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g673 ( .A(n_356), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_356), .A2(n_479), .B1(n_692), .B2(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g783 ( .A(n_356), .Y(n_783) );
OR2x6_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g420 ( .A(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g368 ( .A(n_358), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_364), .B2(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
INVx2_ASAP7_75t_L g511 ( .A(n_363), .Y(n_511) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_SL g389 ( .A(n_367), .Y(n_389) );
BUFx3_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
BUFx3_ASAP7_75t_L g546 ( .A(n_367), .Y(n_546) );
BUFx3_ASAP7_75t_L g577 ( .A(n_367), .Y(n_577) );
BUFx2_ASAP7_75t_L g678 ( .A(n_367), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_375), .B1(n_376), .B2(n_377), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx5_ASAP7_75t_SL g397 ( .A(n_372), .Y(n_397) );
INVx4_ASAP7_75t_L g543 ( .A(n_372), .Y(n_543) );
INVx2_ASAP7_75t_L g582 ( .A(n_372), .Y(n_582) );
INVx11_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx11_ASAP7_75t_L g451 ( .A(n_373), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_377), .A2(n_402), .B1(n_403), .B2(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g788 ( .A(n_378), .Y(n_788) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
XOR2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_522), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_430), .B1(n_431), .B2(n_521), .Y(n_381) );
INVx2_ASAP7_75t_L g521 ( .A(n_382), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_384), .B(n_405), .Y(n_383) );
NOR3xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_394), .C(n_401), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g449 ( .A(n_388), .Y(n_449) );
BUFx3_ASAP7_75t_L g638 ( .A(n_388), .Y(n_638) );
INVx3_ASAP7_75t_L g778 ( .A(n_388), .Y(n_778) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g782 ( .A(n_392), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_397), .Y(n_779) );
INVx4_ASAP7_75t_L g646 ( .A(n_399), .Y(n_646) );
INVx4_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g514 ( .A(n_403), .Y(n_514) );
INVx2_ASAP7_75t_L g549 ( .A(n_403), .Y(n_549) );
INVx2_ASAP7_75t_L g600 ( .A(n_403), .Y(n_600) );
INVx3_ASAP7_75t_L g642 ( .A(n_403), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_415), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B(n_409), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g862 ( .A1(n_407), .A2(n_863), .B(n_864), .Y(n_862) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx4f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g492 ( .A(n_414), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_424), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g609 ( .A(n_419), .Y(n_609) );
BUFx2_ASAP7_75t_L g690 ( .A(n_419), .Y(n_690) );
BUFx2_ASAP7_75t_L g767 ( .A(n_419), .Y(n_767) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g535 ( .A(n_426), .Y(n_535) );
INVx5_ASAP7_75t_L g667 ( .A(n_426), .Y(n_667) );
INVx2_ASAP7_75t_L g765 ( .A(n_426), .Y(n_765) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx4f_ASAP7_75t_L g537 ( .A(n_429), .Y(n_537) );
INVx1_ASAP7_75t_SL g665 ( .A(n_429), .Y(n_665) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B1(n_484), .B2(n_485), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_435), .B(n_454), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_447), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_442), .Y(n_436) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g644 ( .A(n_440), .Y(n_644) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g544 ( .A(n_441), .Y(n_544) );
BUFx3_ASAP7_75t_L g718 ( .A(n_441), .Y(n_718) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_444), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_445), .Y(n_792) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_SL g508 ( .A(n_451), .Y(n_508) );
INVx4_ASAP7_75t_L g676 ( .A(n_451), .Y(n_676) );
OAI21xp33_ASAP7_75t_SL g687 ( .A1(n_451), .A2(n_688), .B(n_689), .Y(n_687) );
INVx4_ASAP7_75t_L g714 ( .A(n_451), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_461), .C(n_472), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_455) );
OA211x2_ASAP7_75t_L g605 ( .A1(n_459), .A2(n_606), .B(n_607), .C(n_608), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_459), .A2(n_622), .B1(n_685), .B2(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g560 ( .A(n_460), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_464), .B2(n_467), .C(n_468), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_464), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g627 ( .A(n_465), .Y(n_627) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g728 ( .A(n_471), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_476), .B2(n_477), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_SL g632 ( .A(n_475), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_477), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_477), .A2(n_632), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g573 ( .A(n_478), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g634 ( .A(n_479), .Y(n_634) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
XOR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_520), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_505), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_495), .C(n_501), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_491), .B1(n_492), .B2(n_493), .C(n_494), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_489), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g613 ( .A(n_511), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_591), .B1(n_651), .B2(n_652), .Y(n_522) );
INVx4_ASAP7_75t_L g651 ( .A(n_523), .Y(n_651) );
XOR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_554), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
XOR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_553), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_528), .B(n_540), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .C(n_538), .Y(n_533) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_547), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
INVx1_ASAP7_75t_L g588 ( .A(n_544), .Y(n_588) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
INVx2_ASAP7_75t_L g818 ( .A(n_546), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVxp67_ASAP7_75t_L g786 ( .A(n_549), .Y(n_786) );
INVx1_ASAP7_75t_SL g589 ( .A(n_555), .Y(n_589) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_556), .B(n_574), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_570), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_560), .A2(n_622), .B1(n_739), .B2(n_740), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_565), .B1(n_566), .B2(n_568), .C(n_569), .Y(n_561) );
OAI221xp5_ASAP7_75t_SL g724 ( .A1(n_562), .A2(n_566), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g741 ( .A1(n_564), .A2(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g652 ( .A(n_592), .Y(n_652) );
OAI22xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_617), .B2(n_650), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
XOR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_616), .Y(n_596) );
NAND4xp75_ASAP7_75t_L g597 ( .A(n_598), .B(n_605), .C(n_610), .D(n_614), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_603), .Y(n_598) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g650 ( .A(n_617), .Y(n_650) );
INVx2_ASAP7_75t_L g649 ( .A(n_618), .Y(n_649) );
AND2x2_ASAP7_75t_SL g618 ( .A(n_619), .B(n_635), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_624), .C(n_630), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_627), .B2(n_628), .C(n_629), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_640), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g841 ( .A(n_653), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_703), .B1(n_704), .B2(n_840), .Y(n_653) );
INVx1_ASAP7_75t_L g840 ( .A(n_654), .Y(n_840) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_680), .Y(n_654) );
INVx1_ASAP7_75t_L g679 ( .A(n_657), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_669), .Y(n_657) );
NOR2xp67_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .C(n_668), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g702 ( .A(n_682), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_694), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .C(n_691), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_699), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_795), .B1(n_838), .B2(n_839), .Y(n_704) );
INVx1_ASAP7_75t_L g838 ( .A(n_705), .Y(n_838) );
OAI22xp5_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_756), .B1(n_793), .B2(n_794), .Y(n_705) );
INVx1_ASAP7_75t_L g793 ( .A(n_706), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_735), .B2(n_755), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g734 ( .A(n_709), .Y(n_734) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_710), .B(n_720), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .Y(n_710) );
NAND2xp33_ASAP7_75t_SL g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
BUFx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .C(n_729), .Y(n_720) );
INVx1_ASAP7_75t_L g755 ( .A(n_735), .Y(n_755) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_754), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_747), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .C(n_744), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g794 ( .A(n_756), .Y(n_794) );
XNOR2x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_774), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B(n_763), .C(n_766), .Y(n_760) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_784), .C(n_789), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_780), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_784) );
INVx2_ASAP7_75t_L g839 ( .A(n_795), .Y(n_839) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_797), .B1(n_821), .B2(n_822), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g820 ( .A(n_798), .Y(n_820) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_810), .Y(n_798) );
NOR3xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_803), .C(n_807), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
XNOR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
NOR4xp75_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .C(n_831), .D(n_835), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_826), .B(n_827), .Y(n_825) );
NAND2xp5_ASAP7_75t_SL g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_845), .B(n_849), .Y(n_844) );
OR2x2_ASAP7_75t_SL g890 ( .A(n_845), .B(n_850), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_846), .Y(n_879) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_847), .B(n_882), .Y(n_885) );
CKINVDCx16_ASAP7_75t_R g882 ( .A(n_848), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
OAI322xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_877), .A3(n_880), .B1(n_883), .B2(n_886), .C1(n_887), .C2(n_888), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
XOR2x2_ASAP7_75t_L g887 ( .A(n_860), .B(n_886), .Y(n_887) );
NAND2x1_ASAP7_75t_SL g860 ( .A(n_861), .B(n_869), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_865), .Y(n_861) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .C(n_868), .Y(n_865) );
NOR2x1_ASAP7_75t_L g869 ( .A(n_870), .B(n_873), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
CKINVDCx16_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
endmodule