module fake_jpeg_16549_n_146 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_40),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_24),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_17),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_49),
.B(n_14),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_18),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_0),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_27),
.A3(n_20),
.B1(n_52),
.B2(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_74),
.B1(n_77),
.B2(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_55),
.C(n_17),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_45),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_27),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_87),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_92),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_20),
.C(n_13),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_57),
.C(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.C(n_104),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_51),
.B1(n_47),
.B2(n_82),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_58),
.C(n_60),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_58),
.B(n_62),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_103),
.B(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_59),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_60),
.B(n_51),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_70),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_67),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_78),
.B1(n_79),
.B2(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_116),
.B1(n_102),
.B2(n_101),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_78),
.B(n_80),
.C(n_83),
.D(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_12),
.A3(n_7),
.B1(n_8),
.B2(n_11),
.C1(n_24),
.C2(n_25),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_94),
.C(n_97),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_108),
.C(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_116),
.B1(n_111),
.B2(n_118),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_129),
.Y(n_135)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_28),
.A3(n_4),
.B1(n_3),
.B2(n_11),
.C(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_132),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_28),
.C(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_136),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_124),
.B(n_123),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_3),
.B(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_119),
.C(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_119),
.Y(n_140)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_141),
.B(n_134),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_143),
.B(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_142),
.Y(n_146)
);


endmodule