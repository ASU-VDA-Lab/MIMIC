module fake_netlist_6_4129_n_4945 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4945);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4945;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_2332;
wire n_3849;
wire n_578;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_3222;
wire n_1387;
wire n_677;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_3030;
wire n_830;
wire n_2838;
wire n_3427;
wire n_852;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_544;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_1660;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_2011;
wire n_564;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_608;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_1290;
wire n_2072;
wire n_1354;
wire n_586;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_604;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_687;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_595;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_2145;
wire n_898;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_925;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_532;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_536;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_581;
wire n_4713;
wire n_4098;
wire n_4476;
wire n_3700;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_648;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_4541;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_552;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_2296;
wire n_3633;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_3331;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_589;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4069;
wire n_2748;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_556;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_3724;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_2552;
wire n_1053;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_858;
wire n_2049;
wire n_956;
wire n_663;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_664;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_2016;
wire n_4470;
wire n_580;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_607;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_974;
wire n_2656;
wire n_2375;
wire n_1934;
wire n_628;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_662;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_533;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_4242;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_545;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_568;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_573;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_1460;
wire n_911;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_633;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_629;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_3340;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_616;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_666;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4563;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_3765;
wire n_4125;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_3639;
wire n_4334;
wire n_659;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_551;
wire n_699;
wire n_4320;
wire n_3884;
wire n_757;
wire n_594;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_2850;
wire n_572;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_530;
wire n_4319;
wire n_3369;
wire n_618;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_612;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_593;
wire n_637;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_2517;
wire n_2713;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_1959;
wire n_3133;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_631;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_623;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_546;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_688;
wire n_1077;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_602;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_587;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_575;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_557;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_3449;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_597;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_621;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_624;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_599;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_543;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_3517;
wire n_4045;
wire n_3893;
wire n_4598;
wire n_2945;
wire n_3061;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_1860;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_566;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_671;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_676;
wire n_832;
wire n_3049;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_1392;
wire n_4495;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_611;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_930;
wire n_2620;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_576;
wire n_2683;
wire n_563;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_626;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_570;
wire n_1789;
wire n_620;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_2334;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_635;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_571;
wire n_2215;
wire n_1884;
wire n_665;
wire n_2055;
wire n_2553;
wire n_632;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_681;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_3079;
wire n_4360;
wire n_540;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_531;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_1003;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_539;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_638;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_577;
wire n_1843;
wire n_619;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_606;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_630;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_549;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_689;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_1988;
wire n_558;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_690;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_678;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_590;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_1634;
wire n_3252;
wire n_627;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_2913;
wire n_840;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_3789;
wire n_605;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_2537;
wire n_4483;
wire n_4661;
wire n_1308;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_1469;
wire n_2650;
wire n_987;
wire n_720;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_656;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_3580;
wire n_2842;
wire n_2335;
wire n_529;
wire n_2307;
wire n_3704;
wire n_684;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_2877;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_562;
wire n_2323;
wire n_2784;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_651;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_983;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_613;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_554;
wire n_1995;
wire n_3751;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1841;
wire n_4660;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_3417;
wire n_4124;
wire n_785;
wire n_609;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_579;
wire n_2789;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_565;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_654;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_584;
wire n_2141;
wire n_548;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_652;
wire n_4604;
wire n_3305;
wire n_1906;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_655;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_591;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_680;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_2814;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_535;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_553;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_679;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_4275;
wire n_1915;
wire n_4283;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_649;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_625;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_1572;
wire n_4308;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_1163;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_2090;
wire n_2603;
wire n_538;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_2108;
wire n_1211;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_2985;
wire n_1978;
wire n_574;
wire n_3792;
wire n_4202;
wire n_3938;
wire n_1446;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_559;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_645;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_541;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_821;
wire n_4372;
wire n_1068;
wire n_982;
wire n_2831;
wire n_932;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_547;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_674;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_702;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_598;
wire n_4169;
wire n_697;
wire n_3271;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_585;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_673;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_542;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_622;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_3148;
wire n_4022;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_657;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_526;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_527;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_600;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_1339;
wire n_2475;
wire n_723;
wire n_3144;
wire n_3244;
wire n_596;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_2357;
wire n_2025;
wire n_4654;
wire n_3640;
wire n_642;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_1618;
wire n_4867;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_3749;
wire n_2942;
wire n_4714;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_617;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_610;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_4182;
wire n_667;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_603;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_4590;
wire n_2543;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_4888;
wire n_1823;
wire n_2479;
wire n_776;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_1456;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_560;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_569;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_3156;
wire n_672;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_636;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_646;
wire n_528;
wire n_1329;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_1759;
wire n_853;
wire n_875;
wire n_1678;
wire n_661;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_555;
wire n_4579;
wire n_669;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4911;
wire n_4436;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_647;
wire n_844;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_3456;
wire n_1537;
wire n_779;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_4142;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_592;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_582;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_588;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g526 ( 
.A(n_68),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_477),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_81),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_494),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_134),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_294),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_296),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_215),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_423),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_200),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_139),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_30),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_246),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_163),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_506),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_177),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_483),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_486),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_67),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_425),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_56),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_84),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_338),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_280),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_40),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_406),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_322),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_457),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_156),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_500),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_377),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_104),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_263),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_149),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_229),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_308),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_90),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_40),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_29),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_75),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_94),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_85),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_94),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_286),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_493),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_309),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_38),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_323),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_502),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_307),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_426),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_313),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_434),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_360),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_121),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_189),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_14),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_21),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_452),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_98),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_293),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_138),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_518),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_141),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_90),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_75),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_124),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_283),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_363),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_400),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_435),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_454),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_357),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_218),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_165),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_275),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_208),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_370),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_227),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_390),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_460),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_272),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_480),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_318),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_231),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_227),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_312),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_401),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_295),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_179),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_160),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_326),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_356),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_283),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_243),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_53),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_107),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_52),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_519),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_64),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_380),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_149),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_378),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_501),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_99),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_233),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_404),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_245),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_43),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_451),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_50),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_156),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_226),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_397),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_10),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_327),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_61),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_158),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_137),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_189),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_275),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_132),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_176),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_35),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_234),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_485),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_419),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_167),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_204),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_447),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_145),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_290),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_154),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_495),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_168),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_41),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_376),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_240),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_9),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_215),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_54),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_164),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_74),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_93),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_487),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_186),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_315),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_219),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_272),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_398),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_251),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_144),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_499),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_488),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_239),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_347),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_430),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_478),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_34),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_241),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_136),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_330),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_358),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_301),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_405),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_131),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_172),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_399),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_89),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_72),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_492),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_173),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_271),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_44),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_133),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_441),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_288),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_53),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_96),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_77),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_163),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_302),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_424),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_105),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_248),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_118),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_136),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_408),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_414),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_348),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_228),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_342),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_17),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_496),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_429),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_178),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_104),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_43),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_50),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_192),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_394),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_113),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_415),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_12),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_211),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_250),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_121),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_161),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_225),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_442),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_465),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_107),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_126),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_214),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_76),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_332),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_135),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_135),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_230),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_59),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_286),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_95),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_521),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_51),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_221),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_42),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_159),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_407),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_240),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_362),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_511),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_371),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_0),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_418),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_462),
.Y(n_770)
);

BUFx5_ASAP7_75t_L g771 ( 
.A(n_194),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_306),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_159),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_469),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_260),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_32),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_448),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_182),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_57),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_79),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_449),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_292),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_119),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_72),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_364),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_35),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_64),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_133),
.Y(n_788)
);

CKINVDCx14_ASAP7_75t_R g789 ( 
.A(n_38),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_164),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_439),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_244),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_196),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_420),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_474),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_343),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_125),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_261),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_1),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_236),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_63),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_30),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_31),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_491),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_221),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_497),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_431),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_51),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_316),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_131),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_204),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_249),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_382),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_22),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_86),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_138),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_241),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_158),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_248),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_132),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_255),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_80),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_79),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_200),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_387),
.Y(n_825)
);

BUFx8_ASAP7_75t_SL g826 ( 
.A(n_250),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_314),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_339),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_109),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_168),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_417),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_208),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_440),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_473),
.Y(n_834)
);

BUFx10_ASAP7_75t_L g835 ( 
.A(n_157),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_436),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_63),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_510),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_54),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_152),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_374),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_453),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_375),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_247),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_37),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_464),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_150),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_266),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_5),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_516),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_174),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_92),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_513),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_379),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_218),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_157),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_279),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_161),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_95),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_36),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_386),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_458),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_350),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_334),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_212),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_205),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_484),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_194),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_86),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_228),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_206),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_359),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_183),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_196),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_289),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_455),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_58),
.Y(n_877)
);

BUFx10_ASAP7_75t_L g878 ( 
.A(n_220),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_58),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_180),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_244),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_388),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_24),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_395),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_233),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_368),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_260),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_212),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_366),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_1),
.Y(n_890)
);

BUFx5_ASAP7_75t_L g891 ( 
.A(n_192),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_3),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_18),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_311),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_211),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_97),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_60),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_46),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_66),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_269),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_466),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_367),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_253),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_181),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_280),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_137),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_335),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_489),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_122),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_461),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_59),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_413),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_261),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_254),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_252),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_463),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_153),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_365),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_57),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_187),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_433),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_445),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_170),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_270),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_443),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_197),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_67),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_39),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_384),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_276),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_427),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_373),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_372),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_337),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_304),
.Y(n_935)
);

BUFx8_ASAP7_75t_SL g936 ( 
.A(n_329),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_291),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_276),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_229),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_105),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_352),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_12),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_39),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_355),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_284),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_85),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_459),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_145),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_344),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_82),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_490),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_219),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_122),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_264),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_361),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_369),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_220),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_42),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_236),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_89),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_155),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_41),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_185),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_321),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_170),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_237),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_14),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_36),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_81),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_381),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_771),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_532),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_771),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_771),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_771),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_771),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_771),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_771),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_575),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_535),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_826),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_771),
.Y(n_982)
);

INVxp33_ASAP7_75t_SL g983 ( 
.A(n_614),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_707),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_891),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_891),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_560),
.Y(n_987)
);

INVxp33_ASAP7_75t_SL g988 ( 
.A(n_647),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_891),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_753),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_936),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_891),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_891),
.Y(n_993)
);

INVxp33_ASAP7_75t_SL g994 ( 
.A(n_708),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_754),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_891),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_563),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_891),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_891),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_632),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_632),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_686),
.Y(n_1002)
);

INVxp33_ASAP7_75t_L g1003 ( 
.A(n_756),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_643),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_643),
.Y(n_1005)
);

CKINVDCx14_ASAP7_75t_R g1006 ( 
.A(n_789),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_875),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_575),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_654),
.Y(n_1009)
);

INVxp33_ASAP7_75t_SL g1010 ( 
.A(n_528),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_710),
.Y(n_1011)
);

INVxp33_ASAP7_75t_L g1012 ( 
.A(n_810),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_710),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_686),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_686),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_618),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_686),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_686),
.Y(n_1018)
);

INVxp33_ASAP7_75t_SL g1019 ( 
.A(n_528),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_743),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_743),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_622),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_743),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_911),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_743),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_752),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_752),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_585),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_530),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_752),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_752),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_623),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_868),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_868),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_583),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

INVxp33_ASAP7_75t_L g1037 ( 
.A(n_548),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_868),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_868),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_586),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_896),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_896),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_896),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_896),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_896),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_909),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_909),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_909),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_621),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_909),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_909),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_526),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_548),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_533),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_620),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_544),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_591),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_546),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_551),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_566),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_599),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_570),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_530),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_556),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_539),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_626),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_547),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_636),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_587),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_565),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_633),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_593),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_639),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_583),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_596),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_598),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_605),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_606),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_608),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_629),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_583),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_613),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_630),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_646),
.B(n_817),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_663),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_640),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_631),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_577),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_841),
.B(n_0),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_642),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_634),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_539),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_539),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_653),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_635),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_666),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_668),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_674),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_556),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_583),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_595),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_613),
.Y(n_1102)
);

CKINVDCx16_ASAP7_75t_R g1103 ( 
.A(n_595),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_676),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_679),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_637),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_684),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_683),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_687),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_716),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_721),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_722),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_733),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_595),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_724),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_735),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_821),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_737),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_701),
.Y(n_1119)
);

INVxp33_ASAP7_75t_SL g1120 ( 
.A(n_536),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_741),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_747),
.Y(n_1122)
);

INVxp33_ASAP7_75t_SL g1123 ( 
.A(n_536),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_760),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_638),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_713),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_761),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_778),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_537),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_788),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_790),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_739),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_801),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_803),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_537),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_812),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_814),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_641),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_823),
.Y(n_1139)
);

CKINVDCx14_ASAP7_75t_R g1140 ( 
.A(n_746),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_830),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_847),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_848),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_568),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_869),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_644),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_682),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_879),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_880),
.Y(n_1149)
);

INVxp33_ASAP7_75t_SL g1150 ( 
.A(n_538),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_583),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_682),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_648),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_890),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_895),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_650),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_538),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_897),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_759),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_898),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_920),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_927),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_939),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_841),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_652),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_841),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_784),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_942),
.Y(n_1168)
);

INVxp33_ASAP7_75t_L g1169 ( 
.A(n_568),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_945),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_950),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_821),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_953),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_552),
.B(n_2),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_541),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_799),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_968),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_829),
.Y(n_1178)
);

INVxp67_ASAP7_75t_SL g1179 ( 
.A(n_908),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_969),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_550),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_555),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_656),
.Y(n_1183)
);

INVxp33_ASAP7_75t_SL g1184 ( 
.A(n_541),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_561),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_562),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_578),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_580),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_912),
.Y(n_1189)
);

INVxp67_ASAP7_75t_SL g1190 ( 
.A(n_584),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_588),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_600),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_612),
.Y(n_1193)
);

INVxp33_ASAP7_75t_SL g1194 ( 
.A(n_559),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_619),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_617),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_627),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_657),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_628),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_559),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_645),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_579),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_564),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_603),
.B(n_2),
.Y(n_1204)
);

INVxp33_ASAP7_75t_SL g1205 ( 
.A(n_564),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_649),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_662),
.Y(n_1207)
);

INVxp33_ASAP7_75t_SL g1208 ( 
.A(n_567),
.Y(n_1208)
);

BUFx2_ASAP7_75t_SL g1209 ( 
.A(n_553),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_821),
.Y(n_1210)
);

INVxp33_ASAP7_75t_SL g1211 ( 
.A(n_567),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_700),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_658),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_703),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_712),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_579),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_723),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_725),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_837),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_L g1220 ( 
.A(n_893),
.B(n_3),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_617),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_659),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_727),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_751),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_873),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_660),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_835),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_769),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_774),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_601),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_785),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_831),
.Y(n_1232)
);

CKINVDCx16_ASAP7_75t_R g1233 ( 
.A(n_835),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_838),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_655),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_655),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_850),
.Y(n_1237)
);

CKINVDCx16_ASAP7_75t_R g1238 ( 
.A(n_835),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_876),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_882),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_884),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_904),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_905),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_571),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_889),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_601),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_664),
.Y(n_1247)
);

INVxp33_ASAP7_75t_SL g1248 ( 
.A(n_571),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_878),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_910),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_918),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_941),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_625),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_603),
.B(n_615),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_625),
.Y(n_1255)
);

INVxp33_ASAP7_75t_SL g1256 ( 
.A(n_572),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_689),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_689),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_770),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_770),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_781),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_878),
.Y(n_1262)
);

INVxp33_ASAP7_75t_SL g1263 ( 
.A(n_572),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_781),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_670),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_864),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_671),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_864),
.Y(n_1268)
);

INVxp33_ASAP7_75t_SL g1269 ( 
.A(n_573),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_901),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_901),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_694),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_694),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_793),
.Y(n_1274)
);

INVxp33_ASAP7_75t_L g1275 ( 
.A(n_793),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_615),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_800),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_711),
.B(n_4),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_800),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_573),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_815),
.Y(n_1281)
);

CKINVDCx14_ASAP7_75t_R g1282 ( 
.A(n_579),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_711),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_815),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_881),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_881),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_887),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_887),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_854),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_854),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_903),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_952),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_903),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_919),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_919),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_928),
.Y(n_1296)
);

INVxp33_ASAP7_75t_SL g1297 ( 
.A(n_576),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_929),
.Y(n_1298)
);

CKINVDCx14_ASAP7_75t_R g1299 ( 
.A(n_672),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_960),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_928),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_929),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_963),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_956),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_878),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_963),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_956),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_646),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_616),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_817),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_926),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_926),
.Y(n_1312)
);

INVxp33_ASAP7_75t_SL g1313 ( 
.A(n_576),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_967),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_940),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_940),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_569),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_651),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_673),
.Y(n_1319)
);

BUFx2_ASAP7_75t_SL g1320 ( 
.A(n_624),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_675),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_677),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_601),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_661),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_719),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_678),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_681),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_690),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_695),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_696),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_601),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_702),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_672),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_589),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_669),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_601),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_704),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_705),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_589),
.Y(n_1339)
);

INVxp33_ASAP7_75t_L g1340 ( 
.A(n_796),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_709),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_680),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_714),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_715),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_720),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_672),
.Y(n_1346)
);

BUFx8_ASAP7_75t_SL g1347 ( 
.A(n_597),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_796),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_796),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_665),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_728),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_796),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_731),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_732),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1152),
.B(n_979),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1002),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1035),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1349),
.A2(n_740),
.B(n_734),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_1350),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1035),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1055),
.B(n_685),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1014),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1035),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1035),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_991),
.Y(n_1365)
);

BUFx12f_ASAP7_75t_L g1366 ( 
.A(n_987),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1015),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1074),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1325),
.Y(n_1369)
);

AND2x2_ASAP7_75t_SL g1370 ( 
.A(n_1204),
.B(n_796),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1164),
.B(n_531),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1074),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_979),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1008),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1074),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1071),
.B(n_1095),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1017),
.Y(n_1377)
);

BUFx8_ASAP7_75t_SL g1378 ( 
.A(n_981),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_978),
.A2(n_949),
.B(n_791),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1018),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1074),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1276),
.B(n_667),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1021),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_980),
.Y(n_1384)
);

BUFx8_ASAP7_75t_L g1385 ( 
.A(n_1129),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1008),
.B(n_791),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1081),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1166),
.B(n_836),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1081),
.Y(n_1389)
);

NOR2x1_ASAP7_75t_L g1390 ( 
.A(n_1089),
.B(n_1323),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1082),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1081),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_978),
.A2(n_949),
.B(n_791),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1016),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_987),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1081),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1100),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1100),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1002),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1100),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_995),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1023),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1349),
.A2(n_744),
.B(n_742),
.Y(n_1403)
);

CKINVDCx6p67_ASAP7_75t_R g1404 ( 
.A(n_1009),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_971),
.A2(n_750),
.B(n_748),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1020),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1100),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1209),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1331),
.B(n_916),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1082),
.B(n_949),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_983),
.A2(n_994),
.B1(n_988),
.B2(n_1140),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1151),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_995),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1029),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_983),
.A2(n_699),
.B1(n_736),
.B2(n_693),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1106),
.B(n_970),
.Y(n_1416)
);

OAI22x1_ASAP7_75t_SL g1417 ( 
.A1(n_997),
.A2(n_607),
.B1(n_610),
.B2(n_597),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1151),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1102),
.B(n_1147),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_997),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1125),
.B(n_688),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1025),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1334),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1151),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1020),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1102),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1283),
.B(n_527),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1034),
.Y(n_1428)
);

NOR2x1_ASAP7_75t_L g1429 ( 
.A(n_1323),
.B(n_758),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1147),
.Y(n_1430)
);

CKINVDCx6p67_ASAP7_75t_R g1431 ( 
.A(n_1049),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1336),
.B(n_527),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1230),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_973),
.A2(n_692),
.B(n_691),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1230),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1000),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_988),
.A2(n_610),
.B1(n_749),
.B2(n_607),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1348),
.B(n_529),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_974),
.A2(n_698),
.B(n_697),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1034),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1230),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1026),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1027),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1043),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1334),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1230),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1289),
.B(n_529),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1309),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1138),
.B(n_706),
.Y(n_1449)
);

OAI22x1_ASAP7_75t_R g1450 ( 
.A1(n_1028),
.A2(n_749),
.B1(n_866),
.B2(n_865),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1246),
.Y(n_1451)
);

AOI22x1_ASAP7_75t_SL g1452 ( 
.A1(n_1028),
.A2(n_866),
.B1(n_870),
.B2(n_865),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1043),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1030),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1031),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1033),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1051),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1290),
.B(n_534),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1036),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1001),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1038),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1051),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1298),
.B(n_534),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1146),
.B(n_717),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1039),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1246),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1323),
.Y(n_1467)
);

OAI22x1_ASAP7_75t_L g1468 ( 
.A1(n_984),
.A2(n_871),
.B1(n_874),
.B2(n_870),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1339),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1339),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_975),
.A2(n_729),
.B(n_718),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1041),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1042),
.Y(n_1473)
);

BUFx8_ASAP7_75t_SL g1474 ( 
.A(n_1040),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1318),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1324),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1044),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1045),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1046),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1335),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1202),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1047),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1048),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1050),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1053),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1053),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1181),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1064),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_976),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1342),
.B(n_730),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1064),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_977),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1016),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1302),
.B(n_540),
.Y(n_1494)
);

INVx5_ASAP7_75t_L g1495 ( 
.A(n_1284),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1182),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1304),
.B(n_540),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1185),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_982),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_985),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1037),
.B(n_542),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_986),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1022),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1099),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_SL g1505 ( 
.A1(n_994),
.A2(n_862),
.B1(n_894),
.B2(n_765),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_989),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1254),
.B(n_738),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1352),
.B(n_542),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1319),
.B(n_745),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1186),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_992),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_993),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1278),
.B(n_757),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1006),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1022),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1032),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1307),
.B(n_543),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_996),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1006),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1284),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_998),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1202),
.Y(n_1523)
);

CKINVDCx11_ASAP7_75t_R g1524 ( 
.A(n_1040),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1004),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_999),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1099),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1321),
.B(n_763),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1144),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1032),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1253),
.A2(n_767),
.B(n_766),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1144),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1196),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1066),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1196),
.Y(n_1535)
);

OAI22x1_ASAP7_75t_L g1536 ( 
.A1(n_990),
.A2(n_874),
.B1(n_877),
.B2(n_871),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1322),
.B(n_772),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1187),
.B(n_543),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1221),
.Y(n_1539)
);

INVx5_ASAP7_75t_L g1540 ( 
.A(n_1284),
.Y(n_1540)
);

INVx5_ASAP7_75t_L g1541 ( 
.A(n_1221),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1005),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1188),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1235),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1235),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1236),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1236),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1277),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1066),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1277),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1255),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1068),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1257),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1258),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1057),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1011),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1259),
.Y(n_1557)
);

BUFx8_ASAP7_75t_L g1558 ( 
.A(n_1244),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1260),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1261),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1264),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1191),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1037),
.B(n_545),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1193),
.Y(n_1564)
);

OAI22x1_ASAP7_75t_SL g1565 ( 
.A1(n_1057),
.A2(n_883),
.B1(n_885),
.B2(n_877),
.Y(n_1565)
);

OAI22x1_ASAP7_75t_R g1566 ( 
.A1(n_1061),
.A2(n_885),
.B1(n_888),
.B2(n_883),
.Y(n_1566)
);

AND2x6_ASAP7_75t_L g1567 ( 
.A(n_1266),
.B(n_726),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1326),
.B(n_777),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1068),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1073),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1013),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1073),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1272),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1268),
.A2(n_764),
.B(n_762),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1273),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1195),
.B(n_545),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1197),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1270),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1271),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1086),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1327),
.B(n_782),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1086),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1199),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1201),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1206),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1274),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1207),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1279),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1320),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1140),
.B(n_549),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1090),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1212),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1214),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1281),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1215),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1328),
.B(n_794),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1217),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1218),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1285),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1223),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1224),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1286),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1329),
.B(n_795),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1090),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1228),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1347),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1153),
.Y(n_1607)
);

BUFx8_ASAP7_75t_SL g1608 ( 
.A(n_1061),
.Y(n_1608)
);

AND2x6_ASAP7_75t_L g1609 ( 
.A(n_1229),
.B(n_755),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1287),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1330),
.B(n_1332),
.Y(n_1611)
);

AND2x6_ASAP7_75t_L g1612 ( 
.A(n_1231),
.B(n_860),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1153),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1337),
.B(n_804),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1232),
.Y(n_1615)
);

BUFx8_ASAP7_75t_L g1616 ( 
.A(n_1216),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1234),
.B(n_549),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1288),
.Y(n_1618)
);

OAI22x1_ASAP7_75t_SL g1619 ( 
.A1(n_1085),
.A2(n_892),
.B1(n_899),
.B2(n_888),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1156),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1291),
.Y(n_1621)
);

AOI22x1_ASAP7_75t_SL g1622 ( 
.A1(n_1085),
.A2(n_899),
.B1(n_900),
.B2(n_892),
.Y(n_1622)
);

BUFx8_ASAP7_75t_SL g1623 ( 
.A(n_1107),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1237),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1293),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1239),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1240),
.Y(n_1627)
);

INVxp33_ASAP7_75t_SL g1628 ( 
.A(n_1156),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1165),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1294),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1169),
.B(n_554),
.Y(n_1631)
);

BUFx12f_ASAP7_75t_L g1632 ( 
.A(n_1165),
.Y(n_1632)
);

INVx6_ASAP7_75t_L g1633 ( 
.A(n_1084),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1241),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1295),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1169),
.B(n_554),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1245),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1250),
.Y(n_1638)
);

INVx5_ASAP7_75t_L g1639 ( 
.A(n_1216),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1251),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1063),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1296),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1275),
.B(n_557),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1183),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1301),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1252),
.Y(n_1646)
);

INVx4_ASAP7_75t_L g1647 ( 
.A(n_1183),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1317),
.B(n_557),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1303),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1347),
.Y(n_1650)
);

BUFx8_ASAP7_75t_L g1651 ( 
.A(n_1333),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1306),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1052),
.Y(n_1653)
);

BUFx8_ASAP7_75t_SL g1654 ( 
.A(n_1107),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1198),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1198),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1054),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1179),
.B(n_558),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1308),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1213),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1056),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1338),
.A2(n_807),
.B(n_806),
.Y(n_1662)
);

BUFx8_ASAP7_75t_SL g1663 ( 
.A(n_1119),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1067),
.B(n_558),
.Y(n_1664)
);

INVx4_ASAP7_75t_L g1665 ( 
.A(n_1213),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1222),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1058),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1222),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1059),
.Y(n_1669)
);

AND2x6_ASAP7_75t_L g1670 ( 
.A(n_1341),
.B(n_938),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1343),
.A2(n_813),
.B(n_809),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1310),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1060),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1062),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1069),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1344),
.A2(n_827),
.B(n_825),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1119),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1226),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1333),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1072),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1345),
.B(n_828),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1675),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1468),
.B(n_900),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_SL g1684 ( 
.A(n_1369),
.B(n_922),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1360),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1524),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1356),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1356),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1399),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1382),
.B(n_1189),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1360),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1364),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1487),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1360),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1364),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1501),
.B(n_1282),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1399),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1419),
.B(n_1373),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1364),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1496),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1498),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1406),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1543),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1562),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1360),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1564),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1501),
.B(n_1351),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1577),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1584),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1419),
.B(n_1075),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1587),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1515),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1592),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1595),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1563),
.B(n_1353),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_SL g1717 ( 
.A(n_1591),
.B(n_934),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1415),
.A2(n_1132),
.B1(n_1159),
.B2(n_1126),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1563),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1373),
.B(n_1076),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1597),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1631),
.B(n_1282),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1626),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1631),
.B(n_1299),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1611),
.B(n_1010),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1409),
.B(n_1299),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1364),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1636),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1634),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1406),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1425),
.Y(n_1731)
);

CKINVDCx16_ASAP7_75t_R g1732 ( 
.A(n_1359),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1638),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1370),
.B(n_1226),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1409),
.B(n_1514),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1409),
.B(n_1514),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1425),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1514),
.B(n_1340),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1646),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1489),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1372),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1489),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1428),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1428),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1492),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1379),
.A2(n_1078),
.B(n_1077),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1440),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1492),
.Y(n_1748)
);

AND2x6_ASAP7_75t_L g1749 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1440),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1444),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1444),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1499),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1372),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1499),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1500),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1453),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1432),
.B(n_1340),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1500),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1502),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1453),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1370),
.B(n_1247),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1474),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1636),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1502),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1506),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1432),
.B(n_1070),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1374),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1467),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1457),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1506),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1643),
.B(n_1088),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1457),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1462),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1462),
.Y(n_1775)
);

CKINVDCx6p67_ASAP7_75t_R g1776 ( 
.A(n_1404),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1420),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1539),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1474),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1420),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1379),
.A2(n_1080),
.B(n_1079),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1539),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1643),
.B(n_1115),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1511),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1432),
.B(n_972),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1539),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1539),
.Y(n_1787)
);

OAI21x1_ASAP7_75t_L g1788 ( 
.A1(n_1434),
.A2(n_1007),
.B(n_1311),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1590),
.Y(n_1789)
);

XOR2xp5_ASAP7_75t_L g1790 ( 
.A(n_1555),
.B(n_1677),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1372),
.Y(n_1791)
);

BUFx8_ASAP7_75t_L g1792 ( 
.A(n_1366),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1539),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1550),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1372),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1438),
.B(n_1247),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1438),
.B(n_1265),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1511),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1522),
.Y(n_1799)
);

XNOR2xp5_ASAP7_75t_L g1800 ( 
.A(n_1505),
.B(n_1126),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1550),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1522),
.Y(n_1802)
);

INVx5_ASAP7_75t_L g1803 ( 
.A(n_1360),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1384),
.B(n_1300),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1374),
.B(n_1083),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1526),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1363),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1447),
.B(n_1265),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1447),
.B(n_1267),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1526),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1436),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1436),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1363),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1524),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1460),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1363),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1463),
.B(n_1497),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1460),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1525),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1463),
.B(n_1267),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1438),
.B(n_1354),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1371),
.B(n_1388),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1525),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1508),
.B(n_1354),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1375),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1391),
.B(n_1087),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1497),
.B(n_1003),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1542),
.Y(n_1828)
);

INVx5_ASAP7_75t_L g1829 ( 
.A(n_1363),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1508),
.B(n_1346),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1355),
.B(n_1386),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1550),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1355),
.B(n_1275),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1508),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1542),
.Y(n_1835)
);

AND2x2_ASAP7_75t_SL g1836 ( 
.A(n_1574),
.B(n_1405),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1550),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1507),
.B(n_1010),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1375),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1556),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1556),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1571),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1371),
.B(n_1388),
.Y(n_1843)
);

BUFx12f_ASAP7_75t_L g1844 ( 
.A(n_1606),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1375),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1633),
.A2(n_1120),
.B1(n_1123),
.B2(n_1019),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1371),
.B(n_833),
.Y(n_1847)
);

CKINVDCx14_ASAP7_75t_R g1848 ( 
.A(n_1515),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1388),
.B(n_834),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1664),
.Y(n_1850)
);

AND2x6_ASAP7_75t_L g1851 ( 
.A(n_1386),
.B(n_1091),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1391),
.B(n_1094),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1550),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1571),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1381),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1427),
.B(n_842),
.Y(n_1856)
);

AND3x2_ASAP7_75t_L g1857 ( 
.A(n_1520),
.B(n_1092),
.C(n_1065),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1608),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1363),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1465),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1512),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1465),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1512),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1477),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1426),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1512),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1458),
.B(n_843),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1381),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1381),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1451),
.Y(n_1870)
);

NAND2x1_ASAP7_75t_L g1871 ( 
.A(n_1392),
.B(n_1407),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1519),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1520),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1519),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1519),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1585),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1572),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1494),
.B(n_846),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1381),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1585),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1477),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1600),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1600),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1624),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1624),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1478),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1667),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1509),
.B(n_853),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1528),
.B(n_574),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1537),
.B(n_574),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1410),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1451),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1478),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1667),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1479),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1667),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1410),
.B(n_1003),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1572),
.Y(n_1898)
);

INVxp33_ASAP7_75t_SL g1899 ( 
.A(n_1411),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1667),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1658),
.B(n_1093),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1674),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1633),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1479),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1674),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1389),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1426),
.B(n_1096),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1430),
.B(n_1097),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1485),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1674),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1467),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1451),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1481),
.B(n_1679),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1674),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1389),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1389),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1362),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1367),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1377),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1608),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1633),
.A2(n_1513),
.B1(n_1376),
.B2(n_1414),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1607),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1607),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1400),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1380),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1476),
.B(n_947),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1467),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1485),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1383),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1485),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1568),
.B(n_581),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1402),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1400),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1581),
.B(n_581),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1485),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1422),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1486),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1430),
.B(n_1098),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1442),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1481),
.B(n_1012),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1443),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1393),
.B(n_1104),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1486),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1400),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1393),
.B(n_1105),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1454),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1400),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1390),
.B(n_1108),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1486),
.Y(n_1949)
);

BUFx8_ASAP7_75t_L g1950 ( 
.A(n_1366),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1455),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1451),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1486),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1596),
.B(n_582),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1658),
.B(n_1103),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1623),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1418),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1660),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1456),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1633),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1418),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1467),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1603),
.B(n_1019),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1459),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1461),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1660),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1451),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1418),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1538),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1614),
.B(n_582),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1418),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1472),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1483),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1424),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1484),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1488),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1681),
.B(n_1120),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1551),
.B(n_1012),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1488),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1658),
.B(n_1639),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1659),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1680),
.B(n_1109),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1488),
.Y(n_1983)
);

AND2x6_ASAP7_75t_L g1984 ( 
.A(n_1538),
.B(n_1110),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1488),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1659),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1639),
.B(n_1114),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1672),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1672),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1551),
.B(n_1312),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1513),
.B(n_1123),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1641),
.B(n_1150),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1678),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1424),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1424),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1491),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1583),
.Y(n_1997)
);

BUFx12f_ASAP7_75t_L g1998 ( 
.A(n_1606),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1491),
.Y(n_1999)
);

BUFx8_ASAP7_75t_L g2000 ( 
.A(n_1395),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1583),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1424),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1491),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1593),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1593),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1598),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1392),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1433),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1433),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1598),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1491),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1601),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1601),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1605),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1605),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1553),
.B(n_1315),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1504),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1504),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1361),
.B(n_590),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1538),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1416),
.B(n_590),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1553),
.B(n_1316),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1615),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1680),
.B(n_1518),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1433),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1615),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1433),
.Y(n_2027)
);

CKINVDCx6p67_ASAP7_75t_R g2028 ( 
.A(n_1404),
.Y(n_2028)
);

CKINVDCx20_ASAP7_75t_R g2029 ( 
.A(n_1555),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1627),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1435),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1627),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1677),
.Y(n_2033)
);

CKINVDCx16_ASAP7_75t_R g2034 ( 
.A(n_1395),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1504),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1557),
.B(n_1135),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1680),
.B(n_1111),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1421),
.B(n_592),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1637),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1434),
.A2(n_1113),
.B(n_1112),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1637),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_SL g2042 ( 
.A1(n_1628),
.A2(n_1132),
.B1(n_1167),
.B2(n_1159),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1523),
.B(n_1157),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1639),
.B(n_1117),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1639),
.B(n_1210),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1640),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1640),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1504),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1435),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1473),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1531),
.A2(n_1118),
.B(n_1116),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1527),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1473),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1435),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1527),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1435),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1473),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1527),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1518),
.B(n_1121),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1473),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1527),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1482),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1532),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1441),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1441),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1441),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1441),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1523),
.B(n_1175),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1449),
.B(n_1150),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1518),
.B(n_1122),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1532),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1482),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1482),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_1623),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1464),
.B(n_592),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1687),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1732),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_1940),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1817),
.B(n_1408),
.Y(n_2079)
);

BUFx4f_ASAP7_75t_L g2080 ( 
.A(n_1776),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1682),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1687),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1942),
.Y(n_2083)
);

BUFx3_ASAP7_75t_L g2084 ( 
.A(n_1698),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1693),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1735),
.B(n_1490),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1736),
.B(n_1405),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_1942),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1700),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1850),
.B(n_1725),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1701),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1942),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1978),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1836),
.A2(n_1405),
.B1(n_1670),
.B2(n_1612),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1831),
.B(n_1358),
.Y(n_2095)
);

NOR3xp33_ASAP7_75t_L g2096 ( 
.A(n_1725),
.B(n_1678),
.C(n_1445),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1702),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1688),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1704),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1705),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1833),
.B(n_1679),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1945),
.Y(n_2102)
);

INVx2_ASAP7_75t_SL g2103 ( 
.A(n_1978),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1707),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1709),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1688),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1689),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1843),
.B(n_1408),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1763),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_L g2110 ( 
.A(n_1984),
.B(n_1670),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1710),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1712),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1714),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1836),
.B(n_1448),
.Y(n_2114)
);

AND2x6_ASAP7_75t_L g2115 ( 
.A(n_1945),
.B(n_1696),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1689),
.Y(n_2116)
);

INVx4_ASAP7_75t_L g2117 ( 
.A(n_1769),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1715),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1697),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1721),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1738),
.B(n_1358),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1723),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_1734),
.A2(n_1471),
.B(n_1439),
.Y(n_2123)
);

AND2x6_ASAP7_75t_L g2124 ( 
.A(n_1945),
.B(n_1648),
.Y(n_2124)
);

INVx4_ASAP7_75t_L g2125 ( 
.A(n_1769),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1697),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1703),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_1897),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1991),
.B(n_1448),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_L g2130 ( 
.A(n_1984),
.B(n_1670),
.Y(n_2130)
);

INVx4_ASAP7_75t_SL g2131 ( 
.A(n_1984),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1838),
.B(n_1358),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1838),
.B(n_1403),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1991),
.B(n_1589),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1698),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1729),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1733),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1703),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_1877),
.Y(n_2139)
);

BUFx10_ASAP7_75t_L g2140 ( 
.A(n_1992),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1711),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1730),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1690),
.B(n_1403),
.Y(n_2143)
);

AOI22x1_ASAP7_75t_L g2144 ( 
.A1(n_1834),
.A2(n_1468),
.B1(n_1536),
.B2(n_1665),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1739),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1789),
.B(n_1591),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_2007),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1730),
.Y(n_2148)
);

OAI21xp33_ASAP7_75t_SL g2149 ( 
.A1(n_1822),
.A2(n_1471),
.B(n_1439),
.Y(n_2149)
);

AND3x1_ASAP7_75t_L g2150 ( 
.A(n_1684),
.B(n_1172),
.C(n_1394),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1769),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2024),
.B(n_1589),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1758),
.B(n_1403),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1731),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1731),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1833),
.B(n_1591),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1827),
.B(n_1613),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1737),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_L g2159 ( 
.A(n_1984),
.B(n_1670),
.Y(n_2159)
);

INVx5_ASAP7_75t_L g2160 ( 
.A(n_1984),
.Y(n_2160)
);

NAND2xp33_ASAP7_75t_L g2161 ( 
.A(n_1851),
.B(n_1670),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1698),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1990),
.Y(n_2163)
);

CKINVDCx20_ASAP7_75t_R g2164 ( 
.A(n_1777),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_SL g2165 ( 
.A(n_1720),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1737),
.Y(n_2166)
);

AO21x2_ASAP7_75t_L g2167 ( 
.A1(n_1734),
.A2(n_1671),
.B(n_1662),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1743),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1711),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2069),
.B(n_1574),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_2024),
.B(n_1613),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1743),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1990),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1744),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2016),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2024),
.B(n_1613),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1744),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2016),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_1768),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1747),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2022),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1768),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2022),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2069),
.B(n_1574),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_1822),
.A2(n_1670),
.B1(n_1612),
.B2(n_1609),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_2007),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2043),
.B(n_1647),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1747),
.Y(n_2188)
);

AND3x2_ASAP7_75t_L g2189 ( 
.A(n_1717),
.B(n_1445),
.C(n_1423),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_L g2190 ( 
.A(n_1851),
.B(n_1609),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1997),
.Y(n_2191)
);

INVx6_ASAP7_75t_L g2192 ( 
.A(n_1792),
.Y(n_2192)
);

INVxp33_ASAP7_75t_L g2193 ( 
.A(n_1804),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2001),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_1711),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1963),
.B(n_1647),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1750),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2004),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_1719),
.B(n_1423),
.Y(n_2199)
);

INVx2_ASAP7_75t_SL g2200 ( 
.A(n_1720),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1963),
.B(n_1647),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1977),
.B(n_1665),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2005),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1750),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1751),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2006),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2010),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_1962),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1977),
.B(n_1476),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2068),
.B(n_1665),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1921),
.B(n_1476),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_1720),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2012),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1751),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_L g2215 ( 
.A(n_1851),
.B(n_1609),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1752),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1746),
.A2(n_1612),
.B1(n_1609),
.B2(n_1567),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_1805),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2013),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_1692),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1752),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2014),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1757),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1757),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_1805),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2015),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1772),
.B(n_1576),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1761),
.Y(n_2228)
);

INVx6_ASAP7_75t_L g2229 ( 
.A(n_1792),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2023),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_R g2231 ( 
.A(n_1848),
.B(n_1666),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1783),
.B(n_1576),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1761),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1770),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1962),
.Y(n_2235)
);

INVx2_ASAP7_75t_SL g2236 ( 
.A(n_1805),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1770),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_1719),
.B(n_1469),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1773),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_1762),
.B(n_1628),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_L g2241 ( 
.A(n_1762),
.B(n_1666),
.C(n_1503),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2026),
.Y(n_2242)
);

NAND2xp33_ASAP7_75t_L g2243 ( 
.A(n_1851),
.B(n_1609),
.Y(n_2243)
);

NOR2x1p5_ASAP7_75t_L g2244 ( 
.A(n_1776),
.B(n_1431),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1773),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_1982),
.Y(n_2246)
);

NAND2x1p5_ASAP7_75t_L g2247 ( 
.A(n_1746),
.B(n_1639),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_R g2248 ( 
.A(n_1848),
.B(n_1650),
.Y(n_2248)
);

BUFx10_ASAP7_75t_L g2249 ( 
.A(n_1992),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1774),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1774),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1775),
.Y(n_2252)
);

BUFx3_ASAP7_75t_L g2253 ( 
.A(n_1826),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2030),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2032),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1834),
.B(n_1576),
.Y(n_2256)
);

NAND2xp33_ASAP7_75t_L g2257 ( 
.A(n_1851),
.B(n_1609),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1775),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2039),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_1728),
.B(n_1493),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1982),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1692),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2041),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1763),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1860),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2046),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1860),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1913),
.B(n_1617),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1862),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1862),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1692),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_R g2272 ( 
.A(n_1779),
.B(n_1650),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1864),
.Y(n_2273)
);

INVx2_ASAP7_75t_SL g2274 ( 
.A(n_1826),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1808),
.B(n_1809),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1864),
.Y(n_2276)
);

OR2x6_ASAP7_75t_L g2277 ( 
.A(n_1844),
.B(n_1516),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_SL g2278 ( 
.A1(n_1899),
.A2(n_1612),
.B1(n_1567),
.B2(n_1176),
.Y(n_2278)
);

BUFx3_ASAP7_75t_L g2279 ( 
.A(n_1826),
.Y(n_2279)
);

INVxp33_ASAP7_75t_L g2280 ( 
.A(n_2042),
.Y(n_2280)
);

AO22x2_ASAP7_75t_L g2281 ( 
.A1(n_1846),
.A2(n_1452),
.B1(n_1622),
.B2(n_1437),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1708),
.B(n_1617),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1728),
.B(n_1517),
.Y(n_2283)
);

AND3x2_ASAP7_75t_L g2284 ( 
.A(n_1898),
.B(n_1470),
.C(n_1469),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_1820),
.B(n_1722),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2047),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1708),
.B(n_1617),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1982),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1881),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1779),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1881),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2037),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_1852),
.Y(n_2293)
);

BUFx10_ASAP7_75t_L g2294 ( 
.A(n_1857),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_1767),
.B(n_1662),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1886),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1886),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1796),
.B(n_1671),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_L g2299 ( 
.A(n_1969),
.B(n_2020),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1692),
.Y(n_2300)
);

AOI21x1_ASAP7_75t_L g2301 ( 
.A1(n_1861),
.A2(n_1866),
.B(n_1863),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_1764),
.B(n_1530),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1893),
.Y(n_2303)
);

INVx4_ASAP7_75t_L g2304 ( 
.A(n_1911),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2037),
.Y(n_2305)
);

NAND2xp33_ASAP7_75t_R g2306 ( 
.A(n_1899),
.B(n_1470),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_1852),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_1764),
.B(n_1549),
.Y(n_2308)
);

INVx5_ASAP7_75t_L g2309 ( 
.A(n_1695),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_1695),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1716),
.B(n_1648),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_1797),
.B(n_1676),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1785),
.B(n_1569),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_1821),
.B(n_1570),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2037),
.Y(n_2315)
);

INVxp33_ASAP7_75t_L g2316 ( 
.A(n_1790),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_1852),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_1907),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1876),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_SL g2320 ( 
.A1(n_1718),
.A2(n_1612),
.B1(n_1567),
.B2(n_1176),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1880),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1893),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_1871),
.Y(n_2323)
);

INVxp67_ASAP7_75t_SL g2324 ( 
.A(n_1903),
.Y(n_2324)
);

OAI21xp33_ASAP7_75t_SL g2325 ( 
.A1(n_1716),
.A2(n_1676),
.B(n_1531),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1888),
.B(n_1648),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2019),
.B(n_1612),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_1969),
.A2(n_1604),
.B1(n_1620),
.B2(n_1582),
.Y(n_2328)
);

INVx6_ASAP7_75t_L g2329 ( 
.A(n_1792),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_1824),
.B(n_1655),
.Y(n_2330)
);

INVxp33_ASAP7_75t_SL g2331 ( 
.A(n_1800),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_1858),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1882),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_1922),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2021),
.B(n_1567),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1895),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_1923),
.B(n_1178),
.C(n_1167),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1724),
.B(n_1629),
.Y(n_2338)
);

NAND2xp33_ASAP7_75t_L g2339 ( 
.A(n_2020),
.B(n_1567),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1883),
.Y(n_2340)
);

INVxp67_ASAP7_75t_SL g2341 ( 
.A(n_1903),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1695),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_1966),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1884),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_1695),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1895),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1726),
.B(n_1668),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_1858),
.Y(n_2348)
);

NAND2xp33_ASAP7_75t_SL g2349 ( 
.A(n_1830),
.B(n_1536),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1872),
.B(n_1644),
.Y(n_2350)
);

INVx5_ASAP7_75t_L g2351 ( 
.A(n_1699),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1885),
.Y(n_2352)
);

INVx3_ASAP7_75t_L g2353 ( 
.A(n_1968),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_1891),
.B(n_1184),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1907),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_1874),
.B(n_1875),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1907),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_1780),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1908),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2038),
.B(n_1567),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1908),
.Y(n_2361)
);

INVx2_ASAP7_75t_SL g2362 ( 
.A(n_1908),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1938),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1904),
.Y(n_2364)
);

AOI22xp33_ASAP7_75t_L g2365 ( 
.A1(n_1746),
.A2(n_1174),
.B1(n_1220),
.B2(n_958),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1904),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_1847),
.A2(n_1849),
.B1(n_1891),
.B2(n_2075),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2059),
.B(n_1475),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1740),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1856),
.B(n_1559),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_1781),
.A2(n_1683),
.B1(n_2051),
.B2(n_2059),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1742),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1745),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_1960),
.B(n_1889),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1867),
.B(n_1559),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1938),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1748),
.Y(n_2377)
);

INVx4_ASAP7_75t_L g2378 ( 
.A(n_1911),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1699),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1938),
.Y(n_2380)
);

AND2x6_ASAP7_75t_L g2381 ( 
.A(n_1926),
.B(n_1124),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1753),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_1780),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1917),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1878),
.B(n_1559),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1918),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1755),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1919),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1925),
.Y(n_2389)
);

AND2x6_ASAP7_75t_L g2390 ( 
.A(n_2059),
.B(n_1127),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_2029),
.Y(n_2391)
);

OAI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_1890),
.A2(n_1431),
.B1(n_1534),
.B2(n_1516),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_1960),
.B(n_1184),
.Y(n_2393)
);

INVx2_ASAP7_75t_SL g2394 ( 
.A(n_2036),
.Y(n_2394)
);

INVx2_ASAP7_75t_SL g2395 ( 
.A(n_2036),
.Y(n_2395)
);

AOI21x1_ASAP7_75t_L g2396 ( 
.A1(n_1756),
.A2(n_1544),
.B(n_1535),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2070),
.B(n_1475),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_1958),
.B(n_1233),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1931),
.B(n_1554),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_1981),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_1934),
.B(n_1554),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1929),
.Y(n_2402)
);

NAND3xp33_ASAP7_75t_L g2403 ( 
.A(n_1683),
.B(n_1024),
.C(n_1200),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_1968),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1932),
.Y(n_2405)
);

AND2x2_ASAP7_75t_SL g2406 ( 
.A(n_2051),
.B(n_1781),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_1954),
.B(n_1194),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_2070),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_1920),
.Y(n_2409)
);

BUFx8_ASAP7_75t_SL g2410 ( 
.A(n_1920),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_1699),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1759),
.Y(n_2412)
);

INVx2_ASAP7_75t_SL g2413 ( 
.A(n_2070),
.Y(n_2413)
);

AND3x2_ASAP7_75t_L g2414 ( 
.A(n_1713),
.B(n_1280),
.C(n_1203),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_1699),
.Y(n_2415)
);

OAI22xp33_ASAP7_75t_L g2416 ( 
.A1(n_1970),
.A2(n_1534),
.B1(n_1580),
.B2(n_1552),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1760),
.Y(n_2417)
);

BUFx10_ASAP7_75t_L g2418 ( 
.A(n_1749),
.Y(n_2418)
);

INVx6_ASAP7_75t_L g2419 ( 
.A(n_1950),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1765),
.Y(n_2420)
);

CKINVDCx20_ASAP7_75t_R g2421 ( 
.A(n_2029),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1766),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_1771),
.Y(n_2423)
);

AND3x2_ASAP7_75t_L g2424 ( 
.A(n_1873),
.B(n_1227),
.C(n_1101),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1784),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_1798),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_1993),
.B(n_1948),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_1799),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1936),
.B(n_1554),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_1802),
.Y(n_2430)
);

INVx4_ASAP7_75t_L g2431 ( 
.A(n_1911),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_L g2432 ( 
.A(n_1901),
.B(n_1651),
.C(n_1616),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_1727),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1806),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1939),
.B(n_1554),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1941),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_1948),
.B(n_1986),
.Y(n_2437)
);

INVx4_ASAP7_75t_L g2438 ( 
.A(n_1927),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2028),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1810),
.Y(n_2440)
);

AND2x2_ASAP7_75t_SL g2441 ( 
.A(n_2051),
.B(n_1238),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2028),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1946),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1951),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1959),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1964),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_1988),
.Y(n_2447)
);

INVx2_ASAP7_75t_SL g2448 ( 
.A(n_1989),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1909),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1965),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_1980),
.B(n_1480),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1972),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1973),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_1948),
.B(n_1305),
.Y(n_2454)
);

INVx2_ASAP7_75t_SL g2455 ( 
.A(n_1811),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_1909),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_1928),
.Y(n_2457)
);

CKINVDCx6p67_ASAP7_75t_R g2458 ( 
.A(n_1844),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1975),
.B(n_1554),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_1980),
.B(n_1480),
.Y(n_2460)
);

AND2x6_ASAP7_75t_L g2461 ( 
.A(n_1812),
.B(n_1128),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1815),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_1818),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_1819),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1823),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_1928),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1930),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1887),
.B(n_1894),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2033),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_1930),
.Y(n_2470)
);

BUFx10_ASAP7_75t_L g2471 ( 
.A(n_1749),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1828),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1835),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_1968),
.Y(n_2474)
);

AND2x4_ASAP7_75t_L g2475 ( 
.A(n_1840),
.B(n_1653),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_1781),
.A2(n_1205),
.B1(n_1208),
.B2(n_1194),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1841),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2033),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_1842),
.Y(n_2479)
);

AND2x6_ASAP7_75t_L g2480 ( 
.A(n_1854),
.B(n_1130),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_1865),
.B(n_1205),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_1935),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_1935),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2265),
.Y(n_2484)
);

OAI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_2090),
.A2(n_1955),
.B1(n_1901),
.B2(n_1219),
.Y(n_2485)
);

INVx2_ASAP7_75t_SL g2486 ( 
.A(n_2139),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2265),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2267),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2267),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2083),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2334),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2090),
.B(n_2196),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2086),
.B(n_1749),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2083),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2269),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2083),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2343),
.Y(n_2497)
);

INVx4_ASAP7_75t_L g2498 ( 
.A(n_2083),
.Y(n_2498)
);

INVx4_ASAP7_75t_L g2499 ( 
.A(n_2102),
.Y(n_2499)
);

OAI22xp33_ASAP7_75t_SL g2500 ( 
.A1(n_2211),
.A2(n_1955),
.B1(n_1211),
.B2(n_1248),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2102),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2094),
.A2(n_2040),
.B1(n_1211),
.B2(n_1248),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2076),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2102),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2076),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2269),
.Y(n_2506)
);

AND2x6_ASAP7_75t_L g2507 ( 
.A(n_2102),
.B(n_1778),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2082),
.Y(n_2508)
);

INVx1_ASAP7_75t_SL g2509 ( 
.A(n_2199),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2238),
.B(n_1686),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2270),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_2358),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2082),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2179),
.B(n_2182),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2394),
.B(n_1987),
.Y(n_2515)
);

HB1xp67_ASAP7_75t_L g2516 ( 
.A(n_2395),
.Y(n_2516)
);

OAI221xp5_ASAP7_75t_L g2517 ( 
.A1(n_2196),
.A2(n_914),
.B1(n_915),
.B2(n_913),
.C(n_906),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2094),
.A2(n_2040),
.B1(n_1256),
.B2(n_1263),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2326),
.B(n_1749),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_2088),
.Y(n_2520)
);

AND2x2_ASAP7_75t_SL g2521 ( 
.A(n_2150),
.B(n_2034),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2147),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2201),
.B(n_1208),
.Y(n_2523)
);

AND2x4_ASAP7_75t_L g2524 ( 
.A(n_2179),
.B(n_2182),
.Y(n_2524)
);

OR2x6_ASAP7_75t_L g2525 ( 
.A(n_2192),
.B(n_1998),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2201),
.B(n_1256),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2202),
.B(n_1263),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2308),
.B(n_1814),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2270),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2253),
.B(n_1987),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2202),
.B(n_1269),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2273),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2273),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2170),
.B(n_1749),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2383),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2184),
.B(n_1778),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2098),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2276),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2276),
.Y(n_2539)
);

INVx4_ASAP7_75t_L g2540 ( 
.A(n_2084),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2187),
.B(n_2210),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2289),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2253),
.B(n_2044),
.Y(n_2543)
);

AND2x4_ASAP7_75t_L g2544 ( 
.A(n_2279),
.B(n_2044),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2291),
.Y(n_2545)
);

INVx4_ASAP7_75t_L g2546 ( 
.A(n_2084),
.Y(n_2546)
);

INVx1_ASAP7_75t_SL g2547 ( 
.A(n_2157),
.Y(n_2547)
);

AO22x2_ASAP7_75t_L g2548 ( 
.A1(n_2211),
.A2(n_1566),
.B1(n_1450),
.B2(n_1956),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2291),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2106),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2374),
.B(n_2132),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2296),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2101),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2106),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2296),
.Y(n_2555)
);

INVxp67_ASAP7_75t_SL g2556 ( 
.A(n_2088),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2107),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2297),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2297),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2303),
.Y(n_2560)
);

OAI21xp33_ASAP7_75t_L g2561 ( 
.A1(n_2311),
.A2(n_1297),
.B(n_1269),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2147),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2279),
.B(n_2045),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2303),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2322),
.Y(n_2565)
);

CKINVDCx16_ASAP7_75t_R g2566 ( 
.A(n_2248),
.Y(n_2566)
);

AND2x4_ASAP7_75t_L g2567 ( 
.A(n_2293),
.B(n_2045),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2322),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2107),
.Y(n_2569)
);

AND2x6_ASAP7_75t_L g2570 ( 
.A(n_2092),
.B(n_1782),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2116),
.Y(n_2571)
);

AND3x1_ASAP7_75t_L g2572 ( 
.A(n_2096),
.B(n_1565),
.C(n_1417),
.Y(n_2572)
);

AND2x2_ASAP7_75t_SL g2573 ( 
.A(n_2080),
.B(n_1654),
.Y(n_2573)
);

INVx8_ASAP7_75t_L g2574 ( 
.A(n_2390),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2441),
.A2(n_1313),
.B1(n_1297),
.B2(n_913),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2469),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2116),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2119),
.Y(n_2578)
);

AO22x2_ASAP7_75t_L g2579 ( 
.A1(n_2241),
.A2(n_2403),
.B1(n_2337),
.B2(n_2129),
.Y(n_2579)
);

INVx4_ASAP7_75t_L g2580 ( 
.A(n_2135),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2209),
.B(n_1178),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2119),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2336),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2146),
.B(n_1219),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2126),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2156),
.B(n_1552),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2336),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2293),
.B(n_1896),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2135),
.B(n_1900),
.Y(n_2589)
);

AO22x2_ASAP7_75t_L g2590 ( 
.A1(n_2129),
.A2(n_2074),
.B1(n_1262),
.B2(n_1249),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2346),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2146),
.B(n_1225),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2374),
.B(n_1782),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2346),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2364),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2092),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2313),
.B(n_1313),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2093),
.B(n_1580),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2147),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2162),
.B(n_1902),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2162),
.B(n_1905),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2364),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2366),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2126),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2147),
.Y(n_2605)
);

BUFx3_ASAP7_75t_L g2606 ( 
.A(n_2077),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2366),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2407),
.B(n_1632),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2127),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2246),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2441),
.A2(n_914),
.B1(n_915),
.B2(n_906),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_SL g2612 ( 
.A(n_2407),
.B(n_1632),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2127),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2292),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2315),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2193),
.B(n_1225),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2369),
.Y(n_2617)
);

INVxp33_ASAP7_75t_L g2618 ( 
.A(n_2398),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2313),
.B(n_1656),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2408),
.B(n_2413),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2260),
.B(n_1656),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2260),
.B(n_2283),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2231),
.Y(n_2623)
);

INVx4_ASAP7_75t_L g2624 ( 
.A(n_2186),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2103),
.B(n_1401),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2138),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2369),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2133),
.A2(n_1914),
.B1(n_1910),
.B2(n_1937),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2283),
.B(n_1401),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2372),
.Y(n_2630)
);

NOR2xp67_ASAP7_75t_L g2631 ( 
.A(n_2246),
.B(n_2071),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2138),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2372),
.Y(n_2633)
);

INVx4_ASAP7_75t_L g2634 ( 
.A(n_2186),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2373),
.Y(n_2635)
);

AND2x6_ASAP7_75t_L g2636 ( 
.A(n_2087),
.B(n_1786),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2373),
.Y(n_2637)
);

AND2x6_ASAP7_75t_L g2638 ( 
.A(n_2153),
.B(n_1786),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2338),
.B(n_1413),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2193),
.B(n_1242),
.Y(n_2640)
);

INVx4_ASAP7_75t_L g2641 ( 
.A(n_2186),
.Y(n_2641)
);

INVx4_ASAP7_75t_L g2642 ( 
.A(n_2186),
.Y(n_2642)
);

INVx2_ASAP7_75t_SL g2643 ( 
.A(n_2427),
.Y(n_2643)
);

INVx8_ASAP7_75t_L g2644 ( 
.A(n_2390),
.Y(n_2644)
);

BUFx6f_ASAP7_75t_L g2645 ( 
.A(n_2220),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2261),
.Y(n_2646)
);

AND3x4_ASAP7_75t_L g2647 ( 
.A(n_2306),
.B(n_1619),
.C(n_1243),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2391),
.B(n_1242),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2377),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2377),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2227),
.B(n_1616),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_L g2652 ( 
.A(n_2134),
.B(n_1243),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2382),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2382),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2285),
.B(n_1413),
.Y(n_2655)
);

AO22x2_ASAP7_75t_L g2656 ( 
.A1(n_2134),
.A2(n_1314),
.B1(n_1292),
.B2(n_1654),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2387),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2387),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2142),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2412),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_2141),
.B(n_1653),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2232),
.B(n_1616),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2220),
.Y(n_2663)
);

INVx6_ASAP7_75t_L g2664 ( 
.A(n_2192),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2142),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2261),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2288),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_L g2668 ( 
.A(n_2302),
.B(n_2275),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2220),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2412),
.Y(n_2670)
);

INVx8_ASAP7_75t_L g2671 ( 
.A(n_2390),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2314),
.B(n_1292),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2417),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2160),
.B(n_1927),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2417),
.Y(n_2675)
);

INVx2_ASAP7_75t_SL g2676 ( 
.A(n_2078),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2143),
.B(n_1787),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2420),
.Y(n_2678)
);

NAND2x1p5_ASAP7_75t_L g2679 ( 
.A(n_2160),
.B(n_1927),
.Y(n_2679)
);

BUFx2_ASAP7_75t_L g2680 ( 
.A(n_2164),
.Y(n_2680)
);

INVx4_ASAP7_75t_L g2681 ( 
.A(n_2288),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2148),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2420),
.Y(n_2683)
);

BUFx3_ASAP7_75t_L g2684 ( 
.A(n_2164),
.Y(n_2684)
);

NOR2x1p5_ASAP7_75t_L g2685 ( 
.A(n_2458),
.B(n_1998),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2422),
.Y(n_2686)
);

INVxp67_ASAP7_75t_L g2687 ( 
.A(n_2282),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2422),
.Y(n_2688)
);

BUFx2_ASAP7_75t_L g2689 ( 
.A(n_2421),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2169),
.B(n_1657),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2423),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2423),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2195),
.B(n_2200),
.Y(n_2693)
);

INVx3_ASAP7_75t_L g2694 ( 
.A(n_2305),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2421),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_2220),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2121),
.B(n_1787),
.Y(n_2697)
);

OR2x2_ASAP7_75t_L g2698 ( 
.A(n_2478),
.B(n_1657),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2425),
.Y(n_2699)
);

INVx1_ASAP7_75t_SL g2700 ( 
.A(n_2275),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2095),
.B(n_1793),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_L g2702 ( 
.A(n_2240),
.B(n_1365),
.Y(n_2702)
);

AND2x6_ASAP7_75t_L g2703 ( 
.A(n_2327),
.B(n_1793),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2148),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2425),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2426),
.Y(n_2706)
);

NAND3x1_ASAP7_75t_L g2707 ( 
.A(n_2240),
.B(n_1663),
.C(n_1950),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2287),
.B(n_1794),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2426),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2393),
.B(n_1365),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2393),
.B(n_1661),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2305),
.Y(n_2712)
);

BUFx4f_ASAP7_75t_L g2713 ( 
.A(n_2192),
.Y(n_2713)
);

INVxp67_ASAP7_75t_L g2714 ( 
.A(n_2256),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2370),
.B(n_1794),
.Y(n_2715)
);

INVx4_ASAP7_75t_L g2716 ( 
.A(n_2390),
.Y(n_2716)
);

AND2x6_ASAP7_75t_L g2717 ( 
.A(n_2335),
.B(n_1801),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2375),
.B(n_1801),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2212),
.B(n_2218),
.Y(n_2719)
);

OAI22xp5_ASAP7_75t_SL g2720 ( 
.A1(n_2331),
.A2(n_923),
.B1(n_924),
.B2(n_917),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2154),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2428),
.Y(n_2722)
);

INVxp67_ASAP7_75t_SL g2723 ( 
.A(n_2262),
.Y(n_2723)
);

NAND2xp33_ASAP7_75t_SL g2724 ( 
.A(n_2231),
.B(n_594),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2428),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2225),
.B(n_1661),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2154),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2385),
.B(n_1832),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2430),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2128),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2155),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_2262),
.Y(n_2732)
);

OAI22xp33_ASAP7_75t_SL g2733 ( 
.A1(n_2144),
.A2(n_923),
.B1(n_924),
.B2(n_917),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2430),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2155),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2262),
.Y(n_2736)
);

BUFx2_ASAP7_75t_L g2737 ( 
.A(n_2454),
.Y(n_2737)
);

NAND2x1p5_ASAP7_75t_L g2738 ( 
.A(n_2160),
.B(n_1937),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2434),
.Y(n_2739)
);

OR2x2_ASAP7_75t_L g2740 ( 
.A(n_2354),
.B(n_1669),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2354),
.B(n_1669),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2262),
.Y(n_2742)
);

AND2x6_ASAP7_75t_L g2743 ( 
.A(n_2360),
.B(n_1832),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2158),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2115),
.B(n_1837),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2158),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2314),
.B(n_1673),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_2271),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_SL g2749 ( 
.A1(n_2280),
.A2(n_943),
.B1(n_946),
.B2(n_930),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2481),
.B(n_1673),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2481),
.B(n_1652),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2140),
.B(n_1385),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2236),
.B(n_1943),
.Y(n_2753)
);

INVx5_ASAP7_75t_L g2754 ( 
.A(n_2160),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2434),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2163),
.B(n_1652),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2410),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2440),
.Y(n_2758)
);

A2O1A1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2325),
.A2(n_1788),
.B(n_1949),
.C(n_1943),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2440),
.Y(n_2760)
);

INVx2_ASAP7_75t_SL g2761 ( 
.A(n_2475),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2166),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2274),
.B(n_1949),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2307),
.B(n_2317),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2166),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2115),
.B(n_2367),
.Y(n_2766)
);

INVxp67_ASAP7_75t_L g2767 ( 
.A(n_2268),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2140),
.B(n_1385),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2115),
.B(n_1837),
.Y(n_2769)
);

INVxp67_ASAP7_75t_L g2770 ( 
.A(n_2437),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2140),
.B(n_1663),
.Y(n_2771)
);

BUFx3_ASAP7_75t_L g2772 ( 
.A(n_2410),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2168),
.Y(n_2773)
);

BUFx6f_ASAP7_75t_L g2774 ( 
.A(n_2271),
.Y(n_2774)
);

AND2x6_ASAP7_75t_L g2775 ( 
.A(n_2355),
.B(n_1853),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2168),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2172),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2172),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2249),
.B(n_1385),
.Y(n_2779)
);

OAI21xp33_ASAP7_75t_L g2780 ( 
.A1(n_2476),
.A2(n_2365),
.B(n_2175),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2174),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2318),
.B(n_2362),
.Y(n_2782)
);

AND2x6_ASAP7_75t_L g2783 ( 
.A(n_2357),
.B(n_1853),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2115),
.B(n_2124),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2235),
.Y(n_2785)
);

INVx4_ASAP7_75t_SL g2786 ( 
.A(n_2124),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2249),
.B(n_1558),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_SL g2788 ( 
.A1(n_2281),
.A2(n_1558),
.B1(n_1651),
.B2(n_943),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2174),
.Y(n_2789)
);

BUFx3_ASAP7_75t_L g2790 ( 
.A(n_2080),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2177),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2177),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2271),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2400),
.B(n_1953),
.Y(n_2794)
);

INVx2_ASAP7_75t_SL g2795 ( 
.A(n_2475),
.Y(n_2795)
);

BUFx6f_ASAP7_75t_L g2796 ( 
.A(n_2271),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2173),
.B(n_1131),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2180),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2180),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2188),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2188),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2197),
.Y(n_2802)
);

AOI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2124),
.A2(n_1953),
.B1(n_1979),
.B2(n_1976),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2197),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2204),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2204),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2178),
.B(n_1133),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2115),
.B(n_1976),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2124),
.A2(n_1979),
.B1(n_1985),
.B2(n_1983),
.Y(n_2809)
);

AND2x6_ASAP7_75t_L g2810 ( 
.A(n_2359),
.B(n_1983),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2300),
.Y(n_2811)
);

OAI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2181),
.A2(n_946),
.B1(n_948),
.B2(n_930),
.Y(n_2812)
);

INVx4_ASAP7_75t_L g2813 ( 
.A(n_2300),
.Y(n_2813)
);

AND2x6_ASAP7_75t_L g2814 ( 
.A(n_2361),
.B(n_1985),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2205),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2124),
.B(n_1996),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2278),
.B(n_1651),
.Y(n_2817)
);

INVx1_ASAP7_75t_SL g2818 ( 
.A(n_2079),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2249),
.B(n_2108),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2400),
.B(n_1996),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2183),
.B(n_1134),
.Y(n_2821)
);

AND2x6_ASAP7_75t_L g2822 ( 
.A(n_2363),
.B(n_2376),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_2079),
.B(n_1558),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2205),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2300),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2371),
.B(n_1999),
.Y(n_2826)
);

INVx2_ASAP7_75t_SL g2827 ( 
.A(n_2475),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2214),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2235),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2353),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2214),
.Y(n_2831)
);

BUFx2_ASAP7_75t_L g2832 ( 
.A(n_2324),
.Y(n_2832)
);

BUFx4f_ASAP7_75t_L g2833 ( 
.A(n_2229),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2341),
.B(n_1136),
.Y(n_2834)
);

AND2x6_ASAP7_75t_L g2835 ( 
.A(n_2380),
.B(n_2449),
.Y(n_2835)
);

BUFx2_ASAP7_75t_L g2836 ( 
.A(n_2189),
.Y(n_2836)
);

AND2x6_ASAP7_75t_L g2837 ( 
.A(n_2449),
.B(n_1999),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2216),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2081),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2216),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2108),
.B(n_1137),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2221),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2371),
.B(n_2003),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2221),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2447),
.B(n_2003),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2223),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2406),
.B(n_2011),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2406),
.B(n_2011),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2223),
.Y(n_2849)
);

NAND3xp33_ASAP7_75t_L g2850 ( 
.A(n_2476),
.B(n_2018),
.C(n_2017),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2224),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2399),
.B(n_2401),
.Y(n_2852)
);

BUFx3_ASAP7_75t_L g2853 ( 
.A(n_2229),
.Y(n_2853)
);

BUFx6f_ASAP7_75t_L g2854 ( 
.A(n_2300),
.Y(n_2854)
);

AND2x6_ASAP7_75t_L g2855 ( 
.A(n_2456),
.B(n_2017),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2310),
.Y(n_2856)
);

INVx1_ASAP7_75t_SL g2857 ( 
.A(n_2347),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2224),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2319),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2330),
.B(n_1139),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2310),
.Y(n_2861)
);

AND2x4_ASAP7_75t_L g2862 ( 
.A(n_2447),
.B(n_2018),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2353),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2228),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2330),
.B(n_1141),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2228),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2347),
.B(n_1378),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2233),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2233),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2114),
.B(n_2061),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2234),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2448),
.B(n_2455),
.Y(n_2872)
);

INVx4_ASAP7_75t_SL g2873 ( 
.A(n_2461),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2234),
.B(n_2035),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2237),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2479),
.B(n_2035),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2152),
.B(n_1142),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2237),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2239),
.Y(n_2879)
);

AND2x6_ASAP7_75t_L g2880 ( 
.A(n_2456),
.B(n_2048),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2239),
.B(n_2048),
.Y(n_2881)
);

BUFx3_ASAP7_75t_L g2882 ( 
.A(n_2229),
.Y(n_2882)
);

NAND2xp33_ASAP7_75t_L g2883 ( 
.A(n_2381),
.B(n_2052),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2245),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2114),
.B(n_2063),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2245),
.Y(n_2886)
);

AND2x4_ASAP7_75t_L g2887 ( 
.A(n_2321),
.B(n_2052),
.Y(n_2887)
);

NAND2x1p5_ASAP7_75t_L g2888 ( 
.A(n_2117),
.B(n_2055),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2328),
.B(n_2071),
.Y(n_2889)
);

NAND2x1p5_ASAP7_75t_L g2890 ( 
.A(n_2117),
.B(n_2055),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2152),
.B(n_1143),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2085),
.Y(n_2892)
);

BUFx2_ASAP7_75t_L g2893 ( 
.A(n_2248),
.Y(n_2893)
);

NAND2x1p5_ASAP7_75t_L g2894 ( 
.A(n_2117),
.B(n_2058),
.Y(n_2894)
);

INVx4_ASAP7_75t_SL g2895 ( 
.A(n_2461),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2250),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2250),
.B(n_2058),
.Y(n_2897)
);

AND2x4_ASAP7_75t_L g2898 ( 
.A(n_2333),
.B(n_2061),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2350),
.B(n_2063),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_2340),
.B(n_1557),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2251),
.B(n_2050),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2251),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2316),
.B(n_1145),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2252),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2185),
.B(n_594),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2252),
.B(n_2053),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2404),
.Y(n_2907)
);

INVxp67_ASAP7_75t_L g2908 ( 
.A(n_2299),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2258),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2258),
.Y(n_2910)
);

BUFx6f_ASAP7_75t_L g2911 ( 
.A(n_2310),
.Y(n_2911)
);

NOR2x1p5_ASAP7_75t_L g2912 ( 
.A(n_2432),
.B(n_1950),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2492),
.B(n_2089),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2754),
.A2(n_2151),
.B(n_2125),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2547),
.B(n_2320),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2492),
.B(n_2091),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2523),
.B(n_2331),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2509),
.Y(n_2918)
);

O2A1O1Ixp33_ASAP7_75t_L g2919 ( 
.A1(n_2597),
.A2(n_2299),
.B(n_2350),
.C(n_2176),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2547),
.B(n_2185),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2523),
.A2(n_2381),
.B1(n_2176),
.B2(n_2171),
.Y(n_2921)
);

INVx2_ASAP7_75t_SL g2922 ( 
.A(n_2491),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_2780),
.A2(n_2217),
.B1(n_2365),
.B2(n_2349),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2541),
.B(n_2097),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2668),
.B(n_2171),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2503),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2526),
.B(n_2099),
.Y(n_2927)
);

AOI22xp33_ASAP7_75t_L g2928 ( 
.A1(n_2780),
.A2(n_2217),
.B1(n_2349),
.B2(n_2339),
.Y(n_2928)
);

A2O1A1Ixp33_ASAP7_75t_SL g2929 ( 
.A1(n_2526),
.A2(n_2161),
.B(n_2130),
.C(n_2159),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2566),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_SL g2931 ( 
.A(n_2668),
.B(n_2100),
.Y(n_2931)
);

NAND2x1p5_ASAP7_75t_L g2932 ( 
.A(n_2490),
.B(n_2378),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2527),
.B(n_2531),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2527),
.A2(n_2208),
.B1(n_2312),
.B2(n_2298),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_L g2935 ( 
.A(n_2622),
.B(n_2280),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2531),
.B(n_2687),
.Y(n_2936)
);

NOR2xp67_ASAP7_75t_L g2937 ( 
.A(n_2486),
.B(n_2439),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2687),
.B(n_2104),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_2872),
.B(n_2105),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2767),
.B(n_2111),
.Y(n_2940)
);

OR2x2_ASAP7_75t_L g2941 ( 
.A(n_2648),
.B(n_2316),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2501),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2505),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2622),
.B(n_2281),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2767),
.B(n_2112),
.Y(n_2945)
);

BUFx4_ASAP7_75t_L g2946 ( 
.A(n_2685),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2872),
.B(n_2113),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2551),
.B(n_2118),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2508),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2819),
.B(n_2120),
.Y(n_2950)
);

BUFx6f_ASAP7_75t_L g2951 ( 
.A(n_2645),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_SL g2952 ( 
.A(n_2818),
.B(n_2122),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2818),
.B(n_2136),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2500),
.B(n_2137),
.Y(n_2954)
);

NAND3xp33_ASAP7_75t_L g2955 ( 
.A(n_2597),
.B(n_2306),
.C(n_2451),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2513),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2551),
.B(n_2145),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2672),
.B(n_2384),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2517),
.A2(n_2339),
.B1(n_2281),
.B2(n_2161),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2747),
.B(n_2714),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2839),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2714),
.B(n_2386),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2741),
.B(n_2388),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2553),
.B(n_2389),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2537),
.Y(n_2965)
);

O2A1O1Ixp33_ASAP7_75t_L g2966 ( 
.A1(n_2517),
.A2(n_2460),
.B(n_2451),
.C(n_2397),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2750),
.B(n_2402),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2581),
.B(n_2460),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2611),
.A2(n_2381),
.B1(n_2215),
.B2(n_2243),
.Y(n_2969)
);

AOI22xp5_ASAP7_75t_SL g2970 ( 
.A1(n_2584),
.A2(n_2264),
.B1(n_2290),
.B2(n_2109),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2751),
.B(n_2405),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2711),
.B(n_2436),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2839),
.Y(n_2973)
);

AND2x2_ASAP7_75t_SL g2974 ( 
.A(n_2502),
.B(n_2110),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_SL g2975 ( 
.A(n_2623),
.B(n_2332),
.Y(n_2975)
);

INVx3_ASAP7_75t_L g2976 ( 
.A(n_2501),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2592),
.B(n_2443),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2700),
.B(n_2444),
.Y(n_2978)
);

AND2x6_ASAP7_75t_SL g2979 ( 
.A(n_2867),
.B(n_2277),
.Y(n_2979)
);

INVxp67_ASAP7_75t_L g2980 ( 
.A(n_2509),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2700),
.B(n_2445),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2550),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2500),
.B(n_2446),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2740),
.B(n_2450),
.Y(n_2984)
);

HB1xp67_ASAP7_75t_L g2985 ( 
.A(n_2497),
.Y(n_2985)
);

BUFx6f_ASAP7_75t_L g2986 ( 
.A(n_2645),
.Y(n_2986)
);

INVx2_ASAP7_75t_SL g2987 ( 
.A(n_2698),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2619),
.B(n_2452),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2554),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2892),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2770),
.B(n_2841),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2892),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2770),
.B(n_2453),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2852),
.B(n_2381),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2611),
.A2(n_2381),
.B1(n_2215),
.B2(n_2243),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2619),
.B(n_2344),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2852),
.B(n_2191),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2557),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2569),
.Y(n_2999)
);

O2A1O1Ixp33_ASAP7_75t_L g3000 ( 
.A1(n_2733),
.A2(n_2397),
.B(n_2368),
.C(n_2298),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_SL g3001 ( 
.A1(n_2788),
.A2(n_2264),
.B1(n_2290),
.B2(n_2348),
.Y(n_3001)
);

INVx1_ASAP7_75t_SL g3002 ( 
.A(n_2512),
.Y(n_3002)
);

NOR2xp67_ASAP7_75t_L g3003 ( 
.A(n_2643),
.B(n_2442),
.Y(n_3003)
);

AOI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2754),
.A2(n_2304),
.B(n_2151),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2571),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2652),
.A2(n_2368),
.B1(n_2312),
.B2(n_2352),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2535),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2484),
.Y(n_3008)
);

AND2x6_ASAP7_75t_SL g3009 ( 
.A(n_2771),
.B(n_2277),
.Y(n_3009)
);

AND2x6_ASAP7_75t_SL g3010 ( 
.A(n_2616),
.B(n_2277),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2593),
.B(n_2194),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2530),
.B(n_2462),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2487),
.Y(n_3013)
);

NAND2xp33_ASAP7_75t_L g3014 ( 
.A(n_2501),
.B(n_2480),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2577),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2593),
.B(n_2198),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2502),
.A2(n_2257),
.B1(n_2190),
.B2(n_2130),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2488),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2489),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2516),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2621),
.B(n_2618),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2834),
.B(n_2203),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2578),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2493),
.A2(n_2908),
.B1(n_2766),
.B2(n_2556),
.Y(n_3024)
);

AND2x4_ASAP7_75t_L g3025 ( 
.A(n_2514),
.B(n_2472),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2756),
.B(n_2206),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2877),
.B(n_2207),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2754),
.A2(n_2431),
.B(n_2151),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2702),
.A2(n_2477),
.B1(n_2463),
.B2(n_2465),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_SL g3030 ( 
.A(n_2713),
.B(n_2409),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2495),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2530),
.B(n_2543),
.Y(n_3032)
);

BUFx3_ASAP7_75t_L g3033 ( 
.A(n_2664),
.Y(n_3033)
);

NAND3xp33_ASAP7_75t_SL g3034 ( 
.A(n_2702),
.B(n_2442),
.C(n_2464),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2891),
.B(n_2213),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2860),
.B(n_2219),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2506),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2737),
.B(n_2639),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2865),
.B(n_2222),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2582),
.Y(n_3040)
);

OAI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2857),
.A2(n_2473),
.B1(n_2230),
.B2(n_2242),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2543),
.B(n_2544),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_L g3043 ( 
.A1(n_2518),
.A2(n_2257),
.B1(n_2190),
.B2(n_2159),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2908),
.B(n_2226),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2518),
.A2(n_2110),
.B1(n_2167),
.B2(n_2295),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_SL g3046 ( 
.A(n_2544),
.B(n_2418),
.Y(n_3046)
);

NOR3x1_ASAP7_75t_L g3047 ( 
.A(n_2485),
.B(n_1149),
.C(n_1148),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2621),
.B(n_2284),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2563),
.B(n_2418),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2899),
.B(n_2254),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2511),
.Y(n_3051)
);

NOR2xp67_ASAP7_75t_L g3052 ( 
.A(n_2903),
.B(n_2255),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2606),
.Y(n_3053)
);

A2O1A1Ixp33_ASAP7_75t_L g3054 ( 
.A1(n_2493),
.A2(n_2149),
.B(n_2295),
.C(n_2263),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2899),
.B(n_2708),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2585),
.Y(n_3056)
);

CKINVDCx8_ASAP7_75t_R g3057 ( 
.A(n_2893),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2708),
.B(n_2259),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2754),
.A2(n_2304),
.B(n_2125),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2614),
.B(n_2266),
.Y(n_3060)
);

INVx4_ASAP7_75t_L g3061 ( 
.A(n_2504),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2615),
.B(n_2286),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2515),
.B(n_2125),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2529),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2604),
.Y(n_3065)
);

NOR3xp33_ASAP7_75t_L g3066 ( 
.A(n_2485),
.B(n_2416),
.C(n_2392),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2757),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2532),
.Y(n_3068)
);

AO22x1_ASAP7_75t_L g3069 ( 
.A1(n_2647),
.A2(n_2000),
.B1(n_954),
.B2(n_957),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_2655),
.B(n_2294),
.Y(n_3070)
);

NAND2xp33_ASAP7_75t_L g3071 ( 
.A(n_2504),
.B(n_2480),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2710),
.B(n_2294),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2556),
.B(n_2304),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2761),
.B(n_2378),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2795),
.B(n_2827),
.Y(n_3075)
);

AOI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2817),
.A2(n_2165),
.B1(n_2167),
.B2(n_2461),
.Y(n_3076)
);

A2O1A1Ixp33_ASAP7_75t_L g3077 ( 
.A1(n_2519),
.A2(n_2889),
.B(n_2561),
.C(n_2766),
.Y(n_3077)
);

NAND3xp33_ASAP7_75t_L g3078 ( 
.A(n_2640),
.B(n_2424),
.C(n_2414),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2504),
.Y(n_3079)
);

OAI22xp5_ASAP7_75t_SL g3080 ( 
.A1(n_2788),
.A2(n_2329),
.B1(n_2419),
.B2(n_962),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2889),
.B(n_2378),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2733),
.A2(n_2480),
.B1(n_2461),
.B2(n_2471),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2533),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2876),
.B(n_2563),
.Y(n_3084)
);

INVxp67_ASAP7_75t_SL g3085 ( 
.A(n_2723),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_2519),
.A2(n_2431),
.B1(n_2438),
.B2(n_2404),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2876),
.B(n_2431),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2567),
.B(n_2438),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2857),
.B(n_2356),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2538),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_2730),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2567),
.B(n_2438),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2620),
.B(n_2418),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2514),
.B(n_2131),
.Y(n_3094)
);

INVx2_ASAP7_75t_SL g3095 ( 
.A(n_2576),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2539),
.Y(n_3096)
);

A2O1A1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2561),
.A2(n_1788),
.B(n_2356),
.C(n_2429),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2620),
.B(n_2693),
.Y(n_3098)
);

AND2x6_ASAP7_75t_L g3099 ( 
.A(n_2784),
.B(n_2131),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2629),
.B(n_2294),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2629),
.B(n_2272),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2542),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2609),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2617),
.A2(n_2461),
.B1(n_2480),
.B2(n_2471),
.Y(n_3104)
);

AOI22xp33_ASAP7_75t_L g3105 ( 
.A1(n_2627),
.A2(n_2480),
.B1(n_2471),
.B2(n_2123),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2832),
.B(n_2165),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_2772),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_2516),
.B(n_2435),
.Y(n_3108)
);

INVx2_ASAP7_75t_SL g3109 ( 
.A(n_2676),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2510),
.Y(n_3110)
);

INVxp67_ASAP7_75t_L g3111 ( 
.A(n_2528),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2667),
.A2(n_2474),
.B1(n_2323),
.B2(n_2468),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2613),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2797),
.B(n_2457),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2807),
.B(n_2457),
.Y(n_3115)
);

AOI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2579),
.A2(n_2123),
.B1(n_2459),
.B2(n_2323),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2626),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2821),
.B(n_2466),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2726),
.B(n_2466),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_SL g3120 ( 
.A(n_2693),
.B(n_2131),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2719),
.B(n_2379),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2545),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2632),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2608),
.B(n_2470),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2549),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2659),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2726),
.B(n_2467),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2630),
.A2(n_2470),
.B1(n_2482),
.B2(n_2467),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2579),
.A2(n_2474),
.B1(n_2060),
.B2(n_2062),
.Y(n_3129)
);

O2A1O1Ixp5_ASAP7_75t_L g3130 ( 
.A1(n_2534),
.A2(n_2301),
.B(n_2483),
.C(n_2482),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2719),
.B(n_2411),
.Y(n_3131)
);

INVx3_ASAP7_75t_L g3132 ( 
.A(n_2490),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2612),
.B(n_2483),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2633),
.B(n_2310),
.Y(n_3134)
);

NOR3xp33_ASAP7_75t_L g3135 ( 
.A(n_2586),
.B(n_1155),
.C(n_1154),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_2859),
.B(n_2329),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2665),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2635),
.B(n_2342),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2637),
.A2(n_2650),
.B1(n_2653),
.B2(n_2649),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2682),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2552),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_2764),
.A2(n_2072),
.B1(n_2073),
.B2(n_2057),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2654),
.B(n_2342),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2657),
.B(n_2342),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2555),
.Y(n_3145)
);

OAI221xp5_ASAP7_75t_L g3146 ( 
.A1(n_2575),
.A2(n_2720),
.B1(n_2823),
.B2(n_2749),
.C(n_2836),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2498),
.Y(n_3147)
);

AND2x6_ASAP7_75t_L g3148 ( 
.A(n_2784),
.B(n_2433),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2704),
.Y(n_3149)
);

AND2x4_ASAP7_75t_SL g3150 ( 
.A(n_2524),
.B(n_2342),
.Y(n_3150)
);

CKINVDCx5p33_ASAP7_75t_R g3151 ( 
.A(n_2525),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2721),
.Y(n_3152)
);

INVx2_ASAP7_75t_SL g3153 ( 
.A(n_2684),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2764),
.B(n_2345),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2658),
.B(n_2345),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2645),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2782),
.B(n_2345),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2558),
.Y(n_3158)
);

NOR3xp33_ASAP7_75t_L g3159 ( 
.A(n_2823),
.B(n_2662),
.C(n_2651),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_2663),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2598),
.B(n_2272),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2660),
.B(n_2345),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2575),
.B(n_2244),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2670),
.B(n_2673),
.Y(n_3164)
);

A2O1A1Ixp33_ASAP7_75t_L g3165 ( 
.A1(n_2870),
.A2(n_1635),
.B(n_1578),
.C(n_1579),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_2664),
.Y(n_3166)
);

INVx4_ASAP7_75t_L g3167 ( 
.A(n_2522),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_2782),
.B(n_2379),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_2524),
.B(n_2379),
.Y(n_3169)
);

BUFx3_ASAP7_75t_L g3170 ( 
.A(n_2853),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2540),
.B(n_2379),
.Y(n_3171)
);

INVxp33_ASAP7_75t_L g3172 ( 
.A(n_2680),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2727),
.Y(n_3173)
);

INVx2_ASAP7_75t_SL g3174 ( 
.A(n_2695),
.Y(n_3174)
);

NAND2x1_ASAP7_75t_L g3175 ( 
.A(n_2507),
.B(n_2498),
.Y(n_3175)
);

O2A1O1Ixp5_ASAP7_75t_L g3176 ( 
.A1(n_2534),
.A2(n_2396),
.B(n_1691),
.C(n_1694),
.Y(n_3176)
);

NOR2xp33_ASAP7_75t_L g3177 ( 
.A(n_2847),
.B(n_2329),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2675),
.B(n_2411),
.Y(n_3178)
);

BUFx3_ASAP7_75t_L g3179 ( 
.A(n_2882),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2625),
.B(n_2419),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2731),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2559),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2847),
.B(n_2419),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_2540),
.B(n_2411),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2678),
.B(n_2411),
.Y(n_3185)
);

NOR3xp33_ASAP7_75t_L g3186 ( 
.A(n_2720),
.B(n_1160),
.C(n_1158),
.Y(n_3186)
);

NAND3xp33_ASAP7_75t_L g3187 ( 
.A(n_2749),
.B(n_2000),
.C(n_773),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2683),
.B(n_2415),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2735),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2546),
.B(n_2415),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_2689),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2744),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2779),
.B(n_1378),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2661),
.B(n_1161),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2848),
.B(n_2415),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2848),
.B(n_2415),
.Y(n_3196)
);

AOI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_2589),
.A2(n_2600),
.B1(n_2601),
.B2(n_2588),
.Y(n_3197)
);

AOI21x1_ASAP7_75t_L g3198 ( 
.A1(n_2697),
.A2(n_1578),
.B(n_1560),
.Y(n_3198)
);

AOI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_2677),
.A2(n_2351),
.B(n_2309),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2560),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_2686),
.A2(n_954),
.B1(n_957),
.B2(n_948),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2564),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2688),
.B(n_2433),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_SL g3204 ( 
.A(n_2546),
.B(n_2433),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2565),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_2691),
.A2(n_961),
.B1(n_965),
.B2(n_959),
.Y(n_3206)
);

AO22x1_ASAP7_75t_L g3207 ( 
.A1(n_2752),
.A2(n_2000),
.B1(n_966),
.B2(n_775),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2580),
.B(n_2433),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2692),
.A2(n_966),
.B1(n_776),
.B2(n_779),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2699),
.B(n_1635),
.Y(n_3210)
);

INVx2_ASAP7_75t_SL g3211 ( 
.A(n_2713),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2705),
.B(n_2706),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_2580),
.B(n_2309),
.Y(n_3213)
);

NAND2xp33_ASAP7_75t_L g3214 ( 
.A(n_2574),
.B(n_2247),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_2709),
.B(n_1635),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2722),
.B(n_1560),
.Y(n_3216)
);

AND2x4_ASAP7_75t_SL g3217 ( 
.A(n_2525),
.B(n_1727),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2725),
.B(n_1579),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_SL g3219 ( 
.A(n_2667),
.B(n_2681),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2729),
.B(n_1971),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_SL g3221 ( 
.A(n_2681),
.B(n_2661),
.Y(n_3221)
);

INVxp67_ASAP7_75t_L g3222 ( 
.A(n_2690),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2734),
.B(n_1971),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2568),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2739),
.B(n_1971),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2690),
.B(n_2309),
.Y(n_3226)
);

OAI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_2610),
.A2(n_2351),
.B1(n_2309),
.B2(n_604),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_2755),
.A2(n_780),
.B1(n_783),
.B2(n_768),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_2758),
.B(n_1974),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2760),
.B(n_1974),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2583),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_2610),
.B(n_2351),
.Y(n_3232)
);

INVx2_ASAP7_75t_SL g3233 ( 
.A(n_2833),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2715),
.B(n_2027),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2646),
.A2(n_2351),
.B1(n_604),
.B2(n_609),
.Y(n_3235)
);

AO22x1_ASAP7_75t_L g3236 ( 
.A1(n_2933),
.A2(n_2752),
.B1(n_2787),
.B2(n_2768),
.Y(n_3236)
);

BUFx12f_ASAP7_75t_L g3237 ( 
.A(n_3053),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_2930),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_3094),
.B(n_3025),
.Y(n_3239)
);

BUFx12f_ASAP7_75t_SL g3240 ( 
.A(n_3180),
.Y(n_3240)
);

NAND3xp33_ASAP7_75t_SL g3241 ( 
.A(n_3066),
.B(n_2787),
.C(n_2768),
.Y(n_3241)
);

BUFx2_ASAP7_75t_L g3242 ( 
.A(n_3007),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_2935),
.A2(n_2548),
.B1(n_2590),
.B2(n_2656),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2936),
.B(n_2900),
.Y(n_3244)
);

AND2x6_ASAP7_75t_SL g3245 ( 
.A(n_3193),
.B(n_2525),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_3033),
.Y(n_3246)
);

BUFx6f_ASAP7_75t_L g3247 ( 
.A(n_2951),
.Y(n_3247)
);

NOR3xp33_ASAP7_75t_L g3248 ( 
.A(n_2917),
.B(n_2724),
.C(n_2812),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2926),
.Y(n_3249)
);

A2O1A1Ixp33_ASAP7_75t_L g3250 ( 
.A1(n_2968),
.A2(n_2885),
.B(n_2883),
.C(n_2850),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2935),
.A2(n_2548),
.B1(n_2590),
.B2(n_2656),
.Y(n_3251)
);

OR2x2_ASAP7_75t_L g3252 ( 
.A(n_2941),
.B(n_2887),
.Y(n_3252)
);

INVx3_ASAP7_75t_L g3253 ( 
.A(n_3094),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3008),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3013),
.Y(n_3255)
);

BUFx6f_ASAP7_75t_L g3256 ( 
.A(n_2951),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_2958),
.B(n_2521),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_2943),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2913),
.B(n_2794),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3018),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3019),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3031),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3037),
.Y(n_3263)
);

BUFx3_ASAP7_75t_L g3264 ( 
.A(n_3166),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3051),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2951),
.Y(n_3266)
);

INVx4_ASAP7_75t_L g3267 ( 
.A(n_2951),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3066),
.A2(n_2600),
.B1(n_2601),
.B2(n_2589),
.Y(n_3268)
);

INVx5_ASAP7_75t_L g3269 ( 
.A(n_2986),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2916),
.B(n_2794),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_2977),
.B(n_2572),
.Y(n_3271)
);

HB1xp67_ASAP7_75t_L g3272 ( 
.A(n_2918),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2949),
.Y(n_3273)
);

NAND2x1p5_ASAP7_75t_L g3274 ( 
.A(n_2922),
.B(n_2833),
.Y(n_3274)
);

AND2x4_ASAP7_75t_SL g3275 ( 
.A(n_2985),
.B(n_2522),
.Y(n_3275)
);

INVx4_ASAP7_75t_L g3276 ( 
.A(n_2986),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3175),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2960),
.B(n_2820),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_3146),
.A2(n_2845),
.B1(n_2862),
.B2(n_2820),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_L g3280 ( 
.A(n_2977),
.B(n_2790),
.Y(n_3280)
);

OAI22xp5_ASAP7_75t_SL g3281 ( 
.A1(n_3001),
.A2(n_2572),
.B1(n_2573),
.B2(n_787),
.Y(n_3281)
);

CKINVDCx8_ASAP7_75t_R g3282 ( 
.A(n_3009),
.Y(n_3282)
);

BUFx3_ASAP7_75t_L g3283 ( 
.A(n_3170),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2956),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_3179),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3164),
.Y(n_3286)
);

INVx3_ASAP7_75t_L g3287 ( 
.A(n_3132),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2965),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2988),
.B(n_2845),
.Y(n_3289)
);

CKINVDCx20_ASAP7_75t_R g3290 ( 
.A(n_3067),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_3025),
.B(n_2786),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2927),
.B(n_2862),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_2985),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3212),
.Y(n_3294)
);

OR2x2_ASAP7_75t_SL g3295 ( 
.A(n_2955),
.B(n_2707),
.Y(n_3295)
);

BUFx12f_ASAP7_75t_SL g3296 ( 
.A(n_3070),
.Y(n_3296)
);

BUFx3_ASAP7_75t_L g3297 ( 
.A(n_3095),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3064),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3068),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_2988),
.B(n_2646),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2948),
.B(n_2718),
.Y(n_3301)
);

OR2x2_ASAP7_75t_SL g3302 ( 
.A(n_3187),
.B(n_2912),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2957),
.B(n_2963),
.Y(n_3303)
);

AND2x4_ASAP7_75t_SL g3304 ( 
.A(n_3061),
.B(n_2522),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3083),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_SL g3306 ( 
.A(n_3021),
.B(n_2666),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_L g3307 ( 
.A(n_2996),
.B(n_2753),
.Y(n_3307)
);

BUFx4f_ASAP7_75t_L g3308 ( 
.A(n_3211),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_2980),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_SL g3310 ( 
.A(n_2996),
.B(n_2666),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3090),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2972),
.B(n_2718),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3096),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2967),
.B(n_2728),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_2944),
.A2(n_2915),
.B1(n_3159),
.B2(n_3042),
.Y(n_3315)
);

OR2x6_ASAP7_75t_L g3316 ( 
.A(n_3233),
.B(n_2574),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2982),
.Y(n_3317)
);

NOR2x1_ASAP7_75t_R g3318 ( 
.A(n_3151),
.B(n_2499),
.Y(n_3318)
);

BUFx12f_ASAP7_75t_L g3319 ( 
.A(n_3107),
.Y(n_3319)
);

A2O1A1Ixp33_ASAP7_75t_L g3320 ( 
.A1(n_2919),
.A2(n_2885),
.B(n_2850),
.C(n_2694),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3102),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_SL g3322 ( 
.A1(n_2970),
.A2(n_2644),
.B1(n_2671),
.B2(n_2574),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3122),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3125),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_2986),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_2989),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2980),
.B(n_2753),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2971),
.B(n_2728),
.Y(n_3328)
);

INVx2_ASAP7_75t_SL g3329 ( 
.A(n_3091),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2998),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3141),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3038),
.B(n_3194),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_2986),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_2999),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2984),
.B(n_2763),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3005),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_2964),
.B(n_2887),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3145),
.Y(n_3338)
);

INVxp67_ASAP7_75t_L g3339 ( 
.A(n_3110),
.Y(n_3339)
);

NAND3xp33_ASAP7_75t_L g3340 ( 
.A(n_3159),
.B(n_1163),
.C(n_1162),
.Y(n_3340)
);

BUFx6f_ASAP7_75t_L g3341 ( 
.A(n_3156),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_3156),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3158),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_2987),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3182),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3200),
.Y(n_3346)
);

INVx2_ASAP7_75t_SL g3347 ( 
.A(n_3002),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3202),
.Y(n_3348)
);

HB1xp67_ASAP7_75t_L g3349 ( 
.A(n_3020),
.Y(n_3349)
);

CKINVDCx5p33_ASAP7_75t_R g3350 ( 
.A(n_3057),
.Y(n_3350)
);

BUFx3_ASAP7_75t_L g3351 ( 
.A(n_3153),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2997),
.B(n_2763),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3015),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_3052),
.B(n_2694),
.Y(n_3354)
);

INVx4_ASAP7_75t_L g3355 ( 
.A(n_3156),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3023),
.Y(n_3356)
);

OR2x6_ASAP7_75t_L g3357 ( 
.A(n_2937),
.B(n_2644),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3205),
.Y(n_3358)
);

INVx3_ASAP7_75t_L g3359 ( 
.A(n_3132),
.Y(n_3359)
);

HB1xp67_ASAP7_75t_L g3360 ( 
.A(n_3020),
.Y(n_3360)
);

BUFx2_ASAP7_75t_L g3361 ( 
.A(n_3191),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3224),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_2991),
.B(n_2712),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3231),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_2938),
.B(n_2940),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3040),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3056),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_3197),
.B(n_2786),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2945),
.B(n_2712),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3060),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3062),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3108),
.B(n_2588),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3065),
.Y(n_3373)
);

INVxp67_ASAP7_75t_L g3374 ( 
.A(n_3111),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3103),
.Y(n_3375)
);

AND2x4_ASAP7_75t_L g3376 ( 
.A(n_3098),
.B(n_2786),
.Y(n_3376)
);

INVx4_ASAP7_75t_L g3377 ( 
.A(n_3156),
.Y(n_3377)
);

AOI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3101),
.A2(n_2822),
.B1(n_2898),
.B2(n_2808),
.Y(n_3378)
);

AND2x4_ASAP7_75t_L g3379 ( 
.A(n_3222),
.B(n_2499),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3111),
.B(n_2785),
.Y(n_3380)
);

CKINVDCx20_ASAP7_75t_R g3381 ( 
.A(n_3174),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3113),
.Y(n_3382)
);

BUFx12f_ASAP7_75t_L g3383 ( 
.A(n_3010),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3100),
.A2(n_2822),
.B1(n_2898),
.B2(n_2808),
.Y(n_3384)
);

INVx5_ASAP7_75t_L g3385 ( 
.A(n_3061),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3108),
.B(n_2536),
.Y(n_3386)
);

AOI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3072),
.A2(n_2822),
.B1(n_2769),
.B2(n_2745),
.Y(n_3387)
);

INVx1_ASAP7_75t_SL g3388 ( 
.A(n_3109),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3117),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_3147),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3123),
.Y(n_3391)
);

INVx3_ASAP7_75t_L g3392 ( 
.A(n_3147),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3022),
.B(n_2536),
.Y(n_3393)
);

INVx5_ASAP7_75t_L g3394 ( 
.A(n_3148),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2962),
.B(n_2924),
.Y(n_3395)
);

NAND3xp33_ASAP7_75t_SL g3396 ( 
.A(n_2966),
.B(n_792),
.C(n_786),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3126),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3036),
.B(n_2697),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3032),
.A2(n_2822),
.B1(n_2905),
.B2(n_2596),
.Y(n_3399)
);

BUFx4f_ASAP7_75t_L g3400 ( 
.A(n_3161),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_2961),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3222),
.B(n_2746),
.Y(n_3402)
);

AND2x6_ASAP7_75t_SL g3403 ( 
.A(n_3048),
.B(n_1168),
.Y(n_3403)
);

CKINVDCx5p33_ASAP7_75t_R g3404 ( 
.A(n_2979),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_3167),
.Y(n_3405)
);

INVx3_ASAP7_75t_L g3406 ( 
.A(n_2932),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3137),
.Y(n_3407)
);

AOI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_3177),
.A2(n_2769),
.B1(n_2745),
.B2(n_2835),
.Y(n_3408)
);

BUFx6f_ASAP7_75t_L g3409 ( 
.A(n_3167),
.Y(n_3409)
);

BUFx3_ASAP7_75t_L g3410 ( 
.A(n_2973),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3140),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3084),
.B(n_2496),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_3172),
.B(n_2785),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_2932),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3039),
.B(n_2677),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_2939),
.B(n_2496),
.Y(n_3416)
);

INVx2_ASAP7_75t_SL g3417 ( 
.A(n_3217),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3149),
.Y(n_3418)
);

CKINVDCx5p33_ASAP7_75t_R g3419 ( 
.A(n_3191),
.Y(n_3419)
);

INVx2_ASAP7_75t_SL g3420 ( 
.A(n_2990),
.Y(n_3420)
);

AND2x6_ASAP7_75t_L g3421 ( 
.A(n_3047),
.B(n_2494),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3152),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3089),
.B(n_2829),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_2947),
.B(n_2494),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3173),
.Y(n_3425)
);

INVx2_ASAP7_75t_SL g3426 ( 
.A(n_2992),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3012),
.B(n_2624),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_3030),
.B(n_2562),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3089),
.B(n_2978),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3181),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3189),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3192),
.Y(n_3432)
);

INVx4_ASAP7_75t_L g3433 ( 
.A(n_3150),
.Y(n_3433)
);

INVx4_ASAP7_75t_L g3434 ( 
.A(n_2942),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2993),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3114),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3029),
.B(n_2562),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3115),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3119),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3118),
.Y(n_3440)
);

OR2x6_ASAP7_75t_L g3441 ( 
.A(n_3003),
.B(n_2644),
.Y(n_3441)
);

CKINVDCx5p33_ASAP7_75t_R g3442 ( 
.A(n_3106),
.Y(n_3442)
);

BUFx3_ASAP7_75t_L g3443 ( 
.A(n_3106),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_SL g3444 ( 
.A1(n_3300),
.A2(n_3077),
.B(n_2929),
.C(n_2983),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_3301),
.A2(n_3214),
.B(n_3081),
.Y(n_3445)
);

O2A1O1Ixp33_ASAP7_75t_L g3446 ( 
.A1(n_3248),
.A2(n_3034),
.B(n_2954),
.C(n_2950),
.Y(n_3446)
);

OAI22x1_ASAP7_75t_L g3447 ( 
.A1(n_3280),
.A2(n_3006),
.B1(n_3257),
.B2(n_3271),
.Y(n_3447)
);

BUFx3_ASAP7_75t_L g3448 ( 
.A(n_3264),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3249),
.Y(n_3449)
);

BUFx6f_ASAP7_75t_L g3450 ( 
.A(n_3269),
.Y(n_3450)
);

INVx3_ASAP7_75t_L g3451 ( 
.A(n_3291),
.Y(n_3451)
);

BUFx2_ASAP7_75t_L g3452 ( 
.A(n_3419),
.Y(n_3452)
);

OAI22xp5_ASAP7_75t_L g3453 ( 
.A1(n_3289),
.A2(n_2959),
.B1(n_3085),
.B2(n_2995),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_3290),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3250),
.A2(n_3055),
.B(n_2925),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3303),
.B(n_3027),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3332),
.B(n_3034),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3338),
.Y(n_3458)
);

BUFx3_ASAP7_75t_L g3459 ( 
.A(n_3283),
.Y(n_3459)
);

AND2x4_ASAP7_75t_L g3460 ( 
.A(n_3291),
.B(n_3120),
.Y(n_3460)
);

O2A1O1Ixp33_ASAP7_75t_L g3461 ( 
.A1(n_3241),
.A2(n_3186),
.B(n_2931),
.C(n_3000),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3338),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3429),
.B(n_2975),
.Y(n_3463)
);

O2A1O1Ixp33_ASAP7_75t_SL g3464 ( 
.A1(n_3310),
.A2(n_3437),
.B(n_3386),
.C(n_3393),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3307),
.B(n_3177),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3343),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3398),
.A2(n_3085),
.B(n_2934),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3396),
.A2(n_2921),
.B(n_2994),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3343),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3415),
.A2(n_3043),
.B(n_3017),
.Y(n_3470)
);

AO22x1_ASAP7_75t_L g3471 ( 
.A1(n_3404),
.A2(n_3136),
.B1(n_3186),
.B2(n_3163),
.Y(n_3471)
);

BUFx4f_ASAP7_75t_SL g3472 ( 
.A(n_3237),
.Y(n_3472)
);

O2A1O1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_3365),
.A2(n_3135),
.B(n_2952),
.C(n_2953),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3395),
.B(n_3035),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3435),
.B(n_2981),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3258),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3273),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3370),
.B(n_3026),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3371),
.B(n_3244),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_3400),
.B(n_3183),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3284),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3243),
.A2(n_3078),
.B1(n_3135),
.B2(n_2974),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3436),
.B(n_3183),
.Y(n_3483)
);

HB1xp67_ASAP7_75t_L g3484 ( 
.A(n_3309),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3436),
.B(n_3201),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3288),
.Y(n_3486)
);

INVx3_ASAP7_75t_L g3487 ( 
.A(n_3253),
.Y(n_3487)
);

OAI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_3315),
.A2(n_2959),
.B1(n_2995),
.B2(n_2969),
.Y(n_3488)
);

AOI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_3312),
.A2(n_3043),
.B(n_3017),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3314),
.A2(n_3071),
.B(n_3014),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3384),
.A2(n_3133),
.B(n_3124),
.C(n_2969),
.Y(n_3491)
);

OAI21xp33_ASAP7_75t_SL g3492 ( 
.A1(n_3328),
.A2(n_2923),
.B(n_2928),
.Y(n_3492)
);

A2O1A1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3378),
.A2(n_3124),
.B(n_3133),
.C(n_2923),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3345),
.Y(n_3494)
);

HB1xp67_ASAP7_75t_L g3495 ( 
.A(n_3293),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_R g3496 ( 
.A(n_3350),
.B(n_2942),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3345),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3346),
.Y(n_3498)
);

HB1xp67_ASAP7_75t_L g3499 ( 
.A(n_3272),
.Y(n_3499)
);

NAND2x1_ASAP7_75t_L g3500 ( 
.A(n_3277),
.B(n_2624),
.Y(n_3500)
);

OR2x6_ASAP7_75t_L g3501 ( 
.A(n_3357),
.B(n_2671),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3320),
.A2(n_3073),
.B(n_3054),
.Y(n_3502)
);

NAND2x1p5_ASAP7_75t_L g3503 ( 
.A(n_3385),
.B(n_2562),
.Y(n_3503)
);

OAI22xp5_ASAP7_75t_L g3504 ( 
.A1(n_3400),
.A2(n_3251),
.B1(n_3442),
.B2(n_3279),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3438),
.B(n_3201),
.Y(n_3505)
);

NOR3xp33_ASAP7_75t_SL g3506 ( 
.A(n_3281),
.B(n_3080),
.C(n_3238),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3438),
.B(n_3206),
.Y(n_3507)
);

INVx3_ASAP7_75t_L g3508 ( 
.A(n_3253),
.Y(n_3508)
);

OR2x6_ASAP7_75t_L g3509 ( 
.A(n_3357),
.B(n_2671),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3240),
.B(n_3069),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_3394),
.A2(n_3045),
.B(n_3105),
.Y(n_3511)
);

AND2x4_ASAP7_75t_L g3512 ( 
.A(n_3239),
.B(n_3376),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3337),
.B(n_3228),
.Y(n_3513)
);

INVx3_ASAP7_75t_L g3514 ( 
.A(n_3405),
.Y(n_3514)
);

INVx2_ASAP7_75t_SL g3515 ( 
.A(n_3308),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3339),
.B(n_3136),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3268),
.A2(n_2928),
.B1(n_3105),
.B2(n_3209),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3292),
.B(n_3041),
.Y(n_3518)
);

INVx4_ASAP7_75t_L g3519 ( 
.A(n_3385),
.Y(n_3519)
);

AND2x4_ASAP7_75t_L g3520 ( 
.A(n_3239),
.B(n_2976),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3421),
.A2(n_3046),
.B1(n_3049),
.B2(n_3041),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3317),
.Y(n_3522)
);

NOR2x1_ASAP7_75t_L g3523 ( 
.A(n_3443),
.B(n_2976),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_R g3524 ( 
.A(n_3381),
.B(n_3079),
.Y(n_3524)
);

AND2x4_ASAP7_75t_L g3525 ( 
.A(n_3376),
.B(n_3079),
.Y(n_3525)
);

A2O1A1Ixp33_ASAP7_75t_L g3526 ( 
.A1(n_3387),
.A2(n_3076),
.B(n_3044),
.C(n_3050),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3440),
.B(n_3058),
.Y(n_3527)
);

BUFx2_ASAP7_75t_L g3528 ( 
.A(n_3242),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3440),
.B(n_3011),
.Y(n_3529)
);

INVxp67_ASAP7_75t_SL g3530 ( 
.A(n_3349),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3335),
.B(n_3016),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3297),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3394),
.A2(n_3045),
.B(n_3004),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3351),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3308),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3326),
.Y(n_3536)
);

AOI21xp5_ASAP7_75t_L g3537 ( 
.A1(n_3394),
.A2(n_3028),
.B(n_2914),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_3368),
.B(n_3160),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3259),
.A2(n_3059),
.B(n_3086),
.Y(n_3539)
);

O2A1O1Ixp33_ASAP7_75t_L g3540 ( 
.A1(n_3374),
.A2(n_2920),
.B(n_3024),
.C(n_3221),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3352),
.B(n_3075),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3330),
.Y(n_3542)
);

O2A1O1Ixp33_ASAP7_75t_L g3543 ( 
.A1(n_3306),
.A2(n_3093),
.B(n_3131),
.C(n_3121),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3278),
.B(n_3207),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3270),
.A2(n_3097),
.B(n_2701),
.Y(n_3545)
);

NOR2xp33_ASAP7_75t_L g3546 ( 
.A(n_3347),
.B(n_3160),
.Y(n_3546)
);

BUFx2_ASAP7_75t_L g3547 ( 
.A(n_3296),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_R g3548 ( 
.A(n_3319),
.B(n_2599),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3286),
.B(n_3127),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_R g3550 ( 
.A(n_3285),
.B(n_2599),
.Y(n_3550)
);

A2O1A1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_3286),
.A2(n_3082),
.B(n_3063),
.C(n_3129),
.Y(n_3551)
);

OAI22x1_ASAP7_75t_L g3552 ( 
.A1(n_3428),
.A2(n_3116),
.B1(n_3142),
.B2(n_3195),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3421),
.A2(n_3383),
.B1(n_3252),
.B2(n_3368),
.Y(n_3553)
);

HB1xp67_ASAP7_75t_L g3554 ( 
.A(n_3360),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_3294),
.A2(n_3082),
.B(n_3092),
.C(n_3088),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3294),
.A2(n_2701),
.B(n_3104),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3346),
.Y(n_3557)
);

OAI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3372),
.A2(n_3139),
.B1(n_3104),
.B2(n_3087),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3439),
.B(n_3195),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3369),
.B(n_3402),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3334),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3348),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_3413),
.B(n_3169),
.Y(n_3563)
);

INVx3_ASAP7_75t_L g3564 ( 
.A(n_3405),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3340),
.A2(n_3196),
.B(n_3157),
.C(n_3168),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3363),
.B(n_3196),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3336),
.Y(n_3567)
);

INVx1_ASAP7_75t_SL g3568 ( 
.A(n_3361),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3348),
.Y(n_3569)
);

BUFx6f_ASAP7_75t_L g3570 ( 
.A(n_3269),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3358),
.Y(n_3571)
);

AOI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_3423),
.A2(n_3219),
.B(n_3199),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3236),
.A2(n_2723),
.B(n_2716),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3421),
.A2(n_3154),
.B1(n_2835),
.B2(n_2717),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3358),
.Y(n_3575)
);

NAND2xp33_ASAP7_75t_L g3576 ( 
.A(n_3421),
.B(n_3099),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3362),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3362),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3327),
.B(n_1170),
.Y(n_3579)
);

CKINVDCx20_ASAP7_75t_R g3580 ( 
.A(n_3282),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_3416),
.B(n_3074),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_SL g3582 ( 
.A1(n_3401),
.A2(n_3410),
.B1(n_3403),
.B2(n_3380),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3353),
.Y(n_3583)
);

O2A1O1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_3354),
.A2(n_3235),
.B(n_3226),
.C(n_3165),
.Y(n_3584)
);

OR2x6_ASAP7_75t_L g3585 ( 
.A(n_3441),
.B(n_3171),
.Y(n_3585)
);

NOR2xp33_ASAP7_75t_L g3586 ( 
.A(n_3388),
.B(n_3216),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3344),
.B(n_3218),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3412),
.B(n_2762),
.Y(n_3588)
);

INVx4_ASAP7_75t_L g3589 ( 
.A(n_3385),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3399),
.A2(n_3234),
.B(n_2843),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3408),
.A2(n_2843),
.B(n_2826),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3277),
.A2(n_2826),
.B(n_3112),
.Y(n_3592)
);

O2A1O1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3420),
.A2(n_1173),
.B(n_1177),
.C(n_1171),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_3245),
.Y(n_3594)
);

BUFx12f_ASAP7_75t_L g3595 ( 
.A(n_3246),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3426),
.A2(n_2829),
.B1(n_3138),
.B2(n_3134),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3364),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3412),
.B(n_2776),
.Y(n_3598)
);

AOI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3416),
.A2(n_798),
.B1(n_802),
.B2(n_797),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_3322),
.A2(n_3144),
.B1(n_3155),
.B2(n_3143),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3356),
.Y(n_3601)
);

NOR3xp33_ASAP7_75t_SL g3602 ( 
.A(n_3364),
.B(n_808),
.C(n_805),
.Y(n_3602)
);

OR2x6_ASAP7_75t_SL g3603 ( 
.A(n_3382),
.B(n_2946),
.Y(n_3603)
);

BUFx6f_ASAP7_75t_L g3604 ( 
.A(n_3269),
.Y(n_3604)
);

NAND2x1p5_ASAP7_75t_L g3605 ( 
.A(n_3433),
.B(n_2599),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3389),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3391),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3406),
.A2(n_2759),
.B(n_2679),
.Y(n_3608)
);

O2A1O1Ixp33_ASAP7_75t_L g3609 ( 
.A1(n_3254),
.A2(n_1180),
.B(n_3190),
.C(n_3184),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3379),
.B(n_2777),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3406),
.A2(n_2679),
.B(n_2674),
.Y(n_3611)
);

O2A1O1Ixp33_ASAP7_75t_L g3612 ( 
.A1(n_3255),
.A2(n_3261),
.B(n_3262),
.C(n_3260),
.Y(n_3612)
);

BUFx8_ASAP7_75t_L g3613 ( 
.A(n_3329),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_SL g3614 ( 
.A(n_3424),
.B(n_2605),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3295),
.B(n_602),
.Y(n_3615)
);

AND2x2_ASAP7_75t_SL g3616 ( 
.A(n_3427),
.B(n_2605),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_SL g3617 ( 
.A(n_3318),
.B(n_2634),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3424),
.B(n_602),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3418),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3422),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3263),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_R g3622 ( 
.A(n_3417),
.B(n_2605),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3441),
.B(n_2634),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3414),
.A2(n_2890),
.B(n_2888),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3287),
.A2(n_2890),
.B(n_2888),
.Y(n_3625)
);

O2A1O1Ixp33_ASAP7_75t_L g3626 ( 
.A1(n_3265),
.A2(n_3208),
.B(n_3204),
.C(n_3213),
.Y(n_3626)
);

BUFx2_ASAP7_75t_L g3627 ( 
.A(n_3274),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_SL g3628 ( 
.A(n_3433),
.B(n_2641),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3379),
.B(n_2789),
.Y(n_3629)
);

O2A1O1Ixp33_ASAP7_75t_SL g3630 ( 
.A1(n_3298),
.A2(n_3232),
.B(n_3162),
.C(n_3185),
.Y(n_3630)
);

CKINVDCx8_ASAP7_75t_R g3631 ( 
.A(n_3405),
.Y(n_3631)
);

CKINVDCx5p33_ASAP7_75t_R g3632 ( 
.A(n_3275),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3431),
.B(n_609),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_L g3634 ( 
.A(n_3432),
.B(n_611),
.Y(n_3634)
);

O2A1O1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3299),
.A2(n_3227),
.B(n_3215),
.C(n_3210),
.Y(n_3635)
);

CKINVDCx20_ASAP7_75t_R g3636 ( 
.A(n_3302),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_L g3637 ( 
.A(n_3373),
.B(n_3375),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3305),
.Y(n_3638)
);

INVx2_ASAP7_75t_SL g3639 ( 
.A(n_3409),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3407),
.B(n_3411),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_3425),
.B(n_611),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3427),
.A2(n_2835),
.B1(n_2703),
.B2(n_2743),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_3311),
.A2(n_3188),
.B1(n_3203),
.B2(n_3178),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3287),
.A2(n_2894),
.B(n_2816),
.Y(n_3644)
);

BUFx4f_ASAP7_75t_L g3645 ( 
.A(n_3409),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3430),
.B(n_3366),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3313),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3366),
.B(n_861),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3367),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3359),
.A2(n_2894),
.B(n_2816),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_3367),
.B(n_2641),
.Y(n_3651)
);

OAI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3461),
.A2(n_2631),
.B(n_2628),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3613),
.Y(n_3653)
);

INVx5_ASAP7_75t_L g3654 ( 
.A(n_3450),
.Y(n_3654)
);

CKINVDCx6p67_ASAP7_75t_R g3655 ( 
.A(n_3448),
.Y(n_3655)
);

AOI222xp33_ASAP7_75t_L g3656 ( 
.A1(n_3517),
.A2(n_851),
.B1(n_822),
.B2(n_819),
.C1(n_816),
.C2(n_820),
.Y(n_3656)
);

NOR2xp67_ASAP7_75t_L g3657 ( 
.A(n_3586),
.B(n_3516),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_SL g3658 ( 
.A(n_3454),
.B(n_3267),
.Y(n_3658)
);

INVx3_ASAP7_75t_L g3659 ( 
.A(n_3450),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3458),
.Y(n_3660)
);

AOI21xp33_ASAP7_75t_L g3661 ( 
.A1(n_3446),
.A2(n_3323),
.B(n_3321),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3462),
.Y(n_3662)
);

AOI222xp33_ASAP7_75t_SL g3663 ( 
.A1(n_3568),
.A2(n_3331),
.B1(n_3324),
.B2(n_832),
.C1(n_818),
.C2(n_839),
.Y(n_3663)
);

INVxp67_ASAP7_75t_SL g3664 ( 
.A(n_3499),
.Y(n_3664)
);

BUFx6f_ASAP7_75t_L g3665 ( 
.A(n_3645),
.Y(n_3665)
);

OAI22x1_ASAP7_75t_L g3666 ( 
.A1(n_3457),
.A2(n_3397),
.B1(n_3434),
.B2(n_3276),
.Y(n_3666)
);

INVx4_ASAP7_75t_L g3667 ( 
.A(n_3450),
.Y(n_3667)
);

BUFx2_ASAP7_75t_L g3668 ( 
.A(n_3528),
.Y(n_3668)
);

INVx5_ASAP7_75t_L g3669 ( 
.A(n_3570),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3479),
.B(n_3397),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3449),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3466),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_3613),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3463),
.B(n_3434),
.Y(n_3674)
);

BUFx3_ASAP7_75t_L g3675 ( 
.A(n_3595),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_3496),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3476),
.Y(n_3677)
);

OAI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3482),
.A2(n_3316),
.B1(n_3392),
.B2(n_3390),
.Y(n_3678)
);

INVx4_ASAP7_75t_L g3679 ( 
.A(n_3570),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3484),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3459),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3474),
.B(n_3247),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3538),
.B(n_3316),
.Y(n_3683)
);

A2O1A1Ixp33_ASAP7_75t_L g3684 ( 
.A1(n_3488),
.A2(n_3304),
.B(n_2631),
.C(n_3130),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3452),
.B(n_3409),
.Y(n_3685)
);

AOI22xp33_ASAP7_75t_L g3686 ( 
.A1(n_3447),
.A2(n_2703),
.B1(n_2743),
.B2(n_2717),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3469),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3531),
.B(n_3247),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3513),
.B(n_3247),
.Y(n_3689)
);

CKINVDCx11_ASAP7_75t_R g3690 ( 
.A(n_3603),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3494),
.Y(n_3691)
);

BUFx2_ASAP7_75t_L g3692 ( 
.A(n_3524),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3497),
.Y(n_3693)
);

BUFx4f_ASAP7_75t_SL g3694 ( 
.A(n_3580),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_3472),
.Y(n_3695)
);

CKINVDCx20_ASAP7_75t_R g3696 ( 
.A(n_3547),
.Y(n_3696)
);

O2A1O1Ixp33_ASAP7_75t_SL g3697 ( 
.A1(n_3565),
.A2(n_3223),
.B(n_3225),
.C(n_3220),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_R g3698 ( 
.A(n_3631),
.B(n_3632),
.Y(n_3698)
);

AND2x4_ASAP7_75t_L g3699 ( 
.A(n_3538),
.B(n_3267),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3456),
.B(n_3256),
.Y(n_3700)
);

AOI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3504),
.A2(n_824),
.B1(n_840),
.B2(n_811),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3636),
.A2(n_845),
.B1(n_849),
.B2(n_844),
.Y(n_3702)
);

BUFx6f_ASAP7_75t_L g3703 ( 
.A(n_3645),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3563),
.B(n_3256),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3560),
.B(n_3256),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3475),
.B(n_3266),
.Y(n_3706)
);

NAND2x1p5_ASAP7_75t_L g3707 ( 
.A(n_3519),
.B(n_3276),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3570),
.Y(n_3708)
);

BUFx6f_ASAP7_75t_L g3709 ( 
.A(n_3604),
.Y(n_3709)
);

INVx3_ASAP7_75t_L g3710 ( 
.A(n_3604),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3579),
.B(n_3618),
.Y(n_3711)
);

BUFx2_ASAP7_75t_L g3712 ( 
.A(n_3550),
.Y(n_3712)
);

OAI22x1_ASAP7_75t_L g3713 ( 
.A1(n_3530),
.A2(n_3377),
.B1(n_3355),
.B2(n_855),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3498),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3477),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3527),
.B(n_3266),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3557),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3529),
.B(n_3266),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_3544),
.B(n_861),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3481),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3486),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3501),
.B(n_3355),
.Y(n_3722)
);

INVx2_ASAP7_75t_SL g3723 ( 
.A(n_3534),
.Y(n_3723)
);

O2A1O1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_3615),
.A2(n_3230),
.B(n_3229),
.C(n_3130),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3541),
.B(n_3478),
.Y(n_3725)
);

INVx5_ASAP7_75t_L g3726 ( 
.A(n_3604),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3483),
.B(n_3325),
.Y(n_3727)
);

AND2x4_ASAP7_75t_L g3728 ( 
.A(n_3501),
.B(n_3377),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3562),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3559),
.B(n_3549),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3569),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3522),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3536),
.Y(n_3733)
);

A2O1A1Ixp33_ASAP7_75t_SL g3734 ( 
.A1(n_3468),
.A2(n_2054),
.B(n_2056),
.C(n_2027),
.Y(n_3734)
);

INVx4_ASAP7_75t_L g3735 ( 
.A(n_3519),
.Y(n_3735)
);

INVx4_ASAP7_75t_L g3736 ( 
.A(n_3589),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3512),
.B(n_3325),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3571),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3525),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3542),
.Y(n_3740)
);

CKINVDCx8_ASAP7_75t_R g3741 ( 
.A(n_3594),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3495),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3575),
.Y(n_3743)
);

INVx5_ASAP7_75t_L g3744 ( 
.A(n_3501),
.Y(n_3744)
);

BUFx2_ASAP7_75t_L g3745 ( 
.A(n_3523),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3577),
.Y(n_3746)
);

NAND2x1p5_ASAP7_75t_L g3747 ( 
.A(n_3589),
.B(n_3325),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3561),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3567),
.Y(n_3749)
);

BUFx2_ASAP7_75t_SL g3750 ( 
.A(n_3649),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3578),
.Y(n_3751)
);

BUFx2_ASAP7_75t_L g3752 ( 
.A(n_3622),
.Y(n_3752)
);

CKINVDCx6p67_ASAP7_75t_R g3753 ( 
.A(n_3532),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3597),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_SL g3755 ( 
.A(n_3473),
.B(n_3333),
.Y(n_3755)
);

INVx3_ASAP7_75t_L g3756 ( 
.A(n_3525),
.Y(n_3756)
);

HB1xp67_ASAP7_75t_L g3757 ( 
.A(n_3554),
.Y(n_3757)
);

BUFx6f_ASAP7_75t_L g3758 ( 
.A(n_3520),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3445),
.A2(n_2642),
.B(n_3176),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3465),
.B(n_863),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3583),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3518),
.A2(n_2703),
.B1(n_2743),
.B2(n_2717),
.Y(n_3762)
);

AO22x1_ASAP7_75t_L g3763 ( 
.A1(n_3648),
.A2(n_856),
.B1(n_857),
.B2(n_852),
.Y(n_3763)
);

AOI22xp33_ASAP7_75t_L g3764 ( 
.A1(n_3480),
.A2(n_2703),
.B1(n_2743),
.B2(n_2717),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3601),
.Y(n_3765)
);

HB1xp67_ASAP7_75t_L g3766 ( 
.A(n_3621),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3606),
.Y(n_3767)
);

INVx2_ASAP7_75t_SL g3768 ( 
.A(n_3548),
.Y(n_3768)
);

HB1xp67_ASAP7_75t_L g3769 ( 
.A(n_3638),
.Y(n_3769)
);

BUFx6f_ASAP7_75t_L g3770 ( 
.A(n_3520),
.Y(n_3770)
);

INVx1_ASAP7_75t_SL g3771 ( 
.A(n_3546),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3647),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3502),
.A2(n_2642),
.B(n_3176),
.Y(n_3773)
);

BUFx6f_ASAP7_75t_L g3774 ( 
.A(n_3515),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3566),
.B(n_3333),
.Y(n_3775)
);

HB1xp67_ASAP7_75t_L g3776 ( 
.A(n_3646),
.Y(n_3776)
);

AND2x4_ASAP7_75t_L g3777 ( 
.A(n_3509),
.B(n_3333),
.Y(n_3777)
);

OR2x6_ASAP7_75t_L g3778 ( 
.A(n_3509),
.B(n_3341),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3467),
.A2(n_2628),
.B(n_2901),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3485),
.B(n_3341),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3640),
.B(n_3341),
.Y(n_3781)
);

OAI22xp5_ASAP7_75t_SL g3782 ( 
.A1(n_3582),
.A2(n_859),
.B1(n_858),
.B2(n_863),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_SL g3783 ( 
.A1(n_3540),
.A2(n_3198),
.B(n_2809),
.Y(n_3783)
);

BUFx12f_ASAP7_75t_L g3784 ( 
.A(n_3535),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3505),
.B(n_3342),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3470),
.A2(n_2906),
.B(n_2901),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3607),
.Y(n_3787)
);

CKINVDCx20_ASAP7_75t_R g3788 ( 
.A(n_3627),
.Y(n_3788)
);

CKINVDCx8_ASAP7_75t_R g3789 ( 
.A(n_3512),
.Y(n_3789)
);

BUFx10_ASAP7_75t_L g3790 ( 
.A(n_3510),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3619),
.Y(n_3791)
);

OR2x6_ASAP7_75t_L g3792 ( 
.A(n_3509),
.B(n_3342),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3620),
.Y(n_3793)
);

HB1xp67_ASAP7_75t_L g3794 ( 
.A(n_3637),
.Y(n_3794)
);

NOR2x1_ASAP7_75t_L g3795 ( 
.A(n_3585),
.B(n_3342),
.Y(n_3795)
);

INVx5_ASAP7_75t_L g3796 ( 
.A(n_3585),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3507),
.B(n_2587),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3612),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3587),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3464),
.Y(n_3800)
);

OR2x6_ASAP7_75t_L g3801 ( 
.A(n_3585),
.B(n_2798),
.Y(n_3801)
);

INVx1_ASAP7_75t_SL g3802 ( 
.A(n_3514),
.Y(n_3802)
);

OR2x2_ASAP7_75t_L g3803 ( 
.A(n_3588),
.B(n_2906),
.Y(n_3803)
);

BUFx2_ASAP7_75t_SL g3804 ( 
.A(n_3623),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3598),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3444),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_3514),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3552),
.A2(n_2814),
.B1(n_2810),
.B2(n_2775),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3643),
.Y(n_3809)
);

NOR2xp33_ASAP7_75t_L g3810 ( 
.A(n_3471),
.B(n_867),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3487),
.Y(n_3811)
);

INVx4_ASAP7_75t_L g3812 ( 
.A(n_3564),
.Y(n_3812)
);

INVxp67_ASAP7_75t_SL g3813 ( 
.A(n_3581),
.Y(n_3813)
);

INVx5_ASAP7_75t_L g3814 ( 
.A(n_3564),
.Y(n_3814)
);

OAI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3553),
.A2(n_3128),
.B1(n_2803),
.B2(n_2809),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3630),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3616),
.Y(n_3817)
);

INVx4_ASAP7_75t_L g3818 ( 
.A(n_3503),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3614),
.Y(n_3819)
);

BUFx2_ASAP7_75t_L g3820 ( 
.A(n_3451),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3599),
.B(n_867),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3521),
.A2(n_3128),
.B1(n_2803),
.B2(n_2520),
.Y(n_3822)
);

CKINVDCx16_ASAP7_75t_R g3823 ( 
.A(n_3617),
.Y(n_3823)
);

BUFx6f_ASAP7_75t_L g3824 ( 
.A(n_3451),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3455),
.B(n_2591),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3610),
.B(n_2594),
.Y(n_3826)
);

BUFx6f_ASAP7_75t_L g3827 ( 
.A(n_3639),
.Y(n_3827)
);

CKINVDCx16_ASAP7_75t_R g3828 ( 
.A(n_3617),
.Y(n_3828)
);

NOR2xp67_ASAP7_75t_SL g3829 ( 
.A(n_3490),
.B(n_3573),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3599),
.B(n_872),
.Y(n_3830)
);

INVx3_ASAP7_75t_L g3831 ( 
.A(n_3487),
.Y(n_3831)
);

CKINVDCx20_ASAP7_75t_R g3832 ( 
.A(n_3506),
.Y(n_3832)
);

INVx3_ASAP7_75t_L g3833 ( 
.A(n_3508),
.Y(n_3833)
);

BUFx2_ASAP7_75t_L g3834 ( 
.A(n_3460),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3460),
.Y(n_3835)
);

BUFx4f_ASAP7_75t_L g3836 ( 
.A(n_3623),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3508),
.Y(n_3837)
);

INVx1_ASAP7_75t_SL g3838 ( 
.A(n_3629),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3651),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3602),
.B(n_2595),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3493),
.B(n_2602),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3489),
.A2(n_2738),
.B(n_2813),
.Y(n_3842)
);

AND2x4_ASAP7_75t_L g3843 ( 
.A(n_3555),
.B(n_2603),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3593),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3574),
.A2(n_2863),
.B1(n_2907),
.B2(n_2830),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3596),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3526),
.B(n_2607),
.Y(n_3847)
);

INVx3_ASAP7_75t_L g3848 ( 
.A(n_3605),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3551),
.Y(n_3849)
);

BUFx2_ASAP7_75t_L g3850 ( 
.A(n_3500),
.Y(n_3850)
);

OAI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3453),
.A2(n_2863),
.B1(n_2907),
.B2(n_2830),
.Y(n_3851)
);

CKINVDCx5p33_ASAP7_75t_R g3852 ( 
.A(n_3633),
.Y(n_3852)
);

OR2x2_ASAP7_75t_L g3853 ( 
.A(n_3491),
.B(n_2765),
.Y(n_3853)
);

BUFx6f_ASAP7_75t_L g3854 ( 
.A(n_3634),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3641),
.Y(n_3855)
);

AND2x4_ASAP7_75t_L g3856 ( 
.A(n_3624),
.B(n_2773),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3591),
.B(n_3492),
.Y(n_3857)
);

BUFx10_ASAP7_75t_L g3858 ( 
.A(n_3628),
.Y(n_3858)
);

INVx1_ASAP7_75t_SL g3859 ( 
.A(n_3628),
.Y(n_3859)
);

BUFx12f_ASAP7_75t_L g3860 ( 
.A(n_3576),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3492),
.B(n_2778),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3600),
.Y(n_3862)
);

INVx5_ASAP7_75t_L g3863 ( 
.A(n_3858),
.Y(n_3863)
);

BUFx2_ASAP7_75t_SL g3864 ( 
.A(n_3788),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_3852),
.B(n_872),
.Y(n_3865)
);

NAND3x1_ASAP7_75t_L g3866 ( 
.A(n_3674),
.B(n_3511),
.C(n_3533),
.Y(n_3866)
);

OAI22x1_ASAP7_75t_L g3867 ( 
.A1(n_3862),
.A2(n_902),
.B1(n_907),
.B2(n_886),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3725),
.B(n_3545),
.Y(n_3868)
);

O2A1O1Ixp33_ASAP7_75t_SL g3869 ( 
.A1(n_3810),
.A2(n_3543),
.B(n_3626),
.C(n_3609),
.Y(n_3869)
);

A2O1A1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_3821),
.A2(n_3584),
.B(n_3572),
.C(n_3635),
.Y(n_3870)
);

AO21x1_ASAP7_75t_L g3871 ( 
.A1(n_3800),
.A2(n_3558),
.B(n_3556),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3760),
.A2(n_3539),
.B(n_3590),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3766),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3689),
.B(n_3642),
.Y(n_3874)
);

A2O1A1Ixp33_ASAP7_75t_L g3875 ( 
.A1(n_3830),
.A2(n_3608),
.B(n_3537),
.C(n_3592),
.Y(n_3875)
);

A2O1A1Ixp33_ASAP7_75t_L g3876 ( 
.A1(n_3701),
.A2(n_3625),
.B(n_3650),
.C(n_3644),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3773),
.A2(n_3611),
.B(n_2881),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3704),
.B(n_4),
.Y(n_3878)
);

NAND3xp33_ASAP7_75t_SL g3879 ( 
.A(n_3656),
.B(n_902),
.C(n_886),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3769),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3786),
.A2(n_2881),
.B(n_2874),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3779),
.A2(n_2897),
.B(n_2874),
.Y(n_3882)
);

BUFx12f_ASAP7_75t_L g3883 ( 
.A(n_3695),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3759),
.A2(n_2897),
.B(n_2813),
.Y(n_3884)
);

O2A1O1Ixp33_ASAP7_75t_SL g3885 ( 
.A1(n_3755),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_3885)
);

BUFx3_ASAP7_75t_L g3886 ( 
.A(n_3696),
.Y(n_3886)
);

OAI21x1_ASAP7_75t_L g3887 ( 
.A1(n_3842),
.A2(n_2738),
.B(n_2781),
.Y(n_3887)
);

INVx3_ASAP7_75t_L g3888 ( 
.A(n_3831),
.Y(n_3888)
);

OAI22x1_ASAP7_75t_L g3889 ( 
.A1(n_3776),
.A2(n_921),
.B1(n_925),
.B2(n_907),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3772),
.Y(n_3890)
);

BUFx6f_ASAP7_75t_L g3891 ( 
.A(n_3665),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3660),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3652),
.A2(n_2669),
.B(n_2663),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3662),
.Y(n_3894)
);

BUFx3_ASAP7_75t_L g3895 ( 
.A(n_3655),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3697),
.A2(n_2669),
.B(n_2663),
.Y(n_3896)
);

O2A1O1Ixp33_ASAP7_75t_SL g3897 ( 
.A1(n_3859),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_3897)
);

OA21x2_ASAP7_75t_L g3898 ( 
.A1(n_3857),
.A2(n_2792),
.B(n_2791),
.Y(n_3898)
);

INVx5_ASAP7_75t_L g3899 ( 
.A(n_3858),
.Y(n_3899)
);

CKINVDCx5p33_ASAP7_75t_R g3900 ( 
.A(n_3694),
.Y(n_3900)
);

BUFx3_ASAP7_75t_L g3901 ( 
.A(n_3784),
.Y(n_3901)
);

NOR2xp33_ASAP7_75t_SL g3902 ( 
.A(n_3741),
.B(n_921),
.Y(n_3902)
);

OAI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3823),
.A2(n_2802),
.B1(n_2806),
.B2(n_2801),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3828),
.A2(n_2846),
.B1(n_2849),
.B2(n_2831),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3672),
.Y(n_3905)
);

AND2x4_ASAP7_75t_L g3906 ( 
.A(n_3744),
.B(n_2858),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3825),
.A2(n_2696),
.B(n_2669),
.Y(n_3907)
);

OAI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3657),
.A2(n_3855),
.B1(n_3854),
.B2(n_3832),
.Y(n_3908)
);

OAI21xp33_ASAP7_75t_L g3909 ( 
.A1(n_3849),
.A2(n_931),
.B(n_925),
.Y(n_3909)
);

OAI21x1_ASAP7_75t_L g3910 ( 
.A1(n_3816),
.A2(n_2866),
.B(n_2864),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3663),
.A2(n_932),
.B1(n_933),
.B2(n_931),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3744),
.B(n_2868),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3687),
.Y(n_3913)
);

CKINVDCx11_ASAP7_75t_R g3914 ( 
.A(n_3690),
.Y(n_3914)
);

O2A1O1Ixp33_ASAP7_75t_L g3915 ( 
.A1(n_3844),
.A2(n_2878),
.B(n_2879),
.C(n_2871),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3730),
.B(n_932),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3691),
.Y(n_3917)
);

O2A1O1Ixp33_ASAP7_75t_SL g3918 ( 
.A1(n_3794),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3847),
.A2(n_2732),
.B(n_2696),
.Y(n_3919)
);

BUFx2_ASAP7_75t_L g3920 ( 
.A(n_3668),
.Y(n_3920)
);

INVx3_ASAP7_75t_L g3921 ( 
.A(n_3831),
.Y(n_3921)
);

AO31x2_ASAP7_75t_L g3922 ( 
.A1(n_3666),
.A2(n_2886),
.A3(n_2896),
.B(n_2884),
.Y(n_3922)
);

INVx3_ASAP7_75t_L g3923 ( 
.A(n_3833),
.Y(n_3923)
);

NAND3xp33_ASAP7_75t_SL g3924 ( 
.A(n_3719),
.B(n_935),
.C(n_933),
.Y(n_3924)
);

O2A1O1Ixp33_ASAP7_75t_SL g3925 ( 
.A1(n_3661),
.A2(n_15),
.B(n_11),
.C(n_13),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3838),
.B(n_935),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3693),
.Y(n_3927)
);

OAI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3854),
.A2(n_944),
.B1(n_951),
.B2(n_937),
.Y(n_3928)
);

O2A1O1Ixp33_ASAP7_75t_L g3929 ( 
.A1(n_3678),
.A2(n_2904),
.B(n_2909),
.C(n_2902),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3854),
.A2(n_2814),
.B1(n_2810),
.B2(n_2775),
.Y(n_3930)
);

A2O1A1Ixp33_ASAP7_75t_L g3931 ( 
.A1(n_3806),
.A2(n_3840),
.B(n_3798),
.C(n_3808),
.Y(n_3931)
);

HB1xp67_ASAP7_75t_L g3932 ( 
.A(n_3757),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3799),
.B(n_937),
.Y(n_3933)
);

O2A1O1Ixp33_ASAP7_75t_L g3934 ( 
.A1(n_3734),
.A2(n_2910),
.B(n_2800),
.C(n_2804),
.Y(n_3934)
);

O2A1O1Ixp33_ASAP7_75t_L g3935 ( 
.A1(n_3840),
.A2(n_2805),
.B(n_2815),
.C(n_2799),
.Y(n_3935)
);

NOR2xp67_ASAP7_75t_SL g3936 ( 
.A(n_3744),
.B(n_2696),
.Y(n_3936)
);

O2A1O1Ixp33_ASAP7_75t_L g3937 ( 
.A1(n_3853),
.A2(n_2828),
.B(n_2838),
.C(n_2824),
.Y(n_3937)
);

OAI22xp5_ASAP7_75t_L g3938 ( 
.A1(n_3771),
.A2(n_3752),
.B1(n_3712),
.B2(n_3817),
.Y(n_3938)
);

O2A1O1Ixp33_ASAP7_75t_SL g3939 ( 
.A1(n_3700),
.A2(n_16),
.B(n_13),
.C(n_15),
.Y(n_3939)
);

A2O1A1Ixp33_ASAP7_75t_L g3940 ( 
.A1(n_3809),
.A2(n_951),
.B(n_955),
.C(n_944),
.Y(n_3940)
);

A2O1A1Ixp33_ASAP7_75t_L g3941 ( 
.A1(n_3686),
.A2(n_964),
.B(n_955),
.C(n_2840),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3805),
.B(n_964),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3711),
.B(n_3692),
.Y(n_3943)
);

O2A1O1Ixp33_ASAP7_75t_SL g3944 ( 
.A1(n_3768),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3782),
.A2(n_2814),
.B1(n_2810),
.B2(n_2775),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3714),
.Y(n_3946)
);

INVx1_ASAP7_75t_SL g3947 ( 
.A(n_3680),
.Y(n_3947)
);

AOI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3684),
.A2(n_2736),
.B(n_2732),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3822),
.A2(n_2736),
.B(n_2732),
.Y(n_3949)
);

CKINVDCx5p33_ASAP7_75t_R g3950 ( 
.A(n_3676),
.Y(n_3950)
);

BUFx12f_ASAP7_75t_L g3951 ( 
.A(n_3790),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3665),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3717),
.Y(n_3953)
);

AOI221x1_ASAP7_75t_L g3954 ( 
.A1(n_3713),
.A2(n_1544),
.B1(n_1546),
.B2(n_1545),
.C(n_1535),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3742),
.Y(n_3955)
);

A2O1A1Ixp33_ASAP7_75t_L g3956 ( 
.A1(n_3813),
.A2(n_2844),
.B(n_2851),
.C(n_2842),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3664),
.B(n_1545),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3670),
.A2(n_2742),
.B(n_2736),
.Y(n_3958)
);

O2A1O1Ixp33_ASAP7_75t_SL g3959 ( 
.A1(n_3819),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_3959)
);

A2O1A1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3829),
.A2(n_2875),
.B(n_2869),
.C(n_2748),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3834),
.B(n_19),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3775),
.B(n_1546),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3841),
.A2(n_2748),
.B(n_2742),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3801),
.A2(n_3789),
.B1(n_3796),
.B2(n_3702),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3729),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3731),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_SL g3967 ( 
.A(n_3658),
.B(n_3099),
.Y(n_3967)
);

OAI21xp33_ASAP7_75t_L g3968 ( 
.A1(n_3846),
.A2(n_1548),
.B(n_1547),
.Y(n_3968)
);

AOI221xp5_ASAP7_75t_SL g3969 ( 
.A1(n_3780),
.A2(n_1586),
.B1(n_1588),
.B2(n_1575),
.C(n_1573),
.Y(n_3969)
);

BUFx10_ASAP7_75t_L g3970 ( 
.A(n_3665),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3738),
.Y(n_3971)
);

OAI21x1_ASAP7_75t_L g3972 ( 
.A1(n_3783),
.A2(n_1548),
.B(n_1547),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_L g3973 ( 
.A1(n_3835),
.A2(n_2814),
.B1(n_2810),
.B2(n_2775),
.Y(n_3973)
);

AOI21x1_ASAP7_75t_L g3974 ( 
.A1(n_3829),
.A2(n_3861),
.B(n_3850),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3835),
.A2(n_2783),
.B1(n_2636),
.B2(n_2638),
.Y(n_3975)
);

INVx4_ASAP7_75t_L g3976 ( 
.A(n_3654),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3843),
.A2(n_2748),
.B(n_2742),
.Y(n_3977)
);

BUFx4f_ASAP7_75t_SL g3978 ( 
.A(n_3753),
.Y(n_3978)
);

AOI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3835),
.A2(n_2783),
.B1(n_2636),
.B2(n_2638),
.Y(n_3979)
);

AOI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3843),
.A2(n_2793),
.B(n_2774),
.Y(n_3980)
);

O2A1O1Ixp33_ASAP7_75t_SL g3981 ( 
.A1(n_3706),
.A2(n_23),
.B(n_20),
.C(n_22),
.Y(n_3981)
);

AOI22xp5_ASAP7_75t_L g3982 ( 
.A1(n_3763),
.A2(n_3099),
.B1(n_3148),
.B2(n_2783),
.Y(n_3982)
);

O2A1O1Ixp33_ASAP7_75t_SL g3983 ( 
.A1(n_3723),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3983)
);

NAND3xp33_ASAP7_75t_L g3984 ( 
.A(n_3797),
.B(n_1575),
.C(n_1573),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_SL g3985 ( 
.A(n_3796),
.B(n_3790),
.Y(n_3985)
);

INVx6_ASAP7_75t_L g3986 ( 
.A(n_3703),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3743),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3856),
.A2(n_2793),
.B(n_2774),
.Y(n_3988)
);

INVx2_ASAP7_75t_SL g3989 ( 
.A(n_3681),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3785),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3737),
.B(n_25),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3796),
.A2(n_2783),
.B1(n_2636),
.B2(n_2638),
.Y(n_3992)
);

OAI22x1_ASAP7_75t_L g3993 ( 
.A1(n_3745),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_3993)
);

OA21x2_ASAP7_75t_L g3994 ( 
.A1(n_3762),
.A2(n_2636),
.B(n_2638),
.Y(n_3994)
);

INVx3_ASAP7_75t_SL g3995 ( 
.A(n_3774),
.Y(n_3995)
);

A2O1A1Ixp33_ASAP7_75t_L g3996 ( 
.A1(n_3724),
.A2(n_2793),
.B(n_2796),
.C(n_2774),
.Y(n_3996)
);

CKINVDCx20_ASAP7_75t_R g3997 ( 
.A(n_3698),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3833),
.Y(n_3998)
);

AOI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3683),
.A2(n_3099),
.B1(n_3148),
.B2(n_1575),
.Y(n_3999)
);

BUFx6f_ASAP7_75t_L g4000 ( 
.A(n_3703),
.Y(n_4000)
);

NOR2x1_ASAP7_75t_R g4001 ( 
.A(n_3653),
.B(n_2796),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3688),
.B(n_1573),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3801),
.A2(n_3836),
.B1(n_3683),
.B2(n_3795),
.Y(n_4003)
);

INVx3_ASAP7_75t_L g4004 ( 
.A(n_3709),
.Y(n_4004)
);

BUFx8_ASAP7_75t_L g4005 ( 
.A(n_3703),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3860),
.A2(n_3099),
.B1(n_3148),
.B2(n_1575),
.Y(n_4006)
);

AO32x2_ASAP7_75t_L g4007 ( 
.A1(n_3851),
.A2(n_28),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_4007)
);

OAI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3739),
.A2(n_2811),
.B1(n_2825),
.B2(n_2796),
.Y(n_4008)
);

AOI22xp33_ASAP7_75t_L g4009 ( 
.A1(n_3739),
.A2(n_3148),
.B1(n_1573),
.B2(n_1588),
.Y(n_4009)
);

AOI211x1_ASAP7_75t_L g4010 ( 
.A1(n_3682),
.A2(n_3705),
.B(n_3727),
.C(n_3718),
.Y(n_4010)
);

NAND2x1_ASAP7_75t_L g4011 ( 
.A(n_3856),
.B(n_2507),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3746),
.Y(n_4012)
);

NOR2xp33_ASAP7_75t_L g4013 ( 
.A(n_3685),
.B(n_31),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3751),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3815),
.A2(n_2825),
.B(n_2811),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3778),
.A2(n_2825),
.B(n_2811),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3824),
.B(n_3758),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3716),
.B(n_1586),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3671),
.B(n_1586),
.Y(n_4019)
);

INVx3_ASAP7_75t_L g4020 ( 
.A(n_3709),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3764),
.A2(n_2856),
.B1(n_2861),
.B2(n_2854),
.Y(n_4021)
);

INVx2_ASAP7_75t_SL g4022 ( 
.A(n_3774),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3778),
.A2(n_2856),
.B(n_2854),
.Y(n_4023)
);

AOI21xp33_ASAP7_75t_L g4024 ( 
.A1(n_3803),
.A2(n_1588),
.B(n_1586),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3754),
.Y(n_4025)
);

OAI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3839),
.A2(n_2507),
.B(n_2837),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3781),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3750),
.Y(n_4028)
);

OAI22x1_ASAP7_75t_L g4029 ( 
.A1(n_3820),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_4029)
);

O2A1O1Ixp33_ASAP7_75t_L g4030 ( 
.A1(n_3826),
.A2(n_1529),
.B(n_2054),
.C(n_2027),
.Y(n_4030)
);

INVx3_ASAP7_75t_L g4031 ( 
.A(n_3709),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3677),
.B(n_1588),
.Y(n_4032)
);

AO22x1_ASAP7_75t_L g4033 ( 
.A1(n_3673),
.A2(n_44),
.B1(n_33),
.B2(n_37),
.Y(n_4033)
);

BUFx12f_ASAP7_75t_L g4034 ( 
.A(n_3774),
.Y(n_4034)
);

A2O1A1Ixp33_ASAP7_75t_L g4035 ( 
.A1(n_3750),
.A2(n_2856),
.B(n_2861),
.C(n_2854),
.Y(n_4035)
);

O2A1O1Ixp33_ASAP7_75t_L g4036 ( 
.A1(n_3845),
.A2(n_1529),
.B(n_2056),
.C(n_2054),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_3675),
.Y(n_4037)
);

O2A1O1Ixp33_ASAP7_75t_L g4038 ( 
.A1(n_3802),
.A2(n_1529),
.B(n_2064),
.C(n_2056),
.Y(n_4038)
);

CKINVDCx5p33_ASAP7_75t_R g4039 ( 
.A(n_3807),
.Y(n_4039)
);

OAI22xp5_ASAP7_75t_L g4040 ( 
.A1(n_3756),
.A2(n_2911),
.B1(n_2861),
.B2(n_1594),
.Y(n_4040)
);

AOI22xp33_ASAP7_75t_L g4041 ( 
.A1(n_3756),
.A2(n_1594),
.B1(n_1602),
.B2(n_1599),
.Y(n_4041)
);

O2A1O1Ixp33_ASAP7_75t_SL g4042 ( 
.A1(n_3848),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_4042)
);

AO32x2_ASAP7_75t_L g4043 ( 
.A1(n_3812),
.A2(n_3667),
.A3(n_3679),
.B1(n_3736),
.B2(n_3735),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_L g4044 ( 
.A1(n_3811),
.A2(n_2065),
.B(n_2064),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_L g4045 ( 
.A(n_3758),
.B(n_45),
.Y(n_4045)
);

CKINVDCx20_ASAP7_75t_R g4046 ( 
.A(n_3758),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3715),
.Y(n_4047)
);

AO31x2_ASAP7_75t_L g4048 ( 
.A1(n_3837),
.A2(n_2895),
.A3(n_2873),
.B(n_2837),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3720),
.Y(n_4049)
);

OAI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3707),
.A2(n_2507),
.B(n_2837),
.Y(n_4050)
);

OAI22x1_ASAP7_75t_L g4051 ( 
.A1(n_3721),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_4051)
);

BUFx10_ASAP7_75t_L g4052 ( 
.A(n_3827),
.Y(n_4052)
);

OAI21x1_ASAP7_75t_SL g4053 ( 
.A1(n_3735),
.A2(n_48),
.B(n_49),
.Y(n_4053)
);

O2A1O1Ixp33_ASAP7_75t_SL g4054 ( 
.A1(n_3848),
.A2(n_56),
.B(n_52),
.C(n_55),
.Y(n_4054)
);

OAI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3732),
.A2(n_2855),
.B(n_2837),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3733),
.B(n_55),
.Y(n_4056)
);

NAND2x1p5_ASAP7_75t_L g4057 ( 
.A(n_3654),
.B(n_2911),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3740),
.B(n_3748),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3749),
.B(n_1594),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3761),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3765),
.B(n_1594),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3767),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3787),
.B(n_1599),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3791),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3793),
.Y(n_4065)
);

OR2x2_ASAP7_75t_L g4066 ( 
.A(n_3804),
.B(n_1599),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_L g4067 ( 
.A1(n_3747),
.A2(n_2065),
.B(n_2064),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3824),
.B(n_1599),
.Y(n_4068)
);

A2O1A1Ixp33_ASAP7_75t_L g4069 ( 
.A1(n_3722),
.A2(n_2911),
.B(n_1610),
.C(n_1618),
.Y(n_4069)
);

OAI21x1_ASAP7_75t_L g4070 ( 
.A1(n_3659),
.A2(n_2065),
.B(n_1691),
.Y(n_4070)
);

OR2x6_ASAP7_75t_L g4071 ( 
.A(n_3804),
.B(n_1602),
.Y(n_4071)
);

O2A1O1Ixp33_ASAP7_75t_L g4072 ( 
.A1(n_3792),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3699),
.B(n_62),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3824),
.Y(n_4074)
);

A2O1A1Ixp33_ASAP7_75t_L g4075 ( 
.A1(n_3722),
.A2(n_3728),
.B(n_3659),
.C(n_3710),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3905),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3990),
.B(n_3699),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3955),
.B(n_3770),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3932),
.B(n_3770),
.Y(n_4079)
);

AOI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3879),
.A2(n_3728),
.B1(n_3777),
.B2(n_3792),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_3872),
.A2(n_3770),
.B1(n_3777),
.B2(n_3812),
.Y(n_4081)
);

NOR2xp33_ASAP7_75t_L g4082 ( 
.A(n_3908),
.B(n_3827),
.Y(n_4082)
);

NAND2xp33_ASAP7_75t_L g4083 ( 
.A(n_3866),
.B(n_3654),
.Y(n_4083)
);

NOR2xp67_ASAP7_75t_SL g4084 ( 
.A(n_3951),
.B(n_3669),
.Y(n_4084)
);

OAI21x1_ASAP7_75t_L g4085 ( 
.A1(n_3974),
.A2(n_3710),
.B(n_3708),
.Y(n_4085)
);

OAI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3911),
.A2(n_3669),
.B1(n_3726),
.B2(n_3818),
.Y(n_4086)
);

INVx4_ASAP7_75t_L g4087 ( 
.A(n_3863),
.Y(n_4087)
);

AOI221xp5_ASAP7_75t_L g4088 ( 
.A1(n_3918),
.A2(n_1610),
.B1(n_1621),
.B2(n_1618),
.C(n_1602),
.Y(n_4088)
);

INVx6_ASAP7_75t_L g4089 ( 
.A(n_4005),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4027),
.B(n_3873),
.Y(n_4090)
);

OAI211xp5_ASAP7_75t_L g4091 ( 
.A1(n_4072),
.A2(n_3679),
.B(n_3667),
.C(n_3708),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_L g4092 ( 
.A(n_3943),
.B(n_3827),
.Y(n_4092)
);

OR2x6_ASAP7_75t_L g4093 ( 
.A(n_3864),
.B(n_3736),
.Y(n_4093)
);

AOI22xp33_ASAP7_75t_SL g4094 ( 
.A1(n_3964),
.A2(n_3899),
.B1(n_3863),
.B2(n_4013),
.Y(n_4094)
);

AND2x4_ASAP7_75t_L g4095 ( 
.A(n_4028),
.B(n_3880),
.Y(n_4095)
);

CKINVDCx20_ASAP7_75t_R g4096 ( 
.A(n_3997),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3890),
.Y(n_4097)
);

OAI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3982),
.A2(n_3726),
.B1(n_3669),
.B2(n_3818),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_3924),
.A2(n_1602),
.B1(n_1618),
.B2(n_1610),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3927),
.Y(n_4100)
);

AOI21xp33_ASAP7_75t_L g4101 ( 
.A1(n_3868),
.A2(n_3814),
.B(n_3726),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_3875),
.A2(n_3814),
.B(n_2895),
.Y(n_4102)
);

OAI21x1_ASAP7_75t_L g4103 ( 
.A1(n_3877),
.A2(n_3919),
.B(n_3948),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3946),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4012),
.Y(n_4105)
);

AOI222xp33_ASAP7_75t_L g4106 ( 
.A1(n_3993),
.A2(n_1625),
.B1(n_1618),
.B2(n_1630),
.C1(n_1621),
.C2(n_1610),
.Y(n_4106)
);

A2O1A1Ixp33_ASAP7_75t_L g4107 ( 
.A1(n_3870),
.A2(n_3814),
.B(n_68),
.C(n_65),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_3909),
.A2(n_3867),
.B1(n_3914),
.B2(n_3871),
.Y(n_4108)
);

INVx3_ASAP7_75t_L g4109 ( 
.A(n_3888),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_4010),
.A2(n_3931),
.B1(n_3945),
.B2(n_3899),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_3874),
.A2(n_1621),
.B1(n_1630),
.B2(n_1625),
.Y(n_4111)
);

AOI21xp33_ASAP7_75t_L g4112 ( 
.A1(n_3889),
.A2(n_1625),
.B(n_1621),
.Y(n_4112)
);

OAI211xp5_ASAP7_75t_L g4113 ( 
.A1(n_3897),
.A2(n_3983),
.B(n_3944),
.C(n_4042),
.Y(n_4113)
);

OAI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_3863),
.A2(n_1625),
.B1(n_1642),
.B2(n_1630),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3899),
.A2(n_1630),
.B1(n_1645),
.B2(n_1642),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3892),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_4014),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_3920),
.B(n_65),
.Y(n_4118)
);

BUFx2_ASAP7_75t_L g4119 ( 
.A(n_3888),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4025),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_3894),
.B(n_66),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_4053),
.A2(n_3985),
.B1(n_3938),
.B2(n_4045),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3865),
.A2(n_1642),
.B1(n_1649),
.B2(n_1645),
.Y(n_4123)
);

O2A1O1Ixp5_ASAP7_75t_L g4124 ( 
.A1(n_4033),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_4124)
);

BUFx6f_ASAP7_75t_L g4125 ( 
.A(n_3895),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_4029),
.A2(n_1642),
.B1(n_1649),
.B2(n_1645),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3913),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3917),
.Y(n_4128)
);

OAI211xp5_ASAP7_75t_L g4129 ( 
.A1(n_4054),
.A2(n_3925),
.B(n_3959),
.C(n_3981),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3953),
.Y(n_4130)
);

OR2x2_ASAP7_75t_L g4131 ( 
.A(n_3947),
.B(n_1645),
.Y(n_4131)
);

AOI22xp33_ASAP7_75t_L g4132 ( 
.A1(n_4051),
.A2(n_1649),
.B1(n_1561),
.B2(n_1532),
.Y(n_4132)
);

INVx1_ASAP7_75t_SL g4133 ( 
.A(n_3995),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3965),
.Y(n_4134)
);

INVx1_ASAP7_75t_SL g4135 ( 
.A(n_4039),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_3878),
.A2(n_1649),
.B1(n_1561),
.B2(n_1532),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3966),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3869),
.A2(n_2873),
.B(n_1561),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_3900),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3971),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_3876),
.A2(n_1561),
.B(n_1533),
.Y(n_4141)
);

OAI22xp5_ASAP7_75t_SL g4142 ( 
.A1(n_3978),
.A2(n_4046),
.B1(n_4037),
.B2(n_4034),
.Y(n_4142)
);

BUFx2_ASAP7_75t_L g4143 ( 
.A(n_3921),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4064),
.B(n_69),
.Y(n_4144)
);

AO221x2_ASAP7_75t_L g4145 ( 
.A1(n_4003),
.A2(n_4074),
.B1(n_3928),
.B2(n_4007),
.C(n_3987),
.Y(n_4145)
);

HB1xp67_ASAP7_75t_L g4146 ( 
.A(n_4047),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4049),
.Y(n_4147)
);

OAI22xp5_ASAP7_75t_L g4148 ( 
.A1(n_4006),
.A2(n_1561),
.B1(n_1533),
.B2(n_74),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_3901),
.A2(n_1533),
.B1(n_2570),
.B2(n_2855),
.Y(n_4149)
);

AOI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_4073),
.A2(n_1533),
.B1(n_2570),
.B2(n_2855),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4060),
.Y(n_4151)
);

CKINVDCx6p67_ASAP7_75t_R g4152 ( 
.A(n_3883),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4062),
.Y(n_4153)
);

BUFx6f_ASAP7_75t_L g4154 ( 
.A(n_3891),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4065),
.B(n_73),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_SL g4156 ( 
.A(n_4075),
.B(n_1482),
.Y(n_4156)
);

BUFx12f_ASAP7_75t_L g4157 ( 
.A(n_3950),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4058),
.Y(n_4158)
);

OAI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_3940),
.A2(n_77),
.B1(n_73),
.B2(n_76),
.Y(n_4159)
);

OAI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_3999),
.A2(n_82),
.B1(n_78),
.B2(n_80),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3957),
.Y(n_4161)
);

AOI22xp33_ASAP7_75t_L g4162 ( 
.A1(n_3991),
.A2(n_2570),
.B1(n_2880),
.B2(n_2855),
.Y(n_4162)
);

OAI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3967),
.A2(n_84),
.B1(n_78),
.B2(n_83),
.Y(n_4163)
);

HB1xp67_ASAP7_75t_L g4164 ( 
.A(n_3921),
.Y(n_4164)
);

O2A1O1Ixp33_ASAP7_75t_SL g4165 ( 
.A1(n_3916),
.A2(n_88),
.B(n_83),
.C(n_87),
.Y(n_4165)
);

OAI221xp5_ASAP7_75t_L g4166 ( 
.A1(n_3942),
.A2(n_91),
.B1(n_87),
.B2(n_88),
.C(n_92),
.Y(n_4166)
);

INVx3_ASAP7_75t_L g4167 ( 
.A(n_3923),
.Y(n_4167)
);

BUFx2_ASAP7_75t_L g4168 ( 
.A(n_3923),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3998),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_L g4170 ( 
.A1(n_3961),
.A2(n_2570),
.B1(n_2880),
.B2(n_1392),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_3898),
.B(n_91),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3922),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_3941),
.A2(n_97),
.B1(n_93),
.B2(n_96),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_3989),
.B(n_3886),
.Y(n_4174)
);

OAI22xp5_ASAP7_75t_L g4175 ( 
.A1(n_3992),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_4175)
);

INVx3_ASAP7_75t_SL g4176 ( 
.A(n_3986),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_3906),
.A2(n_2880),
.B1(n_1392),
.B2(n_1407),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_4022),
.B(n_100),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3922),
.Y(n_4179)
);

AND2x4_ASAP7_75t_L g4180 ( 
.A(n_4004),
.B(n_4020),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_3898),
.B(n_101),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_L g4182 ( 
.A1(n_3906),
.A2(n_2880),
.B1(n_1407),
.B2(n_1397),
.Y(n_4182)
);

INVx4_ASAP7_75t_L g4183 ( 
.A(n_3976),
.Y(n_4183)
);

INVx4_ASAP7_75t_L g4184 ( 
.A(n_3976),
.Y(n_4184)
);

OAI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_3954),
.A2(n_106),
.B1(n_102),
.B2(n_103),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3922),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4002),
.B(n_102),
.Y(n_4187)
);

AO21x2_ASAP7_75t_L g4188 ( 
.A1(n_3907),
.A2(n_3958),
.B(n_3996),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_SL g4189 ( 
.A(n_3902),
.B(n_1495),
.Y(n_4189)
);

NAND2xp33_ASAP7_75t_L g4190 ( 
.A(n_3891),
.B(n_1466),
.Y(n_4190)
);

CKINVDCx20_ASAP7_75t_R g4191 ( 
.A(n_4005),
.Y(n_4191)
);

INVx5_ASAP7_75t_L g4192 ( 
.A(n_4071),
.Y(n_4192)
);

INVx3_ASAP7_75t_L g4193 ( 
.A(n_4052),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_L g4194 ( 
.A1(n_3912),
.A2(n_3893),
.B1(n_3968),
.B2(n_3933),
.Y(n_4194)
);

OAI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_4011),
.A2(n_108),
.B1(n_103),
.B2(n_106),
.Y(n_4195)
);

AND2x4_ASAP7_75t_SL g4196 ( 
.A(n_3970),
.B(n_1466),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3962),
.B(n_108),
.Y(n_4197)
);

HB1xp67_ASAP7_75t_L g4198 ( 
.A(n_3994),
.Y(n_4198)
);

AO221x2_ASAP7_75t_L g4199 ( 
.A1(n_4007),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_4199)
);

BUFx6f_ASAP7_75t_L g4200 ( 
.A(n_3891),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4004),
.B(n_110),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_4018),
.B(n_111),
.Y(n_4202)
);

AND2x4_ASAP7_75t_L g4203 ( 
.A(n_4020),
.B(n_112),
.Y(n_4203)
);

INVxp67_ASAP7_75t_L g4204 ( 
.A(n_3926),
.Y(n_4204)
);

AND2x4_ASAP7_75t_L g4205 ( 
.A(n_4031),
.B(n_113),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4056),
.Y(n_4206)
);

OAI22xp33_ASAP7_75t_L g4207 ( 
.A1(n_4071),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4207)
);

CKINVDCx6p67_ASAP7_75t_R g4208 ( 
.A(n_3970),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4019),
.Y(n_4209)
);

OAI21x1_ASAP7_75t_L g4210 ( 
.A1(n_3910),
.A2(n_1694),
.B(n_1685),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_4031),
.B(n_114),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4043),
.Y(n_4212)
);

AOI22xp33_ASAP7_75t_L g4213 ( 
.A1(n_3912),
.A2(n_1407),
.B1(n_1397),
.B2(n_1368),
.Y(n_4213)
);

AOI21x1_ASAP7_75t_L g4214 ( 
.A1(n_3896),
.A2(n_115),
.B(n_116),
.Y(n_4214)
);

AOI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_3994),
.A2(n_1397),
.B1(n_1412),
.B2(n_1368),
.Y(n_4215)
);

CKINVDCx11_ASAP7_75t_R g4216 ( 
.A(n_4052),
.Y(n_4216)
);

AOI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_3885),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_4217)
);

INVxp67_ASAP7_75t_L g4218 ( 
.A(n_4017),
.Y(n_4218)
);

OAI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_3949),
.A2(n_123),
.B1(n_117),
.B2(n_120),
.Y(n_4219)
);

CKINVDCx5p33_ASAP7_75t_R g4220 ( 
.A(n_3952),
.Y(n_4220)
);

AOI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_3939),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4032),
.Y(n_4222)
);

OAI22xp33_ASAP7_75t_L g4223 ( 
.A1(n_4026),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4059),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_3952),
.B(n_127),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3963),
.B(n_128),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_3952),
.B(n_129),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4061),
.Y(n_4228)
);

OAI22xp5_ASAP7_75t_L g4229 ( 
.A1(n_3930),
.A2(n_140),
.B1(n_130),
.B2(n_134),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4000),
.B(n_130),
.Y(n_4230)
);

CKINVDCx14_ASAP7_75t_R g4231 ( 
.A(n_3986),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4007),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_4043),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4063),
.B(n_140),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4043),
.Y(n_4235)
);

CKINVDCx5p33_ASAP7_75t_R g4236 ( 
.A(n_4000),
.Y(n_4236)
);

BUFx6f_ASAP7_75t_L g4237 ( 
.A(n_4000),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4066),
.B(n_4068),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4044),
.Y(n_4239)
);

AOI21xp33_ASAP7_75t_L g4240 ( 
.A1(n_3935),
.A2(n_141),
.B(n_142),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3972),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_3887),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4076),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4076),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4100),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4104),
.Y(n_4246)
);

INVx1_ASAP7_75t_SL g4247 ( 
.A(n_4135),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4105),
.Y(n_4248)
);

CKINVDCx14_ASAP7_75t_R g4249 ( 
.A(n_4231),
.Y(n_4249)
);

AND2x4_ASAP7_75t_L g4250 ( 
.A(n_4095),
.B(n_3977),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4090),
.B(n_3984),
.Y(n_4251)
);

BUFx2_ASAP7_75t_SL g4252 ( 
.A(n_4191),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4117),
.Y(n_4253)
);

BUFx6f_ASAP7_75t_L g4254 ( 
.A(n_4216),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4120),
.Y(n_4255)
);

INVx2_ASAP7_75t_SL g4256 ( 
.A(n_4125),
.Y(n_4256)
);

BUFx3_ASAP7_75t_L g4257 ( 
.A(n_4089),
.Y(n_4257)
);

BUFx3_ASAP7_75t_L g4258 ( 
.A(n_4089),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4146),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4095),
.B(n_3980),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4097),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4127),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4130),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4078),
.B(n_4067),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4137),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4116),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4128),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4134),
.Y(n_4268)
);

BUFx6f_ASAP7_75t_L g4269 ( 
.A(n_4125),
.Y(n_4269)
);

INVx1_ASAP7_75t_SL g4270 ( 
.A(n_4133),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4140),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4147),
.Y(n_4272)
);

AOI21x1_ASAP7_75t_L g4273 ( 
.A1(n_4084),
.A2(n_3936),
.B(n_3988),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4151),
.Y(n_4274)
);

AOI21xp5_ASAP7_75t_L g4275 ( 
.A1(n_4141),
.A2(n_4030),
.B(n_3960),
.Y(n_4275)
);

OAI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_4107),
.A2(n_3929),
.B(n_4069),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4212),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4153),
.Y(n_4278)
);

OA21x2_ASAP7_75t_L g4279 ( 
.A1(n_4233),
.A2(n_3969),
.B(n_4035),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4235),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4158),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4161),
.Y(n_4282)
);

INVx2_ASAP7_75t_SL g4283 ( 
.A(n_4125),
.Y(n_4283)
);

INVxp67_ASAP7_75t_L g4284 ( 
.A(n_4164),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4169),
.Y(n_4285)
);

BUFx3_ASAP7_75t_L g4286 ( 
.A(n_4157),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4085),
.Y(n_4287)
);

INVxp67_ASAP7_75t_L g4288 ( 
.A(n_4131),
.Y(n_4288)
);

INVx3_ASAP7_75t_L g4289 ( 
.A(n_4183),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_4109),
.B(n_4048),
.Y(n_4290)
);

HB1xp67_ASAP7_75t_L g4291 ( 
.A(n_4179),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4172),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4119),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4186),
.Y(n_4294)
);

INVx2_ASAP7_75t_SL g4295 ( 
.A(n_4180),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4143),
.Y(n_4296)
);

AO21x1_ASAP7_75t_L g4297 ( 
.A1(n_4232),
.A2(n_4021),
.B(n_3904),
.Y(n_4297)
);

BUFx3_ASAP7_75t_L g4298 ( 
.A(n_4152),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4168),
.Y(n_4299)
);

BUFx3_ASAP7_75t_L g4300 ( 
.A(n_4180),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4109),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4209),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4167),
.Y(n_4303)
);

OA21x2_ASAP7_75t_L g4304 ( 
.A1(n_4103),
.A2(n_4242),
.B(n_4232),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4218),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4198),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4167),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4222),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4171),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4224),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4181),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4228),
.Y(n_4312)
);

AOI22xp33_ASAP7_75t_L g4313 ( 
.A1(n_4199),
.A2(n_4166),
.B1(n_4145),
.B2(n_4221),
.Y(n_4313)
);

BUFx3_ASAP7_75t_L g4314 ( 
.A(n_4176),
.Y(n_4314)
);

INVx3_ASAP7_75t_L g4315 ( 
.A(n_4183),
.Y(n_4315)
);

INVx3_ASAP7_75t_L g4316 ( 
.A(n_4184),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4079),
.B(n_4070),
.Y(n_4317)
);

BUFx6f_ASAP7_75t_L g4318 ( 
.A(n_4154),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4077),
.B(n_4024),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4206),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4239),
.Y(n_4321)
);

INVx3_ASAP7_75t_L g4322 ( 
.A(n_4184),
.Y(n_4322)
);

INVx2_ASAP7_75t_SL g4323 ( 
.A(n_4174),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4239),
.Y(n_4324)
);

INVx5_ASAP7_75t_L g4325 ( 
.A(n_4087),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4238),
.Y(n_4326)
);

OA21x2_ASAP7_75t_L g4327 ( 
.A1(n_4102),
.A2(n_3884),
.B(n_4055),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4188),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4144),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4188),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4155),
.Y(n_4331)
);

CKINVDCx6p67_ASAP7_75t_R g4332 ( 
.A(n_4096),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4121),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4121),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4087),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4193),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_4145),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4193),
.Y(n_4338)
);

INVxp33_ASAP7_75t_L g4339 ( 
.A(n_4094),
.Y(n_4339)
);

AND2x2_ASAP7_75t_L g4340 ( 
.A(n_4092),
.B(n_4050),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4214),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_4093),
.Y(n_4342)
);

AND2x2_ASAP7_75t_L g4343 ( 
.A(n_4093),
.B(n_4057),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4241),
.Y(n_4344)
);

BUFx2_ASAP7_75t_L g4345 ( 
.A(n_4220),
.Y(n_4345)
);

HB1xp67_ASAP7_75t_L g4346 ( 
.A(n_4241),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4210),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4187),
.Y(n_4348)
);

BUFx6f_ASAP7_75t_L g4349 ( 
.A(n_4154),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4226),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_4139),
.Y(n_4351)
);

INVx4_ASAP7_75t_L g4352 ( 
.A(n_4208),
.Y(n_4352)
);

AO21x2_ASAP7_75t_L g4353 ( 
.A1(n_4138),
.A2(n_3882),
.B(n_3881),
.Y(n_4353)
);

AND2x4_ASAP7_75t_L g4354 ( 
.A(n_4192),
.B(n_4048),
.Y(n_4354)
);

OAI21xp5_ASAP7_75t_SL g4355 ( 
.A1(n_4108),
.A2(n_4015),
.B(n_3979),
.Y(n_4355)
);

OR2x2_ASAP7_75t_L g4356 ( 
.A(n_4204),
.B(n_3903),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4200),
.Y(n_4357)
);

CKINVDCx5p33_ASAP7_75t_R g4358 ( 
.A(n_4236),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4200),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4211),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4201),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4118),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4202),
.Y(n_4363)
);

OR2x2_ASAP7_75t_L g4364 ( 
.A(n_4234),
.B(n_3956),
.Y(n_4364)
);

AND2x4_ASAP7_75t_L g4365 ( 
.A(n_4192),
.B(n_4048),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4200),
.Y(n_4366)
);

INVxp67_ASAP7_75t_L g4367 ( 
.A(n_4082),
.Y(n_4367)
);

BUFx2_ASAP7_75t_R g4368 ( 
.A(n_4156),
.Y(n_4368)
);

OAI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_4124),
.A2(n_3915),
.B(n_4038),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4237),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4237),
.Y(n_4371)
);

INVxp67_ASAP7_75t_SL g4372 ( 
.A(n_4083),
.Y(n_4372)
);

AND2x4_ASAP7_75t_L g4373 ( 
.A(n_4335),
.B(n_4192),
.Y(n_4373)
);

INVx4_ASAP7_75t_L g4374 ( 
.A(n_4254),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4350),
.B(n_4194),
.Y(n_4375)
);

BUFx3_ASAP7_75t_L g4376 ( 
.A(n_4254),
.Y(n_4376)
);

AOI222xp33_ASAP7_75t_L g4377 ( 
.A1(n_4313),
.A2(n_4217),
.B1(n_4159),
.B2(n_4113),
.C1(n_4129),
.C2(n_4219),
.Y(n_4377)
);

AND2x4_ASAP7_75t_L g4378 ( 
.A(n_4335),
.B(n_4237),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4288),
.B(n_4122),
.Y(n_4379)
);

AO21x2_ASAP7_75t_L g4380 ( 
.A1(n_4328),
.A2(n_4101),
.B(n_4185),
.Y(n_4380)
);

OAI221xp5_ASAP7_75t_L g4381 ( 
.A1(n_4313),
.A2(n_4080),
.B1(n_4081),
.B2(n_4110),
.C(n_4197),
.Y(n_4381)
);

INVx3_ASAP7_75t_SL g4382 ( 
.A(n_4351),
.Y(n_4382)
);

AOI22xp33_ASAP7_75t_L g4383 ( 
.A1(n_4339),
.A2(n_4199),
.B1(n_4173),
.B2(n_4240),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4339),
.A2(n_4223),
.B1(n_4086),
.B2(n_4160),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4301),
.Y(n_4385)
);

AOI22xp33_ASAP7_75t_L g4386 ( 
.A1(n_4337),
.A2(n_4297),
.B1(n_4311),
.B2(n_4309),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4337),
.A2(n_4088),
.B1(n_4163),
.B2(n_4098),
.Y(n_4387)
);

OAI22xp5_ASAP7_75t_L g4388 ( 
.A1(n_4368),
.A2(n_4126),
.B1(n_4132),
.B2(n_4091),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_L g4389 ( 
.A1(n_4309),
.A2(n_4112),
.B1(n_4148),
.B2(n_4175),
.Y(n_4389)
);

AOI22xp33_ASAP7_75t_L g4390 ( 
.A1(n_4311),
.A2(n_4229),
.B1(n_4207),
.B2(n_4106),
.Y(n_4390)
);

AOI22xp33_ASAP7_75t_L g4391 ( 
.A1(n_4276),
.A2(n_4195),
.B1(n_4099),
.B2(n_4123),
.Y(n_4391)
);

AOI221xp5_ASAP7_75t_L g4392 ( 
.A1(n_4360),
.A2(n_4165),
.B1(n_4225),
.B2(n_4230),
.C(n_4227),
.Y(n_4392)
);

HB1xp67_ASAP7_75t_L g4393 ( 
.A(n_4306),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4331),
.B(n_4178),
.Y(n_4394)
);

INVxp67_ASAP7_75t_L g4395 ( 
.A(n_4305),
.Y(n_4395)
);

BUFx8_ASAP7_75t_SL g4396 ( 
.A(n_4254),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_4348),
.A2(n_4367),
.B1(n_4363),
.B2(n_4329),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4300),
.B(n_4203),
.Y(n_4398)
);

AO21x2_ASAP7_75t_L g4399 ( 
.A1(n_4328),
.A2(n_4115),
.B(n_4114),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4243),
.Y(n_4400)
);

OAI211xp5_ASAP7_75t_L g4401 ( 
.A1(n_4355),
.A2(n_4136),
.B(n_4215),
.C(n_4162),
.Y(n_4401)
);

AOI22xp33_ASAP7_75t_L g4402 ( 
.A1(n_4367),
.A2(n_4205),
.B1(n_4111),
.B2(n_4189),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4364),
.A2(n_4142),
.B1(n_4178),
.B2(n_4170),
.Y(n_4403)
);

OAI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4372),
.A2(n_4213),
.B(n_4190),
.Y(n_4404)
);

OAI321xp33_ASAP7_75t_L g4405 ( 
.A1(n_4330),
.A2(n_4150),
.A3(n_4177),
.B1(n_4182),
.B2(n_3975),
.C(n_4008),
.Y(n_4405)
);

AOI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4369),
.A2(n_4009),
.B1(n_4149),
.B2(n_4040),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_4330),
.A2(n_4036),
.B1(n_3937),
.B2(n_3934),
.C(n_4041),
.Y(n_4407)
);

AOI21xp5_ASAP7_75t_L g4408 ( 
.A1(n_4275),
.A2(n_4001),
.B(n_4016),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4260),
.B(n_4196),
.Y(n_4409)
);

AOI221xp5_ASAP7_75t_L g4410 ( 
.A1(n_4282),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.C(n_146),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4319),
.A2(n_3973),
.B1(n_4023),
.B2(n_1412),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_4326),
.B(n_143),
.Y(n_4412)
);

AOI21xp5_ASAP7_75t_L g4413 ( 
.A1(n_4372),
.A2(n_146),
.B(n_147),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4244),
.Y(n_4414)
);

OAI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4342),
.A2(n_150),
.B1(n_147),
.B2(n_148),
.Y(n_4415)
);

OAI211xp5_ASAP7_75t_L g4416 ( 
.A1(n_4356),
.A2(n_152),
.B(n_148),
.C(n_151),
.Y(n_4416)
);

INVx3_ASAP7_75t_L g4417 ( 
.A(n_4314),
.Y(n_4417)
);

OAI22xp5_ASAP7_75t_L g4418 ( 
.A1(n_4249),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_4418)
);

HB1xp67_ASAP7_75t_L g4419 ( 
.A(n_4306),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4340),
.A2(n_1412),
.B1(n_1446),
.B2(n_1368),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4248),
.Y(n_4421)
);

OAI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4342),
.A2(n_162),
.B1(n_155),
.B2(n_160),
.Y(n_4422)
);

INVx3_ASAP7_75t_L g4423 ( 
.A(n_4314),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4302),
.B(n_162),
.Y(n_4424)
);

AOI22xp33_ASAP7_75t_L g4425 ( 
.A1(n_4333),
.A2(n_1446),
.B1(n_1694),
.B2(n_1685),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4334),
.A2(n_4250),
.B1(n_4361),
.B2(n_4362),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4326),
.B(n_165),
.Y(n_4427)
);

OAI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4270),
.A2(n_169),
.B1(n_166),
.B2(n_167),
.Y(n_4428)
);

HB1xp67_ASAP7_75t_L g4429 ( 
.A(n_4284),
.Y(n_4429)
);

INVx3_ASAP7_75t_L g4430 ( 
.A(n_4269),
.Y(n_4430)
);

OAI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4269),
.A2(n_171),
.B1(n_166),
.B2(n_169),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4301),
.Y(n_4432)
);

A2O1A1Ixp33_ASAP7_75t_L g4433 ( 
.A1(n_4249),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4248),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4291),
.Y(n_4435)
);

AOI221xp5_ASAP7_75t_L g4436 ( 
.A1(n_4308),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.C(n_177),
.Y(n_4436)
);

O2A1O1Ixp5_ASAP7_75t_L g4437 ( 
.A1(n_4287),
.A2(n_179),
.B(n_175),
.C(n_178),
.Y(n_4437)
);

OR2x2_ASAP7_75t_L g4438 ( 
.A(n_4259),
.B(n_180),
.Y(n_4438)
);

OR2x6_ASAP7_75t_L g4439 ( 
.A(n_4254),
.B(n_181),
.Y(n_4439)
);

AOI22xp33_ASAP7_75t_L g4440 ( 
.A1(n_4250),
.A2(n_1446),
.B1(n_1807),
.B2(n_1706),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4250),
.B(n_182),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4295),
.B(n_183),
.Y(n_4442)
);

AOI222xp33_ASAP7_75t_L g4443 ( 
.A1(n_4341),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C1(n_187),
.C2(n_188),
.Y(n_4443)
);

AOI222xp33_ASAP7_75t_L g4444 ( 
.A1(n_4341),
.A2(n_184),
.B1(n_188),
.B2(n_190),
.C1(n_191),
.C2(n_193),
.Y(n_4444)
);

AOI22xp33_ASAP7_75t_L g4445 ( 
.A1(n_4352),
.A2(n_1807),
.B1(n_1813),
.B2(n_1706),
.Y(n_4445)
);

BUFx3_ASAP7_75t_L g4446 ( 
.A(n_4358),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_4332),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_4352),
.A2(n_1807),
.B1(n_1813),
.B2(n_1706),
.Y(n_4448)
);

AOI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4298),
.A2(n_1816),
.B1(n_1859),
.B2(n_1813),
.Y(n_4449)
);

AOI221xp5_ASAP7_75t_L g4450 ( 
.A1(n_4310),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.C(n_195),
.Y(n_4450)
);

INVx4_ASAP7_75t_L g4451 ( 
.A(n_4298),
.Y(n_4451)
);

OA21x2_ASAP7_75t_L g4452 ( 
.A1(n_4287),
.A2(n_195),
.B(n_197),
.Y(n_4452)
);

O2A1O1Ixp33_ASAP7_75t_L g4453 ( 
.A1(n_4251),
.A2(n_201),
.B(n_198),
.C(n_199),
.Y(n_4453)
);

AOI22xp5_ASAP7_75t_L g4454 ( 
.A1(n_4353),
.A2(n_201),
.B1(n_198),
.B2(n_199),
.Y(n_4454)
);

OAI21x1_ASAP7_75t_L g4455 ( 
.A1(n_4321),
.A2(n_1859),
.B(n_1816),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4312),
.B(n_202),
.Y(n_4456)
);

AOI211xp5_ASAP7_75t_L g4457 ( 
.A1(n_4247),
.A2(n_205),
.B(n_202),
.C(n_203),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4291),
.Y(n_4458)
);

OAI22xp33_ASAP7_75t_SL g4459 ( 
.A1(n_4325),
.A2(n_4323),
.B1(n_4345),
.B2(n_4284),
.Y(n_4459)
);

O2A1O1Ixp33_ASAP7_75t_SL g4460 ( 
.A1(n_4256),
.A2(n_207),
.B(n_203),
.C(n_206),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4245),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_4257),
.A2(n_1859),
.B1(n_1870),
.B2(n_1816),
.Y(n_4462)
);

AOI22xp33_ASAP7_75t_L g4463 ( 
.A1(n_4258),
.A2(n_1892),
.B1(n_1912),
.B2(n_1870),
.Y(n_4463)
);

AOI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4258),
.A2(n_1892),
.B1(n_1912),
.B2(n_1870),
.Y(n_4464)
);

OAI22xp5_ASAP7_75t_L g4465 ( 
.A1(n_4269),
.A2(n_210),
.B1(n_207),
.B2(n_209),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_4303),
.Y(n_4466)
);

INVx3_ASAP7_75t_L g4467 ( 
.A(n_4269),
.Y(n_4467)
);

CKINVDCx5p33_ASAP7_75t_R g4468 ( 
.A(n_4351),
.Y(n_4468)
);

AO31x2_ASAP7_75t_L g4469 ( 
.A1(n_4294),
.A2(n_213),
.A3(n_209),
.B(n_210),
.Y(n_4469)
);

AOI221xp5_ASAP7_75t_L g4470 ( 
.A1(n_4320),
.A2(n_4253),
.B1(n_4255),
.B2(n_4246),
.C(n_4272),
.Y(n_4470)
);

AOI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4353),
.A2(n_216),
.B1(n_213),
.B2(n_214),
.Y(n_4471)
);

OAI211xp5_ASAP7_75t_L g4472 ( 
.A1(n_4304),
.A2(n_222),
.B(n_216),
.C(n_217),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4338),
.B(n_217),
.Y(n_4473)
);

AOI22xp33_ASAP7_75t_L g4474 ( 
.A1(n_4264),
.A2(n_4327),
.B1(n_4252),
.B2(n_4317),
.Y(n_4474)
);

OAI221xp5_ASAP7_75t_L g4475 ( 
.A1(n_4283),
.A2(n_4286),
.B1(n_4281),
.B2(n_4296),
.C(n_4293),
.Y(n_4475)
);

OAI22xp5_ASAP7_75t_L g4476 ( 
.A1(n_4273),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_4476)
);

OAI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4358),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_SL g4478 ( 
.A(n_4325),
.B(n_1541),
.Y(n_4478)
);

OAI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4336),
.A2(n_231),
.B1(n_226),
.B2(n_230),
.Y(n_4479)
);

AOI211xp5_ASAP7_75t_L g4480 ( 
.A1(n_4343),
.A2(n_235),
.B(n_232),
.C(n_234),
.Y(n_4480)
);

OAI211xp5_ASAP7_75t_L g4481 ( 
.A1(n_4304),
.A2(n_238),
.B(n_235),
.C(n_237),
.Y(n_4481)
);

INVxp67_ASAP7_75t_L g4482 ( 
.A(n_4262),
.Y(n_4482)
);

BUFx6f_ASAP7_75t_L g4483 ( 
.A(n_4286),
.Y(n_4483)
);

HB1xp67_ASAP7_75t_L g4484 ( 
.A(n_4304),
.Y(n_4484)
);

OAI22xp5_ASAP7_75t_L g4485 ( 
.A1(n_4370),
.A2(n_243),
.B1(n_239),
.B2(n_242),
.Y(n_4485)
);

OAI22xp33_ASAP7_75t_SL g4486 ( 
.A1(n_4325),
.A2(n_246),
.B1(n_242),
.B2(n_245),
.Y(n_4486)
);

AOI221xp5_ASAP7_75t_L g4487 ( 
.A1(n_4274),
.A2(n_247),
.B1(n_249),
.B2(n_251),
.C(n_252),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4303),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4263),
.Y(n_4489)
);

OR2x2_ASAP7_75t_L g4490 ( 
.A(n_4267),
.B(n_253),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4400),
.Y(n_4491)
);

OAI33xp33_ASAP7_75t_L g4492 ( 
.A1(n_4428),
.A2(n_4344),
.A3(n_4265),
.B1(n_4278),
.B2(n_4294),
.B3(n_4271),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4484),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4414),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4385),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4432),
.Y(n_4496)
);

OR2x2_ASAP7_75t_L g4497 ( 
.A(n_4379),
.B(n_4299),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4466),
.Y(n_4498)
);

AND2x4_ASAP7_75t_L g4499 ( 
.A(n_4417),
.B(n_4423),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4488),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4375),
.B(n_4397),
.Y(n_4501)
);

NAND2x1_ASAP7_75t_L g4502 ( 
.A(n_4373),
.B(n_4289),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4489),
.Y(n_4503)
);

BUFx3_ASAP7_75t_L g4504 ( 
.A(n_4396),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4417),
.B(n_4315),
.Y(n_4505)
);

AND2x4_ASAP7_75t_L g4506 ( 
.A(n_4423),
.B(n_4435),
.Y(n_4506)
);

INVx3_ASAP7_75t_L g4507 ( 
.A(n_4451),
.Y(n_4507)
);

INVx6_ASAP7_75t_L g4508 ( 
.A(n_4374),
.Y(n_4508)
);

AOI22xp33_ASAP7_75t_L g4509 ( 
.A1(n_4377),
.A2(n_4327),
.B1(n_4279),
.B2(n_4324),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4421),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4386),
.B(n_4285),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4395),
.B(n_4473),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4409),
.B(n_4315),
.Y(n_4513)
);

INVx4_ASAP7_75t_L g4514 ( 
.A(n_4374),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4461),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4429),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_4398),
.B(n_4316),
.Y(n_4517)
);

AND2x4_ASAP7_75t_SL g4518 ( 
.A(n_4451),
.B(n_4316),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4434),
.Y(n_4519)
);

NAND2x1_ASAP7_75t_L g4520 ( 
.A(n_4373),
.B(n_4322),
.Y(n_4520)
);

BUFx2_ASAP7_75t_L g4521 ( 
.A(n_4376),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4426),
.B(n_4322),
.Y(n_4522)
);

AND2x4_ASAP7_75t_SL g4523 ( 
.A(n_4441),
.B(n_4318),
.Y(n_4523)
);

INVxp67_ASAP7_75t_SL g4524 ( 
.A(n_4393),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4482),
.Y(n_4525)
);

INVx3_ASAP7_75t_L g4526 ( 
.A(n_4483),
.Y(n_4526)
);

OAI211xp5_ASAP7_75t_L g4527 ( 
.A1(n_4457),
.A2(n_4383),
.B(n_4480),
.C(n_4433),
.Y(n_4527)
);

AND2x4_ASAP7_75t_L g4528 ( 
.A(n_4458),
.B(n_4441),
.Y(n_4528)
);

OR2x2_ASAP7_75t_L g4529 ( 
.A(n_4394),
.B(n_4261),
.Y(n_4529)
);

BUFx3_ASAP7_75t_L g4530 ( 
.A(n_4483),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4419),
.Y(n_4531)
);

NOR2xp33_ASAP7_75t_L g4532 ( 
.A(n_4483),
.B(n_4371),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4469),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4469),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4469),
.Y(n_4535)
);

INVx5_ASAP7_75t_L g4536 ( 
.A(n_4439),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4452),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4452),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4430),
.Y(n_4539)
);

NOR2x1_ASAP7_75t_SL g4540 ( 
.A(n_4439),
.B(n_4325),
.Y(n_4540)
);

INVx5_ASAP7_75t_L g4541 ( 
.A(n_4439),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4490),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4430),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4412),
.Y(n_4544)
);

OR2x2_ASAP7_75t_L g4545 ( 
.A(n_4438),
.B(n_4266),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_4446),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_4381),
.B(n_4357),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4467),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4470),
.B(n_4266),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4427),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4467),
.B(n_4378),
.Y(n_4551)
);

CKINVDCx11_ASAP7_75t_R g4552 ( 
.A(n_4382),
.Y(n_4552)
);

BUFx2_ASAP7_75t_L g4553 ( 
.A(n_4447),
.Y(n_4553)
);

INVx3_ASAP7_75t_L g4554 ( 
.A(n_4378),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4442),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4399),
.Y(n_4556)
);

BUFx6f_ASAP7_75t_L g4557 ( 
.A(n_4478),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4474),
.B(n_4359),
.Y(n_4558)
);

INVxp67_ASAP7_75t_L g4559 ( 
.A(n_4424),
.Y(n_4559)
);

BUFx6f_ASAP7_75t_L g4560 ( 
.A(n_4456),
.Y(n_4560)
);

HB1xp67_ASAP7_75t_L g4561 ( 
.A(n_4399),
.Y(n_4561)
);

AND2x4_ASAP7_75t_L g4562 ( 
.A(n_4380),
.B(n_4277),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4380),
.B(n_4366),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4440),
.B(n_4307),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4475),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4455),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4437),
.Y(n_4567)
);

INVx2_ASAP7_75t_SL g4568 ( 
.A(n_4468),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4404),
.B(n_4307),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4454),
.Y(n_4570)
);

NOR4xp25_ASAP7_75t_SL g4571 ( 
.A(n_4459),
.B(n_4349),
.C(n_4318),
.D(n_4346),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4454),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4471),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4471),
.B(n_4268),
.Y(n_4574)
);

HB1xp67_ASAP7_75t_L g4575 ( 
.A(n_4472),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4476),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4481),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4479),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4486),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4418),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4392),
.B(n_4268),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4491),
.Y(n_4582)
);

OAI221xp5_ASAP7_75t_L g4583 ( 
.A1(n_4527),
.A2(n_4384),
.B1(n_4391),
.B2(n_4387),
.C(n_4413),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4551),
.B(n_4318),
.Y(n_4584)
);

NAND3xp33_ASAP7_75t_SL g4585 ( 
.A(n_4575),
.B(n_4453),
.C(n_4416),
.Y(n_4585)
);

CKINVDCx6p67_ASAP7_75t_R g4586 ( 
.A(n_4536),
.Y(n_4586)
);

OAI22xp5_ASAP7_75t_L g4587 ( 
.A1(n_4572),
.A2(n_4390),
.B1(n_4388),
.B2(n_4389),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4508),
.Y(n_4588)
);

HB1xp67_ASAP7_75t_L g4589 ( 
.A(n_4493),
.Y(n_4589)
);

NAND3xp33_ASAP7_75t_L g4590 ( 
.A(n_4572),
.B(n_4575),
.C(n_4509),
.Y(n_4590)
);

NAND3xp33_ASAP7_75t_L g4591 ( 
.A(n_4509),
.B(n_4444),
.C(n_4443),
.Y(n_4591)
);

AOI22xp33_ASAP7_75t_L g4592 ( 
.A1(n_4570),
.A2(n_4487),
.B1(n_4410),
.B2(n_4450),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_4508),
.Y(n_4593)
);

INVx3_ASAP7_75t_L g4594 ( 
.A(n_4514),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4494),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4503),
.Y(n_4596)
);

AOI22xp33_ASAP7_75t_L g4597 ( 
.A1(n_4570),
.A2(n_4573),
.B1(n_4501),
.B2(n_4576),
.Y(n_4597)
);

AOI22xp33_ASAP7_75t_L g4598 ( 
.A1(n_4576),
.A2(n_4436),
.B1(n_4465),
.B2(n_4431),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4508),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4521),
.B(n_4318),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4499),
.B(n_4349),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4499),
.B(n_4349),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4530),
.Y(n_4603)
);

AND2x2_ASAP7_75t_SL g4604 ( 
.A(n_4567),
.B(n_4402),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4530),
.Y(n_4605)
);

AOI211xp5_ASAP7_75t_L g4606 ( 
.A1(n_4577),
.A2(n_4415),
.B(n_4422),
.C(n_4477),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4515),
.Y(n_4607)
);

NAND3xp33_ASAP7_75t_L g4608 ( 
.A(n_4567),
.B(n_4460),
.C(n_4485),
.Y(n_4608)
);

OAI22xp5_ASAP7_75t_L g4609 ( 
.A1(n_4536),
.A2(n_4403),
.B1(n_4408),
.B2(n_4406),
.Y(n_4609)
);

AOI22xp33_ASAP7_75t_L g4610 ( 
.A1(n_4579),
.A2(n_4565),
.B1(n_4492),
.B2(n_4547),
.Y(n_4610)
);

OAI222xp33_ASAP7_75t_L g4611 ( 
.A1(n_4536),
.A2(n_4406),
.B1(n_4411),
.B2(n_4277),
.C1(n_4280),
.C2(n_4321),
.Y(n_4611)
);

NAND3xp33_ASAP7_75t_L g4612 ( 
.A(n_4536),
.B(n_4541),
.C(n_4571),
.Y(n_4612)
);

NAND3xp33_ASAP7_75t_L g4613 ( 
.A(n_4541),
.B(n_4401),
.C(n_4420),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_L g4614 ( 
.A(n_4504),
.B(n_4405),
.Y(n_4614)
);

OAI22xp5_ASAP7_75t_L g4615 ( 
.A1(n_4541),
.A2(n_4425),
.B1(n_4354),
.B2(n_4365),
.Y(n_4615)
);

OAI211xp5_ASAP7_75t_L g4616 ( 
.A1(n_4541),
.A2(n_4407),
.B(n_4448),
.C(n_4445),
.Y(n_4616)
);

NAND4xp75_ASAP7_75t_L g4617 ( 
.A(n_4563),
.B(n_4327),
.C(n_4279),
.D(n_4324),
.Y(n_4617)
);

OAI33xp33_ASAP7_75t_L g4618 ( 
.A1(n_4537),
.A2(n_4280),
.A3(n_4292),
.B1(n_256),
.B2(n_257),
.B3(n_258),
.Y(n_4618)
);

OAI221xp5_ASAP7_75t_L g4619 ( 
.A1(n_4547),
.A2(n_4449),
.B1(n_4463),
.B2(n_4462),
.C(n_4464),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4493),
.Y(n_4620)
);

INVxp67_ASAP7_75t_L g4621 ( 
.A(n_4540),
.Y(n_4621)
);

OAI31xp33_ASAP7_75t_L g4622 ( 
.A1(n_4581),
.A2(n_4365),
.A3(n_4354),
.B(n_4290),
.Y(n_4622)
);

OAI33xp33_ASAP7_75t_L g4623 ( 
.A1(n_4538),
.A2(n_254),
.A3(n_255),
.B1(n_256),
.B2(n_257),
.B3(n_258),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4499),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4542),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4578),
.B(n_4560),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4580),
.A2(n_4347),
.B1(n_4365),
.B2(n_4354),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4580),
.A2(n_4347),
.B1(n_4279),
.B2(n_4290),
.Y(n_4628)
);

AOI221xp5_ASAP7_75t_L g4629 ( 
.A1(n_4578),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_4629)
);

NOR2xp33_ASAP7_75t_L g4630 ( 
.A(n_4504),
.B(n_259),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4524),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4526),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4526),
.Y(n_4633)
);

OAI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4511),
.A2(n_262),
.B(n_265),
.Y(n_4634)
);

CKINVDCx14_ASAP7_75t_R g4635 ( 
.A(n_4552),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4524),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4546),
.Y(n_4637)
);

AOI22xp33_ASAP7_75t_SL g4638 ( 
.A1(n_4560),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4574),
.A2(n_267),
.B(n_268),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4545),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4505),
.B(n_268),
.Y(n_4641)
);

AOI21xp5_ASAP7_75t_L g4642 ( 
.A1(n_4549),
.A2(n_269),
.B(n_270),
.Y(n_4642)
);

NAND4xp25_ASAP7_75t_L g4643 ( 
.A(n_4559),
.B(n_271),
.C(n_273),
.D(n_274),
.Y(n_4643)
);

AOI31xp33_ASAP7_75t_L g4644 ( 
.A1(n_4568),
.A2(n_273),
.A3(n_274),
.B(n_277),
.Y(n_4644)
);

OA21x2_ASAP7_75t_L g4645 ( 
.A1(n_4556),
.A2(n_277),
.B(n_278),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4589),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4601),
.B(n_4554),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4624),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4602),
.B(n_4554),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4586),
.B(n_4514),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4589),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4620),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4594),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4631),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4642),
.B(n_4560),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4636),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4594),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4637),
.B(n_4514),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4588),
.B(n_4507),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4626),
.B(n_4531),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4593),
.B(n_4507),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4599),
.B(n_4506),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4645),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4590),
.B(n_4531),
.Y(n_4664)
);

NOR2xp67_ASAP7_75t_L g4665 ( 
.A(n_4612),
.B(n_4568),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4645),
.Y(n_4666)
);

INVxp67_ASAP7_75t_L g4667 ( 
.A(n_4614),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4621),
.B(n_4506),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4582),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4603),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4642),
.B(n_4560),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4584),
.B(n_4506),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4605),
.B(n_4518),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4639),
.B(n_4559),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4632),
.B(n_4518),
.Y(n_4675)
);

BUFx2_ASAP7_75t_L g4676 ( 
.A(n_4635),
.Y(n_4676)
);

INVxp67_ASAP7_75t_SL g4677 ( 
.A(n_4621),
.Y(n_4677)
);

AOI22xp33_ASAP7_75t_L g4678 ( 
.A1(n_4591),
.A2(n_4569),
.B1(n_4558),
.B2(n_4522),
.Y(n_4678)
);

NAND2x1p5_ASAP7_75t_L g4679 ( 
.A(n_4639),
.B(n_4502),
.Y(n_4679)
);

OR2x2_ASAP7_75t_L g4680 ( 
.A(n_4625),
.B(n_4516),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4633),
.B(n_4539),
.Y(n_4681)
);

NOR2xp33_ASAP7_75t_L g4682 ( 
.A(n_4583),
.B(n_4552),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4595),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4600),
.Y(n_4684)
);

OR2x2_ASAP7_75t_L g4685 ( 
.A(n_4640),
.B(n_4533),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4677),
.B(n_4610),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4676),
.B(n_4604),
.Y(n_4687)
);

AOI22xp33_ASAP7_75t_L g4688 ( 
.A1(n_4667),
.A2(n_4585),
.B1(n_4604),
.B2(n_4587),
.Y(n_4688)
);

INVx4_ASAP7_75t_L g4689 ( 
.A(n_4676),
.Y(n_4689)
);

NOR2x1p5_ASAP7_75t_L g4690 ( 
.A(n_4655),
.B(n_4585),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4678),
.B(n_4597),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4668),
.Y(n_4692)
);

BUFx3_ASAP7_75t_L g4693 ( 
.A(n_4650),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4646),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4672),
.B(n_4627),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4684),
.B(n_4608),
.Y(n_4696)
);

AOI33xp33_ASAP7_75t_L g4697 ( 
.A1(n_4670),
.A2(n_4592),
.A3(n_4598),
.B1(n_4638),
.B2(n_4606),
.B3(n_4629),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4668),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4646),
.Y(n_4699)
);

AOI22xp33_ASAP7_75t_L g4700 ( 
.A1(n_4682),
.A2(n_4609),
.B1(n_4613),
.B2(n_4592),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4672),
.B(n_4520),
.Y(n_4701)
);

OAI31xp33_ASAP7_75t_L g4702 ( 
.A1(n_4679),
.A2(n_4611),
.A3(n_4616),
.B(n_4643),
.Y(n_4702)
);

AOI22xp5_ASAP7_75t_L g4703 ( 
.A1(n_4665),
.A2(n_4618),
.B1(n_4623),
.B2(n_4616),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4651),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4651),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4668),
.Y(n_4706)
);

BUFx3_ASAP7_75t_L g4707 ( 
.A(n_4650),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4684),
.B(n_4644),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4666),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_SL g4710 ( 
.A(n_4679),
.B(n_4546),
.Y(n_4710)
);

OAI31xp33_ASAP7_75t_L g4711 ( 
.A1(n_4679),
.A2(n_4611),
.A3(n_4615),
.B(n_4562),
.Y(n_4711)
);

OAI22xp5_ASAP7_75t_L g4712 ( 
.A1(n_4674),
.A2(n_4634),
.B1(n_4638),
.B2(n_4628),
.Y(n_4712)
);

HB1xp67_ASAP7_75t_L g4713 ( 
.A(n_4709),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4689),
.B(n_4673),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4689),
.B(n_4673),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_4689),
.B(n_4670),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4694),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4687),
.B(n_4658),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4687),
.B(n_4658),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4692),
.B(n_4659),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4694),
.Y(n_4721)
);

AND2x4_ASAP7_75t_L g4722 ( 
.A(n_4692),
.B(n_4652),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4698),
.B(n_4659),
.Y(n_4723)
);

INVx3_ASAP7_75t_L g4724 ( 
.A(n_4698),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4701),
.B(n_4662),
.Y(n_4725)
);

AND2x2_ASAP7_75t_SL g4726 ( 
.A(n_4688),
.B(n_4671),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4699),
.Y(n_4727)
);

INVx2_ASAP7_75t_SL g4728 ( 
.A(n_4706),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4706),
.Y(n_4729)
);

HB1xp67_ASAP7_75t_L g4730 ( 
.A(n_4709),
.Y(n_4730)
);

NAND5xp2_ASAP7_75t_L g4731 ( 
.A(n_4718),
.B(n_4700),
.C(n_4702),
.D(n_4686),
.E(n_4691),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4725),
.B(n_4661),
.Y(n_4732)
);

NAND4xp25_ASAP7_75t_L g4733 ( 
.A(n_4719),
.B(n_4696),
.C(n_4697),
.D(n_4693),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4724),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4714),
.B(n_4661),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4715),
.B(n_4693),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4713),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4713),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4720),
.B(n_4664),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4730),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4724),
.B(n_4707),
.Y(n_4741)
);

NAND4xp25_ASAP7_75t_SL g4742 ( 
.A(n_4716),
.B(n_4703),
.C(n_4711),
.D(n_4708),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4728),
.B(n_4690),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4723),
.B(n_4707),
.Y(n_4744)
);

INVx3_ASAP7_75t_L g4745 ( 
.A(n_4722),
.Y(n_4745)
);

INVx1_ASAP7_75t_SL g4746 ( 
.A(n_4730),
.Y(n_4746)
);

AND2x4_ASAP7_75t_SL g4747 ( 
.A(n_4722),
.B(n_4546),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4728),
.Y(n_4748)
);

INVx1_ASAP7_75t_SL g4749 ( 
.A(n_4741),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4745),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4735),
.B(n_4701),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4732),
.B(n_4662),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4746),
.Y(n_4753)
);

NOR2x1_ASAP7_75t_L g4754 ( 
.A(n_4745),
.B(n_4710),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4736),
.B(n_4726),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4744),
.B(n_4695),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4748),
.B(n_4726),
.Y(n_4757)
);

OR2x2_ASAP7_75t_L g4758 ( 
.A(n_4739),
.B(n_4664),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4734),
.B(n_4722),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4756),
.B(n_4747),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4750),
.Y(n_4761)
);

OR2x2_ASAP7_75t_L g4762 ( 
.A(n_4758),
.B(n_4733),
.Y(n_4762)
);

OAI211xp5_ASAP7_75t_L g4763 ( 
.A1(n_4757),
.A2(n_4743),
.B(n_4746),
.C(n_4737),
.Y(n_4763)
);

INVxp67_ASAP7_75t_SL g4764 ( 
.A(n_4754),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4751),
.B(n_4729),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4759),
.Y(n_4766)
);

AOI221xp5_ASAP7_75t_L g4767 ( 
.A1(n_4753),
.A2(n_4731),
.B1(n_4742),
.B2(n_4712),
.C(n_4743),
.Y(n_4767)
);

INVxp67_ASAP7_75t_L g4768 ( 
.A(n_4755),
.Y(n_4768)
);

AOI221xp5_ASAP7_75t_L g4769 ( 
.A1(n_4767),
.A2(n_4731),
.B1(n_4742),
.B2(n_4738),
.C(n_4740),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4764),
.B(n_4752),
.Y(n_4770)
);

OAI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4768),
.A2(n_4749),
.B(n_4753),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4761),
.Y(n_4772)
);

OAI22xp5_ASAP7_75t_L g4773 ( 
.A1(n_4762),
.A2(n_4760),
.B1(n_4660),
.B2(n_4663),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4763),
.Y(n_4774)
);

OAI322xp33_ASAP7_75t_L g4775 ( 
.A1(n_4766),
.A2(n_4729),
.A3(n_4727),
.B1(n_4721),
.B2(n_4717),
.C1(n_4705),
.C2(n_4704),
.Y(n_4775)
);

NAND5xp2_ASAP7_75t_SL g4776 ( 
.A(n_4767),
.B(n_4695),
.C(n_4675),
.D(n_4647),
.E(n_4649),
.Y(n_4776)
);

AOI221xp5_ASAP7_75t_L g4777 ( 
.A1(n_4767),
.A2(n_4656),
.B1(n_4654),
.B2(n_4663),
.C(n_4657),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4765),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4769),
.A2(n_4657),
.B(n_4653),
.Y(n_4779)
);

NOR2xp67_ASAP7_75t_L g4780 ( 
.A(n_4778),
.B(n_4653),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4774),
.B(n_4656),
.Y(n_4781)
);

AOI211x1_ASAP7_75t_L g4782 ( 
.A1(n_4771),
.A2(n_4683),
.B(n_4669),
.C(n_4675),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4770),
.B(n_4553),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4773),
.Y(n_4784)
);

AND2x2_ASAP7_75t_L g4785 ( 
.A(n_4772),
.B(n_4647),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4785),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4780),
.B(n_4777),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4783),
.B(n_4648),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4782),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4781),
.Y(n_4790)
);

AOI21xp33_ASAP7_75t_SL g4791 ( 
.A1(n_4784),
.A2(n_4630),
.B(n_4776),
.Y(n_4791)
);

O2A1O1Ixp33_ASAP7_75t_L g4792 ( 
.A1(n_4779),
.A2(n_4775),
.B(n_4683),
.C(n_4561),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4787),
.Y(n_4793)
);

XOR2xp5_ASAP7_75t_L g4794 ( 
.A(n_4786),
.B(n_4546),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_SL g4795 ( 
.A(n_4791),
.B(n_4649),
.Y(n_4795)
);

AOI22xp33_ASAP7_75t_L g4796 ( 
.A1(n_4789),
.A2(n_4681),
.B1(n_4685),
.B2(n_4680),
.Y(n_4796)
);

OAI322xp33_ASAP7_75t_L g4797 ( 
.A1(n_4788),
.A2(n_4685),
.A3(n_4680),
.B1(n_4556),
.B2(n_4596),
.C1(n_4607),
.C2(n_4681),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4792),
.B(n_4641),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4790),
.Y(n_4799)
);

XNOR2xp5_ASAP7_75t_L g4800 ( 
.A(n_4786),
.B(n_4523),
.Y(n_4800)
);

A2O1A1Ixp33_ASAP7_75t_L g4801 ( 
.A1(n_4792),
.A2(n_4622),
.B(n_4562),
.C(n_4532),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4787),
.Y(n_4802)
);

INVx1_ASAP7_75t_SL g4803 ( 
.A(n_4787),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4786),
.B(n_4525),
.Y(n_4804)
);

XOR2x2_ASAP7_75t_L g4805 ( 
.A(n_4788),
.B(n_4617),
.Y(n_4805)
);

AO22x2_ASAP7_75t_L g4806 ( 
.A1(n_4794),
.A2(n_4543),
.B1(n_4548),
.B2(n_4539),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4796),
.B(n_4528),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4800),
.B(n_4528),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4804),
.B(n_4555),
.Y(n_4809)
);

AOI22xp5_ASAP7_75t_L g4810 ( 
.A1(n_4803),
.A2(n_4798),
.B1(n_4802),
.B2(n_4793),
.Y(n_4810)
);

INVx6_ASAP7_75t_L g4811 ( 
.A(n_4799),
.Y(n_4811)
);

NOR3xp33_ASAP7_75t_L g4812 ( 
.A(n_4801),
.B(n_4512),
.C(n_4534),
.Y(n_4812)
);

NOR2xp33_ASAP7_75t_L g4813 ( 
.A(n_4797),
.B(n_4543),
.Y(n_4813)
);

NAND3xp33_ASAP7_75t_L g4814 ( 
.A(n_4805),
.B(n_4557),
.C(n_4535),
.Y(n_4814)
);

AOI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4795),
.A2(n_4550),
.B(n_4544),
.Y(n_4815)
);

XNOR2x2_ASAP7_75t_L g4816 ( 
.A(n_4803),
.B(n_4548),
.Y(n_4816)
);

NOR2xp33_ASAP7_75t_L g4817 ( 
.A(n_4795),
.B(n_4497),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4804),
.B(n_4517),
.Y(n_4818)
);

XNOR2x2_ASAP7_75t_L g4819 ( 
.A(n_4803),
.B(n_4619),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4794),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4807),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4818),
.Y(n_4822)
);

INVx1_ASAP7_75t_SL g4823 ( 
.A(n_4816),
.Y(n_4823)
);

AOI322xp5_ASAP7_75t_L g4824 ( 
.A1(n_4817),
.A2(n_4495),
.A3(n_4496),
.B1(n_4498),
.B2(n_4500),
.C1(n_4519),
.C2(n_4510),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4812),
.B(n_4813),
.Y(n_4825)
);

CKINVDCx5p33_ASAP7_75t_R g4826 ( 
.A(n_4810),
.Y(n_4826)
);

AOI221xp5_ASAP7_75t_L g4827 ( 
.A1(n_4814),
.A2(n_4523),
.B1(n_4510),
.B2(n_4519),
.C(n_4566),
.Y(n_4827)
);

OAI221xp5_ASAP7_75t_SL g4828 ( 
.A1(n_4808),
.A2(n_4529),
.B1(n_4564),
.B2(n_4513),
.C(n_284),
.Y(n_4828)
);

INVx1_ASAP7_75t_SL g4829 ( 
.A(n_4811),
.Y(n_4829)
);

NOR3xp33_ASAP7_75t_L g4830 ( 
.A(n_4820),
.B(n_279),
.C(n_281),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4809),
.Y(n_4831)
);

AOI211xp5_ASAP7_75t_L g4832 ( 
.A1(n_4815),
.A2(n_282),
.B(n_285),
.C(n_287),
.Y(n_4832)
);

AOI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_4806),
.A2(n_1495),
.B1(n_1521),
.B2(n_1540),
.Y(n_4833)
);

NAND4xp25_ASAP7_75t_L g4834 ( 
.A(n_4806),
.B(n_297),
.C(n_298),
.D(n_299),
.Y(n_4834)
);

XNOR2xp5_ASAP7_75t_L g4835 ( 
.A(n_4819),
.B(n_300),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4807),
.Y(n_4836)
);

NOR3xp33_ASAP7_75t_L g4837 ( 
.A(n_4821),
.B(n_303),
.C(n_305),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_SL g4838 ( 
.A(n_4826),
.B(n_1495),
.Y(n_4838)
);

AOI211x1_ASAP7_75t_SL g4839 ( 
.A1(n_4825),
.A2(n_310),
.B(n_317),
.C(n_319),
.Y(n_4839)
);

NOR2x1_ASAP7_75t_L g4840 ( 
.A(n_4834),
.B(n_4823),
.Y(n_4840)
);

AND2x4_ASAP7_75t_L g4841 ( 
.A(n_4822),
.B(n_320),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_SL g4842 ( 
.A(n_4829),
.B(n_1495),
.Y(n_4842)
);

NOR3xp33_ASAP7_75t_L g4843 ( 
.A(n_4836),
.B(n_324),
.C(n_325),
.Y(n_4843)
);

BUFx3_ASAP7_75t_L g4844 ( 
.A(n_4831),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4830),
.B(n_328),
.Y(n_4845)
);

A2O1A1Ixp33_ASAP7_75t_L g4846 ( 
.A1(n_4832),
.A2(n_331),
.B(n_333),
.C(n_336),
.Y(n_4846)
);

NOR3xp33_ASAP7_75t_L g4847 ( 
.A(n_4828),
.B(n_340),
.C(n_341),
.Y(n_4847)
);

NOR3xp33_ASAP7_75t_L g4848 ( 
.A(n_4833),
.B(n_345),
.C(n_346),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_SL g4849 ( 
.A(n_4827),
.B(n_1495),
.Y(n_4849)
);

NOR2xp33_ASAP7_75t_SL g4850 ( 
.A(n_4824),
.B(n_1521),
.Y(n_4850)
);

NAND3xp33_ASAP7_75t_SL g4851 ( 
.A(n_4829),
.B(n_349),
.C(n_351),
.Y(n_4851)
);

NOR2x1_ASAP7_75t_L g4852 ( 
.A(n_4835),
.B(n_353),
.Y(n_4852)
);

NOR2x1_ASAP7_75t_L g4853 ( 
.A(n_4835),
.B(n_354),
.Y(n_4853)
);

AOI22xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4844),
.A2(n_1521),
.B1(n_1540),
.B2(n_1466),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4852),
.Y(n_4855)
);

AOI221xp5_ASAP7_75t_SL g4856 ( 
.A1(n_4849),
.A2(n_383),
.B1(n_385),
.B2(n_389),
.C(n_391),
.Y(n_4856)
);

NOR4xp75_ASAP7_75t_L g4857 ( 
.A(n_4845),
.B(n_392),
.C(n_393),
.D(n_396),
.Y(n_4857)
);

AOI221xp5_ASAP7_75t_L g4858 ( 
.A1(n_4847),
.A2(n_2067),
.B1(n_2066),
.B2(n_2049),
.C(n_2031),
.Y(n_4858)
);

XNOR2xp5_ASAP7_75t_L g4859 ( 
.A(n_4840),
.B(n_402),
.Y(n_4859)
);

O2A1O1Ixp33_ASAP7_75t_L g4860 ( 
.A1(n_4846),
.A2(n_403),
.B(n_409),
.C(n_410),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4841),
.Y(n_4861)
);

AOI221xp5_ASAP7_75t_SL g4862 ( 
.A1(n_4838),
.A2(n_411),
.B1(n_412),
.B2(n_416),
.C(n_421),
.Y(n_4862)
);

AOI221x1_ASAP7_75t_L g4863 ( 
.A1(n_4848),
.A2(n_422),
.B1(n_428),
.B2(n_432),
.C(n_437),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4859),
.Y(n_4864)
);

NAND5xp2_ASAP7_75t_L g4865 ( 
.A(n_4856),
.B(n_4850),
.C(n_4837),
.D(n_4843),
.E(n_4853),
.Y(n_4865)
);

AOI322xp5_ASAP7_75t_L g4866 ( 
.A1(n_4855),
.A2(n_4851),
.A3(n_4842),
.B1(n_4839),
.B2(n_4841),
.C1(n_444),
.C2(n_446),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4861),
.B(n_438),
.Y(n_4867)
);

NOR2x1_ASAP7_75t_L g4868 ( 
.A(n_4860),
.B(n_450),
.Y(n_4868)
);

NOR3xp33_ASAP7_75t_L g4869 ( 
.A(n_4858),
.B(n_4862),
.C(n_4854),
.Y(n_4869)
);

XOR2xp5_ASAP7_75t_L g4870 ( 
.A(n_4857),
.B(n_456),
.Y(n_4870)
);

XNOR2xp5_ASAP7_75t_L g4871 ( 
.A(n_4863),
.B(n_467),
.Y(n_4871)
);

AND3x2_ASAP7_75t_L g4872 ( 
.A(n_4855),
.B(n_468),
.C(n_470),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4872),
.Y(n_4873)
);

AO22x2_ASAP7_75t_L g4874 ( 
.A1(n_4864),
.A2(n_471),
.B1(n_476),
.B2(n_479),
.Y(n_4874)
);

AOI22xp5_ASAP7_75t_L g4875 ( 
.A1(n_4870),
.A2(n_1839),
.B1(n_2066),
.B2(n_2049),
.Y(n_4875)
);

AND4x1_ASAP7_75t_L g4876 ( 
.A(n_4868),
.B(n_498),
.C(n_505),
.D(n_507),
.Y(n_4876)
);

NOR4xp25_ASAP7_75t_L g4877 ( 
.A(n_4867),
.B(n_508),
.C(n_509),
.D(n_512),
.Y(n_4877)
);

NOR3xp33_ASAP7_75t_L g4878 ( 
.A(n_4865),
.B(n_514),
.C(n_517),
.Y(n_4878)
);

AOI211xp5_ASAP7_75t_L g4879 ( 
.A1(n_4871),
.A2(n_522),
.B(n_523),
.C(n_1879),
.Y(n_4879)
);

OAI211xp5_ASAP7_75t_L g4880 ( 
.A1(n_4866),
.A2(n_1892),
.B(n_1967),
.C(n_1952),
.Y(n_4880)
);

OR5x1_ASAP7_75t_L g4881 ( 
.A(n_4869),
.B(n_1967),
.C(n_1952),
.D(n_1912),
.E(n_2067),
.Y(n_4881)
);

NOR4xp25_ASAP7_75t_L g4882 ( 
.A(n_4864),
.B(n_1868),
.C(n_2031),
.D(n_2025),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4873),
.B(n_1541),
.Y(n_4883)
);

AND3x2_ASAP7_75t_L g4884 ( 
.A(n_4878),
.B(n_1868),
.C(n_2031),
.Y(n_4884)
);

OAI22xp5_ASAP7_75t_L g4885 ( 
.A1(n_4875),
.A2(n_1868),
.B1(n_2025),
.B2(n_2009),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4876),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4879),
.Y(n_4887)
);

HB1xp67_ASAP7_75t_L g4888 ( 
.A(n_4877),
.Y(n_4888)
);

NAND3x1_ASAP7_75t_L g4889 ( 
.A(n_4880),
.B(n_1855),
.C(n_2009),
.Y(n_4889)
);

HB1xp67_ASAP7_75t_L g4890 ( 
.A(n_4874),
.Y(n_4890)
);

OAI22xp5_ASAP7_75t_SL g4891 ( 
.A1(n_4881),
.A2(n_1855),
.B1(n_2009),
.B2(n_2008),
.Y(n_4891)
);

NOR3xp33_ASAP7_75t_L g4892 ( 
.A(n_4888),
.B(n_4882),
.C(n_4874),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4890),
.Y(n_4893)
);

OAI22xp5_ASAP7_75t_L g4894 ( 
.A1(n_4886),
.A2(n_2025),
.B1(n_1855),
.B2(n_1869),
.Y(n_4894)
);

OAI222xp33_ASAP7_75t_L g4895 ( 
.A1(n_4887),
.A2(n_1803),
.B1(n_1829),
.B2(n_1396),
.C1(n_1398),
.C2(n_1357),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4883),
.Y(n_4896)
);

INVx2_ASAP7_75t_L g4897 ( 
.A(n_4893),
.Y(n_4897)
);

XNOR2x1_ASAP7_75t_L g4898 ( 
.A(n_4896),
.B(n_4884),
.Y(n_4898)
);

XNOR2x1_ASAP7_75t_L g4899 ( 
.A(n_4894),
.B(n_4885),
.Y(n_4899)
);

INVxp67_ASAP7_75t_SL g4900 ( 
.A(n_4892),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_4895),
.Y(n_4901)
);

XNOR2x2_ASAP7_75t_L g4902 ( 
.A(n_4897),
.B(n_4889),
.Y(n_4902)
);

XNOR2xp5_ASAP7_75t_L g4903 ( 
.A(n_4900),
.B(n_4891),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4898),
.Y(n_4904)
);

AND3x4_ASAP7_75t_L g4905 ( 
.A(n_4901),
.B(n_1845),
.C(n_2008),
.Y(n_4905)
);

OAI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4904),
.A2(n_4899),
.B1(n_1869),
.B2(n_1879),
.Y(n_4906)
);

CKINVDCx20_ASAP7_75t_R g4907 ( 
.A(n_4903),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4905),
.A2(n_1845),
.B(n_2002),
.Y(n_4908)
);

OAI22xp5_ASAP7_75t_SL g4909 ( 
.A1(n_4902),
.A2(n_1839),
.B1(n_2002),
.B2(n_1995),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4907),
.B(n_1839),
.Y(n_4910)
);

AOI22xp5_ASAP7_75t_L g4911 ( 
.A1(n_4909),
.A2(n_1839),
.B1(n_1995),
.B2(n_1994),
.Y(n_4911)
);

AOI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4906),
.A2(n_1795),
.B1(n_1995),
.B2(n_1994),
.Y(n_4912)
);

AOI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4910),
.A2(n_4908),
.B(n_1869),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4912),
.B(n_4911),
.Y(n_4914)
);

XNOR2xp5_ASAP7_75t_L g4915 ( 
.A(n_4910),
.B(n_1825),
.Y(n_4915)
);

OA22x2_ASAP7_75t_L g4916 ( 
.A1(n_4911),
.A2(n_1825),
.B1(n_1961),
.B2(n_1957),
.Y(n_4916)
);

AOI222xp33_ASAP7_75t_SL g4917 ( 
.A1(n_4915),
.A2(n_1825),
.B1(n_1961),
.B2(n_1957),
.C1(n_1947),
.C2(n_1944),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4916),
.Y(n_4918)
);

XNOR2xp5_ASAP7_75t_L g4919 ( 
.A(n_4913),
.B(n_1825),
.Y(n_4919)
);

BUFx6f_ASAP7_75t_L g4920 ( 
.A(n_4914),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4915),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4915),
.Y(n_4922)
);

AOI222xp33_ASAP7_75t_L g4923 ( 
.A1(n_4915),
.A2(n_1994),
.B1(n_1961),
.B2(n_1957),
.C1(n_1947),
.C2(n_1944),
.Y(n_4923)
);

HB1xp67_ASAP7_75t_L g4924 ( 
.A(n_4915),
.Y(n_4924)
);

CKINVDCx20_ASAP7_75t_R g4925 ( 
.A(n_4914),
.Y(n_4925)
);

AOI22xp5_ASAP7_75t_SL g4926 ( 
.A1(n_4925),
.A2(n_1994),
.B1(n_1961),
.B2(n_1957),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_SL g4927 ( 
.A(n_4920),
.B(n_1947),
.Y(n_4927)
);

AOI22xp5_ASAP7_75t_SL g4928 ( 
.A1(n_4919),
.A2(n_1947),
.B1(n_1944),
.B2(n_1933),
.Y(n_4928)
);

OA22x2_ASAP7_75t_L g4929 ( 
.A1(n_4918),
.A2(n_1944),
.B1(n_1933),
.B2(n_1924),
.Y(n_4929)
);

NAND2xp33_ASAP7_75t_SL g4930 ( 
.A(n_4920),
.B(n_1795),
.Y(n_4930)
);

AND2x2_ASAP7_75t_L g4931 ( 
.A(n_4924),
.B(n_1795),
.Y(n_4931)
);

OAI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4921),
.A2(n_1803),
.B(n_1829),
.Y(n_4932)
);

OAI221xp5_ASAP7_75t_SL g4933 ( 
.A1(n_4922),
.A2(n_1791),
.B1(n_1924),
.B2(n_1916),
.C(n_1915),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_SL g4934 ( 
.A(n_4917),
.B(n_1791),
.Y(n_4934)
);

XNOR2xp5_ASAP7_75t_L g4935 ( 
.A(n_4931),
.B(n_4923),
.Y(n_4935)
);

HB1xp67_ASAP7_75t_L g4936 ( 
.A(n_4927),
.Y(n_4936)
);

AOI22x1_ASAP7_75t_L g4937 ( 
.A1(n_4932),
.A2(n_1791),
.B1(n_1924),
.B2(n_1916),
.Y(n_4937)
);

XNOR2xp5_ASAP7_75t_L g4938 ( 
.A(n_4930),
.B(n_1754),
.Y(n_4938)
);

NOR3xp33_ASAP7_75t_L g4939 ( 
.A(n_4934),
.B(n_1357),
.C(n_1387),
.Y(n_4939)
);

CKINVDCx14_ASAP7_75t_R g4940 ( 
.A(n_4928),
.Y(n_4940)
);

OR2x6_ASAP7_75t_L g4941 ( 
.A(n_4936),
.B(n_4929),
.Y(n_4941)
);

AOI221xp5_ASAP7_75t_L g4942 ( 
.A1(n_4940),
.A2(n_4933),
.B1(n_4926),
.B2(n_1791),
.C(n_1869),
.Y(n_4942)
);

AOI221xp5_ASAP7_75t_L g4943 ( 
.A1(n_4939),
.A2(n_1741),
.B1(n_1916),
.B2(n_1915),
.C(n_1906),
.Y(n_4943)
);

AOI21xp5_ASAP7_75t_L g4944 ( 
.A1(n_4941),
.A2(n_4935),
.B(n_4938),
.Y(n_4944)
);

AOI22xp5_ASAP7_75t_L g4945 ( 
.A1(n_4944),
.A2(n_4942),
.B1(n_4943),
.B2(n_4937),
.Y(n_4945)
);


endmodule