module fake_jpeg_7735_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_45),
.Y(n_50)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_24),
.B1(n_35),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_20),
.B1(n_28),
.B2(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_37),
.B1(n_24),
.B2(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_18),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_34),
.B1(n_32),
.B2(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_82),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_96),
.B1(n_32),
.B2(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_28),
.B1(n_65),
.B2(n_44),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_20),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_29),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_90),
.Y(n_125)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_106),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_29),
.B(n_31),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_111),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_56),
.C(n_57),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_64),
.C(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_97),
.B1(n_28),
.B2(n_50),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_38),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_36),
.C(n_42),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_130),
.C(n_131),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_135),
.B1(n_143),
.B2(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_41),
.C(n_42),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_41),
.C(n_42),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_104),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_153),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_97),
.B1(n_53),
.B2(n_93),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_121),
.B1(n_123),
.B2(n_93),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_144),
.B1(n_115),
.B2(n_123),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_41),
.C(n_45),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_106),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_31),
.B(n_30),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_115),
.B(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_53),
.B1(n_45),
.B2(n_38),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_38),
.B1(n_21),
.B2(n_26),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_148),
.B1(n_124),
.B2(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_33),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_150),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_21),
.B1(n_26),
.B2(n_23),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_33),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_45),
.B1(n_21),
.B2(n_26),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_19),
.B(n_17),
.C(n_16),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_17),
.B(n_19),
.C(n_118),
.Y(n_172)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_108),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_166),
.C(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_175),
.B1(n_176),
.B2(n_180),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_110),
.B1(n_104),
.B2(n_125),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_185),
.B1(n_138),
.B2(n_142),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_181),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_17),
.B(n_19),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_183),
.B(n_150),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_144),
.B1(n_152),
.B2(n_128),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_145),
.B1(n_136),
.B2(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_124),
.B1(n_120),
.B2(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_147),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_124),
.B1(n_120),
.B2(n_21),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_26),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_23),
.B1(n_33),
.B2(n_25),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_78),
.B1(n_21),
.B2(n_23),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_172),
.B1(n_173),
.B2(n_159),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_139),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_199),
.C(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_201),
.B(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_207),
.B1(n_17),
.B2(n_29),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_86),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_203),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_23),
.B1(n_33),
.B2(n_25),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_154),
.B1(n_113),
.B2(n_72),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_183),
.B1(n_158),
.B2(n_117),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_77),
.B1(n_72),
.B2(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_188),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_0),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_0),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_185),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_1),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_221),
.C(n_224),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_160),
.C(n_159),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_117),
.C(n_77),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_19),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_19),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_19),
.C(n_17),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_240),
.Y(n_259)
);

OAI22x1_ASAP7_75t_SL g237 ( 
.A1(n_188),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_201),
.C(n_212),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_29),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_210),
.C(n_211),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_242),
.B(n_250),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_202),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_196),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_239),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_195),
.Y(n_247)
);

XOR2x2_ASAP7_75t_SL g250 ( 
.A(n_230),
.B(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_214),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_216),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_254),
.A2(n_7),
.B(n_15),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_195),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_245),
.C(n_263),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_223),
.B1(n_222),
.B2(n_218),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_225),
.B1(n_238),
.B2(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_270),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_229),
.C(n_226),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_205),
.B1(n_193),
.B2(n_215),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_280),
.B1(n_249),
.B2(n_9),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_246),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_205),
.B(n_194),
.C(n_233),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_275),
.B1(n_281),
.B2(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_244),
.B1(n_255),
.B2(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_9),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_297),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_250),
.C(n_242),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_6),
.B(n_15),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_257),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_296),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_270),
.C(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_276),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_11),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_271),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_299),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_279),
.B1(n_249),
.B2(n_11),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_6),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_1),
.C(n_2),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_286),
.B(n_12),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_14),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_320),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_290),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_294),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_299),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_321),
.A2(n_327),
.B(n_284),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_298),
.C(n_300),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_288),
.B(n_14),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_284),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_305),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_313),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_332),
.Y(n_333)
);

A2O1A1O1Ixp25_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_323),
.B(n_322),
.C(n_4),
.D(n_5),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.C(n_3),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_338)
);

AOI221xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_4),
.B1(n_5),
.B2(n_29),
.C(n_335),
.Y(n_339)
);


endmodule