module real_aes_8871_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g532 ( .A(n_1), .Y(n_532) );
INVx1_ASAP7_75t_L g197 ( .A(n_2), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_3), .A2(n_38), .B1(n_159), .B2(n_474), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g138 ( .A1(n_4), .A2(n_139), .B(n_146), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_5), .B(n_132), .Y(n_523) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_7), .A2(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_39), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_8), .B(n_39), .Y(n_448) );
INVx1_ASAP7_75t_L g156 ( .A(n_9), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_10), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g137 ( .A(n_11), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_12), .B(n_169), .Y(n_469) );
INVx1_ASAP7_75t_L g244 ( .A(n_13), .Y(n_244) );
INVx1_ASAP7_75t_L g527 ( .A(n_14), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_15), .B(n_133), .Y(n_508) );
AO32x2_ASAP7_75t_L g489 ( .A1(n_16), .A2(n_132), .A3(n_166), .B1(n_490), .B2(n_494), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_17), .B(n_159), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_18), .B(n_185), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_19), .B(n_133), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_20), .A2(n_49), .B1(n_159), .B2(n_474), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_21), .B(n_139), .Y(n_209) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_22), .A2(n_74), .B1(n_159), .B2(n_169), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_23), .B(n_159), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_24), .B(n_130), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_25), .A2(n_242), .B(n_243), .C(n_245), .Y(n_241) );
OAI222xp33_ASAP7_75t_L g453 ( .A1(n_26), .A2(n_454), .B1(n_741), .B2(n_747), .C1(n_748), .C2(n_750), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_26), .Y(n_747) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_27), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_28), .B(n_162), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_29), .B(n_154), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_30), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_31), .Y(n_750) );
INVx1_ASAP7_75t_L g175 ( .A(n_32), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_33), .B(n_162), .Y(n_487) );
INVx2_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_35), .B(n_159), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_36), .B(n_162), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_37), .A2(n_144), .B(n_149), .C(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g173 ( .A(n_40), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_41), .B(n_154), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_42), .B(n_159), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_43), .A2(n_84), .B1(n_216), .B2(n_474), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_44), .B(n_159), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_45), .B(n_159), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_46), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_47), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_48), .B(n_139), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_50), .A2(n_59), .B1(n_159), .B2(n_169), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_51), .A2(n_149), .B1(n_169), .B2(n_171), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_52), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_53), .B(n_159), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_54), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_55), .B(n_159), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_56), .A2(n_153), .B(n_155), .C(n_158), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_57), .Y(n_262) );
INVx1_ASAP7_75t_L g147 ( .A(n_58), .Y(n_147) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_61), .A2(n_120), .B1(n_121), .B2(n_440), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_61), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_62), .B(n_159), .Y(n_533) );
INVx1_ASAP7_75t_L g136 ( .A(n_63), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
AO32x2_ASAP7_75t_L g499 ( .A1(n_65), .A2(n_132), .A3(n_224), .B1(n_494), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g544 ( .A(n_66), .Y(n_544) );
INVx1_ASAP7_75t_L g482 ( .A(n_67), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_SL g184 ( .A1(n_68), .A2(n_158), .B(n_185), .C(n_186), .Y(n_184) );
INVxp67_ASAP7_75t_L g187 ( .A(n_69), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_70), .B(n_169), .Y(n_483) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_72), .Y(n_179) );
INVx1_ASAP7_75t_L g255 ( .A(n_73), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_75), .A2(n_144), .B(n_149), .C(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_76), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_77), .B(n_169), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_78), .B(n_198), .Y(n_212) );
INVx2_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_80), .B(n_185), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_81), .B(n_169), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_82), .A2(n_144), .B(n_149), .C(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
OR2x2_ASAP7_75t_L g445 ( .A(n_83), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g456 ( .A(n_83), .B(n_447), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_85), .A2(n_98), .B1(n_169), .B2(n_170), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_86), .B(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_87), .A2(n_100), .B1(n_113), .B2(n_754), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_88), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_89), .A2(n_144), .B(n_149), .C(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_90), .Y(n_234) );
INVx1_ASAP7_75t_L g183 ( .A(n_91), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_92), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_93), .B(n_198), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_94), .B(n_169), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_95), .B(n_132), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_97), .A2(n_139), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_SL g754 ( .A(n_102), .Y(n_754) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g447 ( .A(n_108), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g458 ( .A(n_109), .B(n_447), .Y(n_458) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_109), .B(n_446), .Y(n_749) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_452), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g753 ( .A(n_116), .Y(n_753) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_442), .B(n_449), .Y(n_118) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_123), .A2(n_455), .B1(n_457), .B2(n_459), .Y(n_454) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g441 ( .A(n_124), .Y(n_441) );
AND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_362), .C(n_407), .Y(n_124) );
NOR4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_285), .C(n_326), .D(n_343), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_189), .B(n_205), .C(n_247), .Y(n_126) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_128), .B(n_190), .Y(n_189) );
NOR4xp25_ASAP7_75t_L g309 ( .A(n_128), .B(n_303), .C(n_310), .D(n_316), .Y(n_309) );
AND2x2_ASAP7_75t_L g382 ( .A(n_128), .B(n_271), .Y(n_382) );
AND2x2_ASAP7_75t_L g401 ( .A(n_128), .B(n_347), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_128), .B(n_396), .Y(n_410) );
AND2x2_ASAP7_75t_L g423 ( .A(n_128), .B(n_204), .Y(n_423) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_SL g268 ( .A(n_129), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_129), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g325 ( .A(n_129), .B(n_164), .Y(n_325) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_129), .B(n_271), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_129), .B(n_164), .Y(n_340) );
AND2x2_ASAP7_75t_L g349 ( .A(n_129), .B(n_274), .Y(n_349) );
BUFx2_ASAP7_75t_L g372 ( .A(n_129), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_129), .B(n_180), .Y(n_376) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_138), .B(n_161), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_131), .B(n_219), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_131), .B(n_494), .C(n_510), .Y(n_509) );
AO21x1_ASAP7_75t_L g547 ( .A1(n_131), .A2(n_510), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_132), .A2(n_181), .B(n_188), .Y(n_180) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_132), .A2(n_515), .B(n_523), .Y(n_514) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_134), .B(n_135), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx2_ASAP7_75t_L g238 ( .A(n_139), .Y(n_238) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_140), .B(n_144), .Y(n_177) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g522 ( .A(n_141), .Y(n_522) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
INVx1_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
INVx1_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_143), .Y(n_157) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
INVx4_ASAP7_75t_SL g160 ( .A(n_144), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_144), .A2(n_467), .B(n_471), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_144), .A2(n_481), .B(n_484), .Y(n_480) );
BUFx3_ASAP7_75t_L g494 ( .A(n_144), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_144), .A2(n_516), .B(n_519), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_144), .A2(n_526), .B(n_530), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_152), .C(n_160), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_148), .A2(n_160), .B(n_183), .C(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_148), .A2(n_160), .B(n_240), .C(n_241), .Y(n_239) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx3_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g474 ( .A(n_150), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_153), .A2(n_472), .B(n_473), .Y(n_471) );
O2A1O1Ixp5_ASAP7_75t_L g543 ( .A1(n_153), .A2(n_531), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx4_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_154), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g500 ( .A1(n_154), .A2(n_157), .B1(n_501), .B2(n_502), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_154), .A2(n_492), .B1(n_511), .B2(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_157), .B(n_187), .Y(n_186) );
INVx5_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_SL g481 ( .A1(n_158), .A2(n_198), .B(n_482), .C(n_483), .Y(n_481) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_159), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g167 ( .A1(n_160), .A2(n_168), .B1(n_176), .B2(n_177), .Y(n_167) );
INVx1_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx2_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_162), .A2(n_237), .B(n_246), .Y(n_236) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_162), .A2(n_466), .B(n_475), .Y(n_465) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_162), .A2(n_480), .B(n_487), .Y(n_479) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
AND2x2_ASAP7_75t_L g204 ( .A(n_164), .B(n_180), .Y(n_204) );
BUFx2_ASAP7_75t_L g278 ( .A(n_164), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_164), .A2(n_311), .B1(n_313), .B2(n_314), .Y(n_310) );
OR2x2_ASAP7_75t_L g332 ( .A(n_164), .B(n_192), .Y(n_332) );
AND2x2_ASAP7_75t_L g396 ( .A(n_164), .B(n_274), .Y(n_396) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g264 ( .A(n_165), .B(n_192), .Y(n_264) );
AND2x2_ASAP7_75t_L g271 ( .A(n_165), .B(n_180), .Y(n_271) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_165), .Y(n_313) );
OR2x2_ASAP7_75t_L g348 ( .A(n_165), .B(n_191), .Y(n_348) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_178), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_166), .B(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_166), .A2(n_193), .B(n_201), .Y(n_192) );
INVx2_ASAP7_75t_L g217 ( .A(n_166), .Y(n_217) );
INVx2_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g174 ( .A(n_172), .Y(n_174) );
INVx4_ASAP7_75t_L g242 ( .A(n_172), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_177), .A2(n_194), .B(n_195), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_177), .A2(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g267 ( .A(n_180), .Y(n_267) );
INVx3_ASAP7_75t_L g276 ( .A(n_180), .Y(n_276) );
BUFx2_ASAP7_75t_L g300 ( .A(n_180), .Y(n_300) );
AND2x2_ASAP7_75t_L g333 ( .A(n_180), .B(n_268), .Y(n_333) );
INVx1_ASAP7_75t_L g470 ( .A(n_185), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_189), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_418) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_204), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_191), .B(n_276), .Y(n_280) );
INVx1_ASAP7_75t_L g308 ( .A(n_191), .Y(n_308) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g274 ( .A(n_192), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .C(n_200), .Y(n_196) );
INVx2_ASAP7_75t_L g492 ( .A(n_198), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_198), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_198), .A2(n_541), .B(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_200), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_203), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_203), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
NAND2x1_ASAP7_75t_SL g205 ( .A(n_206), .B(n_220), .Y(n_205) );
AND2x2_ASAP7_75t_L g284 ( .A(n_206), .B(n_235), .Y(n_284) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_206), .Y(n_358) );
AND2x2_ASAP7_75t_L g385 ( .A(n_206), .B(n_305), .Y(n_385) );
AND2x2_ASAP7_75t_L g393 ( .A(n_206), .B(n_355), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_206), .B(n_250), .Y(n_420) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g251 ( .A(n_207), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g269 ( .A(n_207), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
INVx1_ASAP7_75t_L g296 ( .A(n_207), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_207), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_207), .B(n_253), .Y(n_329) );
OR2x2_ASAP7_75t_L g367 ( .A(n_207), .B(n_322), .Y(n_367) );
AOI32xp33_ASAP7_75t_L g379 ( .A1(n_207), .A2(n_380), .A3(n_383), .B1(n_384), .B2(n_385), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_207), .B(n_355), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_207), .B(n_315), .Y(n_430) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_210), .B(n_217), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_214), .A2(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g245 ( .A(n_216), .Y(n_245) );
INVx1_ASAP7_75t_L g260 ( .A(n_217), .Y(n_260) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_217), .A2(n_525), .B(n_534), .Y(n_524) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_217), .A2(n_539), .B(n_546), .Y(n_538) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g341 ( .A(n_221), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
INVx1_ASAP7_75t_L g303 ( .A(n_222), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_222), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_222), .B(n_252), .Y(n_322) );
AND2x2_ASAP7_75t_L g355 ( .A(n_222), .B(n_331), .Y(n_355) );
AND2x2_ASAP7_75t_L g392 ( .A(n_222), .B(n_253), .Y(n_392) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_223), .B(n_252), .Y(n_282) );
AND2x2_ASAP7_75t_L g289 ( .A(n_223), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g330 ( .A(n_223), .B(n_331), .Y(n_330) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_231), .Y(n_227) );
INVx2_ASAP7_75t_L g306 ( .A(n_235), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_235), .B(n_252), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_235), .B(n_297), .Y(n_378) );
INVx1_ASAP7_75t_L g400 ( .A(n_235), .Y(n_400) );
INVx1_ASAP7_75t_L g417 ( .A(n_235), .Y(n_417) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g270 ( .A(n_236), .B(n_252), .Y(n_270) );
AND2x2_ASAP7_75t_L g292 ( .A(n_236), .B(n_253), .Y(n_292) );
INVx1_ASAP7_75t_L g331 ( .A(n_236), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_242), .B(n_244), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_242), .A2(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g529 ( .A(n_242), .Y(n_529) );
AOI221x1_ASAP7_75t_SL g247 ( .A1(n_248), .A2(n_263), .B1(n_269), .B2(n_271), .C(n_272), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_248), .A2(n_336), .B1(n_403), .B2(n_404), .Y(n_402) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND2x2_ASAP7_75t_L g294 ( .A(n_249), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g389 ( .A(n_249), .B(n_269), .Y(n_389) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g345 ( .A(n_250), .B(n_270), .Y(n_345) );
INVx1_ASAP7_75t_L g357 ( .A(n_251), .Y(n_357) );
AND2x2_ASAP7_75t_L g368 ( .A(n_251), .B(n_355), .Y(n_368) );
AND2x2_ASAP7_75t_L g435 ( .A(n_251), .B(n_330), .Y(n_435) );
INVx2_ASAP7_75t_L g297 ( .A(n_252), .Y(n_297) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_260), .B(n_261), .Y(n_253) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_264), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_265), .B(n_348), .Y(n_351) );
INVx3_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_266), .A2(n_387), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NOR2xp33_ASAP7_75t_SL g409 ( .A(n_269), .B(n_295), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_270), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g361 ( .A(n_270), .B(n_289), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_270), .B(n_296), .Y(n_438) );
AND2x2_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g374 ( .A(n_271), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B(n_281), .Y(n_272) );
NAND2x1_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_274), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g323 ( .A(n_274), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g335 ( .A(n_274), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_274), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g359 ( .A(n_275), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_275), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_275), .B(n_278), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_278), .A2(n_317), .B(n_347), .C(n_349), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_278), .A2(n_365), .B1(n_368), .B2(n_369), .C(n_373), .Y(n_364) );
AND2x2_ASAP7_75t_L g360 ( .A(n_279), .B(n_313), .Y(n_360) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g320 ( .A(n_284), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g391 ( .A(n_284), .B(n_392), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_293), .C(n_318), .Y(n_285) );
NAND3xp33_ASAP7_75t_SL g404 ( .A(n_286), .B(n_405), .C(n_406), .Y(n_404) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
OR2x2_ASAP7_75t_L g377 ( .A(n_288), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .B1(n_301), .B2(n_307), .C(n_309), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_295), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_300), .A2(n_357), .B1(n_358), .B2(n_359), .Y(n_356) );
OR2x2_ASAP7_75t_L g437 ( .A(n_300), .B(n_348), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVxp67_ASAP7_75t_L g411 ( .A(n_303), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_305), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g312 ( .A(n_306), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_308), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_308), .B(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_308), .B(n_375), .Y(n_414) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g428 ( .A(n_317), .B(n_348), .Y(n_428) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g406 ( .A(n_323), .Y(n_406) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI322xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_332), .A3(n_333), .B1(n_334), .B2(n_337), .C1(n_339), .C2(n_341), .Y(n_326) );
OAI322xp33_ASAP7_75t_L g408 ( .A1(n_327), .A2(n_409), .A3(n_410), .B1(n_411), .B2(n_412), .C1(n_413), .C2(n_415), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx4_ASAP7_75t_L g342 ( .A(n_329), .Y(n_342) );
AND2x2_ASAP7_75t_L g403 ( .A(n_329), .B(n_355), .Y(n_403) );
AND2x2_ASAP7_75t_L g416 ( .A(n_329), .B(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_332), .Y(n_427) );
INVx1_ASAP7_75t_L g405 ( .A(n_333), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OR2x2_ASAP7_75t_L g339 ( .A(n_335), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g422 ( .A(n_335), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_335), .B(n_376), .Y(n_433) );
OR2x2_ASAP7_75t_L g366 ( .A(n_338), .B(n_367), .Y(n_366) );
INVxp33_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
OAI221xp5_ASAP7_75t_SL g343 ( .A1(n_342), .A2(n_344), .B1(n_346), .B2(n_350), .C(n_352), .Y(n_343) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_342), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g426 ( .A(n_342), .Y(n_426) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI322xp5_ASAP7_75t_L g390 ( .A1(n_349), .A2(n_374), .A3(n_391), .B1(n_393), .B2(n_394), .C1(n_397), .C2(n_401), .Y(n_390) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B1(n_360), .B2(n_361), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_386), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_364), .B(n_379), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_367), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NAND2xp33_ASAP7_75t_SL g384 ( .A(n_370), .B(n_381), .Y(n_384) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OAI322xp33_ASAP7_75t_L g424 ( .A1(n_372), .A2(n_425), .A3(n_427), .B1(n_428), .B2(n_429), .C1(n_431), .C2(n_434), .Y(n_424) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_382), .B(n_430), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_388), .B(n_390), .C(n_402), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_418), .C(n_424), .D(n_436), .Y(n_407) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_441), .A2(n_742), .B1(n_745), .B2(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_449), .A2(n_453), .B(n_751), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g744 ( .A(n_456), .Y(n_744) );
INVx6_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g745 ( .A(n_458), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_459), .Y(n_746) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_663), .Y(n_459) );
NAND5xp2_ASAP7_75t_L g460 ( .A(n_461), .B(n_582), .C(n_597), .D(n_623), .E(n_645), .Y(n_460) );
NOR2xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_562), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_503), .B1(n_535), .B2(n_551), .C(n_552), .Y(n_462) );
NOR2xp33_ASAP7_75t_SL g463 ( .A(n_464), .B(n_495), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_464), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g739 ( .A(n_464), .Y(n_739) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
INVx1_ASAP7_75t_L g579 ( .A(n_465), .Y(n_579) );
AND2x2_ASAP7_75t_L g581 ( .A(n_465), .B(n_489), .Y(n_581) );
AND2x2_ASAP7_75t_L g591 ( .A(n_465), .B(n_488), .Y(n_591) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_465), .Y(n_609) );
INVx1_ASAP7_75t_L g619 ( .A(n_465), .Y(n_619) );
OR2x2_ASAP7_75t_L g657 ( .A(n_465), .B(n_556), .Y(n_657) );
INVx2_ASAP7_75t_L g707 ( .A(n_465), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_465), .B(n_555), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_470), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_477), .B(n_488), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_478), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_478), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_478), .B(n_579), .Y(n_639) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_479), .Y(n_497) );
INVx2_ASAP7_75t_L g556 ( .A(n_479), .Y(n_556) );
OR2x2_ASAP7_75t_L g618 ( .A(n_479), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g557 ( .A(n_488), .B(n_499), .Y(n_557) );
AND2x2_ASAP7_75t_L g574 ( .A(n_488), .B(n_554), .Y(n_574) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g498 ( .A(n_489), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g577 ( .A(n_489), .Y(n_577) );
AND2x2_ASAP7_75t_L g706 ( .A(n_489), .B(n_707), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_492), .A2(n_520), .B(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_492), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_494), .A2(n_540), .B(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
AND2x2_ASAP7_75t_L g669 ( .A(n_496), .B(n_557), .Y(n_669) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g670 ( .A(n_497), .B(n_581), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_498), .A2(n_638), .B(n_640), .C(n_642), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_498), .B(n_638), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_498), .A2(n_568), .B1(n_711), .B2(n_712), .C(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
INVx1_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_499), .Y(n_599) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
AND2x2_ASAP7_75t_L g616 ( .A(n_505), .B(n_561), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_505), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_506), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g708 ( .A(n_506), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g740 ( .A(n_506), .Y(n_740) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
AND2x2_ASAP7_75t_L g596 ( .A(n_507), .B(n_550), .Y(n_596) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_507), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g612 ( .A(n_507), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_513), .B(n_652), .Y(n_687) );
INVx1_ASAP7_75t_SL g691 ( .A(n_513), .Y(n_691) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
INVx3_ASAP7_75t_L g550 ( .A(n_514), .Y(n_550) );
AND2x2_ASAP7_75t_L g561 ( .A(n_514), .B(n_538), .Y(n_561) );
AND2x2_ASAP7_75t_L g583 ( .A(n_514), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_622), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_514), .B(n_560), .Y(n_709) );
INVx2_ASAP7_75t_L g531 ( .A(n_522), .Y(n_531) );
AND2x2_ASAP7_75t_L g549 ( .A(n_524), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g560 ( .A(n_524), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_524), .B(n_538), .Y(n_585) );
AND2x2_ASAP7_75t_L g621 ( .A(n_524), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_549), .Y(n_536) );
INVx1_ASAP7_75t_L g601 ( .A(n_537), .Y(n_601) );
AND2x2_ASAP7_75t_L g643 ( .A(n_537), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_537), .B(n_564), .Y(n_649) );
AOI21xp5_ASAP7_75t_SL g723 ( .A1(n_537), .A2(n_555), .B(n_578), .Y(n_723) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
OR2x2_ASAP7_75t_L g566 ( .A(n_538), .B(n_547), .Y(n_566) );
AND2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_550), .Y(n_613) );
INVx2_ASAP7_75t_L g622 ( .A(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g728 ( .A(n_538), .Y(n_728) );
AND2x2_ASAP7_75t_L g652 ( .A(n_547), .B(n_622), .Y(n_652) );
INVx1_ASAP7_75t_L g677 ( .A(n_547), .Y(n_677) );
AND2x2_ASAP7_75t_L g586 ( .A(n_549), .B(n_570), .Y(n_586) );
AND2x2_ASAP7_75t_L g598 ( .A(n_549), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g716 ( .A(n_549), .Y(n_716) );
INVx2_ASAP7_75t_L g606 ( .A(n_550), .Y(n_606) );
AND2x2_ASAP7_75t_L g644 ( .A(n_550), .B(n_560), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_550), .B(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_557), .B(n_558), .Y(n_552) );
AND2x2_ASAP7_75t_L g659 ( .A(n_553), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g713 ( .A(n_553), .Y(n_713) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
BUFx2_ASAP7_75t_L g732 ( .A(n_554), .Y(n_732) );
BUFx2_ASAP7_75t_L g603 ( .A(n_555), .Y(n_603) );
AND2x2_ASAP7_75t_L g705 ( .A(n_555), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g688 ( .A(n_556), .Y(n_688) );
AND2x4_ASAP7_75t_L g615 ( .A(n_557), .B(n_578), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_557), .B(n_639), .Y(n_651) );
AOI32xp33_ASAP7_75t_L g575 ( .A1(n_558), .A2(n_576), .A3(n_578), .B1(n_580), .B2(n_581), .Y(n_575) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx3_ASAP7_75t_L g564 ( .A(n_559), .Y(n_564) );
OR2x2_ASAP7_75t_L g700 ( .A(n_559), .B(n_656), .Y(n_700) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g569 ( .A(n_560), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g676 ( .A(n_560), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g568 ( .A(n_561), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_561), .B(n_570), .Y(n_580) );
INVx1_ASAP7_75t_L g701 ( .A(n_561), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_561), .B(n_676), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_567), .B(n_571), .C(n_575), .Y(n_562) );
OAI322xp33_ASAP7_75t_L g671 ( .A1(n_563), .A2(n_608), .A3(n_672), .B1(n_674), .B2(n_678), .C1(n_679), .C2(n_683), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVxp67_ASAP7_75t_L g636 ( .A(n_564), .Y(n_636) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g690 ( .A(n_566), .B(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_566), .B(n_606), .Y(n_737) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g629 ( .A(n_569), .Y(n_629) );
OR2x2_ASAP7_75t_L g715 ( .A(n_570), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_573), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g624 ( .A(n_574), .B(n_603), .Y(n_624) );
AND2x2_ASAP7_75t_L g695 ( .A(n_574), .B(n_608), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_574), .B(n_682), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_576), .A2(n_583), .B1(n_586), .B2(n_587), .C(n_592), .Y(n_582) );
OR2x2_ASAP7_75t_L g593 ( .A(n_576), .B(n_589), .Y(n_593) );
AND2x2_ASAP7_75t_L g681 ( .A(n_576), .B(n_682), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g720 ( .A1(n_576), .A2(n_606), .A3(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_577), .B(n_613), .C(n_636), .Y(n_654) );
AND2x2_ASAP7_75t_L g680 ( .A(n_577), .B(n_673), .Y(n_680) );
INVxp67_ASAP7_75t_L g660 ( .A(n_578), .Y(n_660) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_581), .B(n_633), .Y(n_689) );
INVx2_ASAP7_75t_L g699 ( .A(n_581), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_581), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g668 ( .A(n_584), .Y(n_668) );
OR2x2_ASAP7_75t_L g594 ( .A(n_585), .B(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_587), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_590), .Y(n_673) );
AND2x2_ASAP7_75t_L g632 ( .A(n_591), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g678 ( .A(n_591), .Y(n_678) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_591), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AOI21xp33_ASAP7_75t_SL g617 ( .A1(n_593), .A2(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g711 ( .A(n_596), .B(n_621), .Y(n_711) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_610), .C(n_617), .Y(n_597) );
AND2x2_ASAP7_75t_L g641 ( .A(n_599), .B(n_609), .Y(n_641) );
INVx2_ASAP7_75t_L g656 ( .A(n_599), .Y(n_656) );
OR2x2_ASAP7_75t_L g694 ( .A(n_599), .B(n_657), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_599), .B(n_737), .Y(n_736) );
AOI211xp5_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_602), .B(n_604), .C(n_607), .Y(n_600) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_603), .B(n_641), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_604), .A2(n_699), .B(n_723), .C(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_605), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g662 ( .A(n_606), .B(n_652), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_606), .Y(n_667) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVxp33_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
AND2x2_ASAP7_75t_L g697 ( .A(n_613), .B(n_676), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_618), .A2(n_680), .B(n_681), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g698 ( .A1(n_620), .A2(n_699), .A3(n_700), .B1(n_701), .B2(n_702), .C1(n_704), .C2(n_708), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_630), .B2(n_634), .C(n_637), .Y(n_623) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g675 ( .A(n_628), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g719 ( .A(n_632), .Y(n_719) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_635), .B(n_655), .Y(n_721) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g684 ( .A(n_644), .B(n_652), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_652), .C(n_653), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_648), .A2(n_665), .B1(n_669), .B2(n_670), .C(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_652), .B(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_658), .B2(n_661), .Y(n_653) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_SL g682 ( .A(n_657), .Y(n_682) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_685), .C(n_710), .D(n_720), .E(n_730), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_668), .Y(n_665) );
NOR4xp25_ASAP7_75t_L g738 ( .A(n_667), .B(n_673), .C(n_739), .D(n_740), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_670), .A2(n_731), .B1(n_733), .B2(n_735), .C(n_738), .Y(n_730) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g729 ( .A(n_676), .Y(n_729) );
OAI322xp33_ASAP7_75t_L g686 ( .A1(n_680), .A2(n_687), .A3(n_688), .B1(n_689), .B2(n_690), .C1(n_692), .C2(n_696), .Y(n_686) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_698), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g731 ( .A(n_706), .B(n_732), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
endmodule