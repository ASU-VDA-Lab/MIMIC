module fake_jpeg_227_n_58 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_58);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_16),
.B(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_17),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_18),
.C(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_18),
.C(n_4),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_18),
.B(n_1),
.C(n_2),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_0),
.C(n_3),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_0),
.C(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_40),
.B1(n_6),
.B2(n_7),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_5),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_49),
.B1(n_9),
.B2(n_12),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_5),
.C(n_6),
.Y(n_53)
);

OAI321xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_52),
.B2(n_49),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_53),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_12),
.Y(n_58)
);


endmodule