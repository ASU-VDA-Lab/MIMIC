module fake_netlist_6_1876_n_1246 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1246);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1246;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_95),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_54),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_44),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_21),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_66),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_55),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_125),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_148),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_63),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_116),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_76),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_163),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_47),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_56),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_31),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_84),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_74),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_86),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_152),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_57),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_78),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_104),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_138),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_45),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_33),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_83),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_179),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_161),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_131),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_181),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_166),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_184),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_132),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_158),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_19),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_121),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_105),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_80),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_72),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_114),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_107),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_29),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_119),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_96),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_43),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_106),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_6),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_128),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_43),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_44),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_130),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_162),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_67),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_174),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_35),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_120),
.Y(n_308)
);

BUFx2_ASAP7_75t_SL g309 ( 
.A(n_180),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_108),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_19),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_269),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_256),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_193),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_232),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_194),
.B(n_1),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_200),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_193),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_191),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_200),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_231),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_222),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_197),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_194),
.B(n_2),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_207),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_211),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_287),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_289),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_233),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_289),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_231),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_307),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_196),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_207),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_307),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_201),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_198),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_214),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_240),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_213),
.B(n_3),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_221),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_219),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_219),
.Y(n_365)
);

BUFx6f_ASAP7_75t_SL g366 ( 
.A(n_282),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_263),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_224),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_213),
.B(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_209),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_228),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_238),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_212),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_252),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_254),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_215),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_255),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_247),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_263),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_216),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_258),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_276),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_273),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_280),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_276),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_286),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_286),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_281),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_295),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_285),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_295),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_217),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_282),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_220),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_304),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_195),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_195),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_327),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_364),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_334),
.B(n_202),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_333),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_R g414 ( 
.A(n_349),
.B(n_225),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_364),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_356),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_354),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_358),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_370),
.Y(n_423)
);

CKINVDCx8_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_332),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_371),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_376),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_309),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_379),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_344),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_321),
.B(n_282),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_365),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_383),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_396),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_325),
.A2(n_283),
.B1(n_270),
.B2(n_291),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

NOR2x1_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_245),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_350),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_314),
.B(n_245),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_326),
.B(n_331),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_365),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_316),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_366),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_330),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_334),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_366),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_319),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_357),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_318),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_440),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_288),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_346),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_420),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_468),
.B(n_322),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_406),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_206),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_468),
.B(n_463),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_429),
.B(n_400),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_444),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_416),
.B(n_381),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_418),
.B(n_312),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_404),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_426),
.B(n_324),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_335),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_428),
.B(n_288),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_322),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_414),
.B(n_453),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_339),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_444),
.Y(n_507)
);

NOR2x1p5_ASAP7_75t_L g508 ( 
.A(n_467),
.B(n_244),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_405),
.B(n_336),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_437),
.B(n_362),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_441),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_438),
.A2(n_439),
.B1(n_448),
.B2(n_443),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_406),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_347),
.B1(n_341),
.B2(n_353),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_226),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_454),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_229),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_403),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_433),
.B(n_206),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_202),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_453),
.B(n_203),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_464),
.B(n_203),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_467),
.B(n_204),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_433),
.A2(n_253),
.B1(n_293),
.B2(n_294),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_469),
.B(n_234),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_460),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_431),
.A2(n_351),
.B1(n_352),
.B2(n_218),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_431),
.A2(n_206),
.B1(n_218),
.B2(n_306),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_408),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_472),
.B(n_204),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_471),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_412),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_516),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_479),
.B(n_412),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_417),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_475),
.B(n_417),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_518),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_502),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_502),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_516),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_476),
.A2(n_503),
.B1(n_475),
.B2(n_518),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_421),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_495),
.B(n_421),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_517),
.B(n_423),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_503),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_482),
.B(n_447),
.C(n_422),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_423),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_433),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_498),
.B(n_430),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_497),
.B(n_430),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_473),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_432),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_524),
.B(n_432),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_525),
.B(n_435),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_525),
.B(n_435),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_476),
.B(n_466),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_476),
.A2(n_218),
.B1(n_206),
.B2(n_250),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_499),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_473),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_531),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_531),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_501),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_510),
.B(n_442),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_520),
.B(n_442),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_507),
.Y(n_582)
);

AOI221xp5_ASAP7_75t_SL g583 ( 
.A1(n_490),
.A2(n_218),
.B1(n_250),
.B2(n_306),
.C(n_456),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_532),
.B(n_445),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_474),
.B(n_445),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_474),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_518),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_466),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_478),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_491),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_477),
.B(n_433),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_541),
.B(n_446),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_504),
.B(n_446),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_532),
.B(n_250),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_406),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_494),
.B(n_235),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_494),
.B(n_237),
.Y(n_597)
);

AOI22x1_ASAP7_75t_L g598 ( 
.A1(n_484),
.A2(n_205),
.B1(n_208),
.B2(n_275),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_494),
.B(n_496),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_537),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_494),
.B(n_239),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_496),
.B(n_241),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_496),
.B(n_242),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_496),
.B(n_243),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_527),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_500),
.B(n_246),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_535),
.B(n_461),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_532),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_500),
.B(n_249),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_540),
.B(n_461),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_537),
.B(n_484),
.Y(n_615)
);

AO22x1_ASAP7_75t_L g616 ( 
.A1(n_476),
.A2(n_533),
.B1(n_503),
.B2(n_303),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_488),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_500),
.B(n_259),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_507),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_489),
.B(n_455),
.Y(n_622)
);

NAND2x1_ASAP7_75t_L g623 ( 
.A(n_480),
.B(n_481),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_521),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_488),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_521),
.A2(n_382),
.B1(n_395),
.B2(n_393),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_500),
.B(n_260),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_493),
.B(n_262),
.Y(n_630)
);

BUFx5_ASAP7_75t_L g631 ( 
.A(n_503),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_493),
.B(n_265),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_534),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_542),
.B(n_266),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_476),
.A2(n_503),
.B1(n_522),
.B2(n_530),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_515),
.A2(n_306),
.B(n_250),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_529),
.B(n_455),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_513),
.B(n_205),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_542),
.B(n_267),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_542),
.B(n_271),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_480),
.B(n_274),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_577),
.A2(n_615),
.B(n_589),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_577),
.A2(n_519),
.B(n_486),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_549),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_615),
.A2(n_486),
.B(n_484),
.Y(n_645)
);

BUFx4f_ASAP7_75t_L g646 ( 
.A(n_625),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_599),
.A2(n_486),
.B(n_505),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_618),
.Y(n_648)
);

OAI22x1_ASAP7_75t_L g649 ( 
.A1(n_544),
.A2(n_355),
.B1(n_325),
.B2(n_328),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_624),
.Y(n_650)
);

CKINVDCx10_ASAP7_75t_R g651 ( 
.A(n_571),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_582),
.A2(n_492),
.B(n_485),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_569),
.A2(n_526),
.B(n_534),
.C(n_521),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_554),
.A2(n_481),
.B(n_480),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_554),
.A2(n_481),
.B(n_480),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_611),
.A2(n_483),
.B(n_481),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_476),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_582),
.A2(n_492),
.B(n_485),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_556),
.B(n_513),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_641),
.A2(n_492),
.B(n_485),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_588),
.A2(n_521),
.B(n_530),
.C(n_512),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_578),
.A2(n_521),
.B(n_530),
.C(n_538),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_633),
.Y(n_665)
);

BUFx12f_ASAP7_75t_L g666 ( 
.A(n_581),
.Y(n_666)
);

BUFx6f_ASAP7_75t_SL g667 ( 
.A(n_564),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_549),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_575),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_546),
.A2(n_539),
.B(n_508),
.C(n_483),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_596),
.A2(n_492),
.B(n_485),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_556),
.B(n_483),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_547),
.B(n_489),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_592),
.B(n_483),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_634),
.A2(n_640),
.B(n_639),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_593),
.B(n_424),
.C(n_434),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_592),
.B(n_507),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_635),
.A2(n_601),
.B(n_597),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_550),
.A2(n_508),
.B(n_514),
.C(n_367),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_563),
.B(n_507),
.Y(n_681)
);

NOR2x1_ASAP7_75t_L g682 ( 
.A(n_548),
.B(n_507),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_563),
.B(n_489),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_603),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_562),
.A2(n_393),
.B(n_367),
.C(n_382),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_555),
.B(n_489),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_635),
.A2(n_485),
.B(n_492),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_562),
.B(n_503),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_593),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_631),
.B(n_277),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_565),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_590),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_603),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_586),
.B(n_385),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_604),
.A2(n_487),
.B(n_306),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_561),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_559),
.B(n_424),
.C(n_434),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_572),
.B(n_385),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_551),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_605),
.A2(n_487),
.B(n_301),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_591),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_574),
.A2(n_390),
.B(n_389),
.C(n_391),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_610),
.B(n_395),
.Y(n_704)
);

OAI21xp33_ASAP7_75t_L g705 ( 
.A1(n_557),
.A2(n_328),
.B(n_355),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_559),
.A2(n_208),
.B(n_310),
.C(n_308),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_600),
.A2(n_487),
.B(n_278),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_602),
.A2(n_487),
.B(n_279),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_610),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_623),
.A2(n_487),
.B(n_98),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_606),
.A2(n_487),
.B(n_305),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_560),
.B(n_340),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_610),
.B(n_290),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_566),
.A2(n_292),
.B1(n_297),
.B2(n_300),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_567),
.A2(n_348),
.B1(n_342),
.B2(n_343),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_340),
.Y(n_716)
);

OA21x2_ASAP7_75t_L g717 ( 
.A1(n_583),
.A2(n_88),
.B(n_187),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_587),
.A2(n_348),
.B(n_345),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_608),
.A2(n_85),
.B(n_109),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_607),
.A2(n_612),
.B(n_545),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_613),
.A2(n_82),
.B(n_185),
.Y(n_721)
);

BUFx4f_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_619),
.A2(n_79),
.B(n_183),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_568),
.B(n_342),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_629),
.A2(n_77),
.B(n_177),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_585),
.B(n_434),
.Y(n_726)
);

BUFx4_ASAP7_75t_SL g727 ( 
.A(n_590),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_609),
.B(n_404),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_630),
.A2(n_345),
.B(n_343),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_625),
.B(n_415),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_632),
.A2(n_458),
.B(n_415),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_626),
.A2(n_59),
.B(n_176),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_595),
.A2(n_458),
.B(n_58),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_626),
.B(n_5),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_584),
.A2(n_53),
.B1(n_167),
.B2(n_165),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_638),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_553),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_710),
.A2(n_621),
.B(n_580),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_690),
.A2(n_552),
.B(n_558),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_552),
.B(n_558),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_669),
.B(n_617),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_646),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_689),
.B(n_584),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_698),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_660),
.B(n_638),
.Y(n_745)
);

CKINVDCx11_ASAP7_75t_R g746 ( 
.A(n_666),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_661),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_661),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_645),
.A2(n_579),
.B(n_594),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_688),
.A2(n_570),
.B1(n_628),
.B2(n_637),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_676),
.B(n_697),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_687),
.A2(n_594),
.B(n_636),
.Y(n_752)
);

OAI22x1_ASAP7_75t_L g753 ( 
.A1(n_715),
.A2(n_628),
.B1(n_598),
.B2(n_627),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_644),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_687),
.A2(n_732),
.B(n_647),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_642),
.A2(n_570),
.B(n_614),
.C(n_558),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_616),
.Y(n_757)
);

OAI21xp33_ASAP7_75t_L g758 ( 
.A1(n_712),
.A2(n_620),
.B(n_9),
.Y(n_758)
);

AO31x2_ASAP7_75t_L g759 ( 
.A1(n_642),
.A2(n_631),
.A3(n_620),
.B(n_558),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_675),
.A2(n_552),
.B(n_620),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_679),
.A2(n_656),
.B(n_655),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_645),
.A2(n_631),
.B(n_620),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_699),
.B(n_631),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_668),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_702),
.B(n_552),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_707),
.A2(n_708),
.B(n_681),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_680),
.A2(n_631),
.B(n_10),
.C(n_11),
.Y(n_767)
);

O2A1O1Ixp5_ASAP7_75t_L g768 ( 
.A1(n_672),
.A2(n_631),
.B(n_68),
.C(n_73),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_677),
.A2(n_52),
.B(n_164),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_724),
.B(n_8),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_662),
.A2(n_671),
.B(n_647),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_684),
.Y(n_772)
);

AOI21x1_ASAP7_75t_L g773 ( 
.A1(n_679),
.A2(n_62),
.B(n_160),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_643),
.A2(n_51),
.B(n_159),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_643),
.A2(n_657),
.B(n_659),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_653),
.A2(n_49),
.B(n_155),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_646),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_648),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_720),
.A2(n_48),
.B(n_154),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_658),
.B(n_172),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_696),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_674),
.A2(n_153),
.B(n_151),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_695),
.A2(n_147),
.B(n_146),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_700),
.A2(n_143),
.B(n_142),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_719),
.A2(n_141),
.B(n_139),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_722),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_654),
.A2(n_134),
.B(n_133),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_650),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_665),
.B(n_683),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_736),
.A2(n_10),
.A3(n_11),
.B(n_13),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_705),
.B(n_13),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_652),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_SL g793 ( 
.A(n_691),
.B(n_14),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_664),
.A2(n_670),
.B(n_663),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_673),
.B(n_14),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_709),
.B(n_15),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_722),
.B(n_129),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_709),
.B(n_15),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_692),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_651),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_713),
.A2(n_127),
.B(n_126),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_682),
.A2(n_122),
.B(n_118),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_778),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_743),
.A2(n_701),
.B1(n_716),
.B2(n_728),
.Y(n_804)
);

INVx3_ASAP7_75t_SL g805 ( 
.A(n_799),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_777),
.B(n_704),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_743),
.B(n_686),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_799),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_777),
.B(n_730),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_745),
.B(n_694),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_788),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_744),
.B(n_685),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_786),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_761),
.A2(n_735),
.B(n_706),
.C(n_733),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_754),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_741),
.B(n_714),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_766),
.A2(n_711),
.B(n_723),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_765),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_754),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_750),
.A2(n_703),
.B1(n_730),
.B2(n_731),
.Y(n_821)
);

NOR2x1_ASAP7_75t_SL g822 ( 
.A(n_742),
.B(n_734),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_739),
.A2(n_725),
.B(n_721),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_764),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_764),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_792),
.Y(n_826)
);

AOI222xp33_ASAP7_75t_L g827 ( 
.A1(n_791),
.A2(n_649),
.B1(n_718),
.B2(n_726),
.C1(n_667),
.C2(n_729),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_791),
.A2(n_770),
.B1(n_729),
.B2(n_797),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_SL g829 ( 
.A1(n_756),
.A2(n_733),
.B(n_693),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_772),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_772),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_760),
.A2(n_737),
.B(n_731),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_786),
.B(n_730),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_758),
.A2(n_727),
.B1(n_717),
.B2(n_667),
.C(n_20),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_717),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_781),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_741),
.B(n_16),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_747),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_740),
.A2(n_794),
.B(n_756),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_787),
.A2(n_115),
.B(n_113),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_789),
.B(n_16),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_796),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_775),
.A2(n_112),
.B(n_111),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_751),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_795),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_757),
.B(n_22),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_747),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_753),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_742),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_767),
.B(n_23),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_767),
.B(n_24),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_780),
.A2(n_798),
.B(n_768),
.C(n_797),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_748),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_780),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_793),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_748),
.Y(n_856)
);

BUFx6f_ASAP7_75t_SL g857 ( 
.A(n_742),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_836),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_816),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_821),
.A2(n_765),
.B1(n_763),
.B2(n_800),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_820),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_824),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_830),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_828),
.A2(n_765),
.B1(n_782),
.B2(n_769),
.Y(n_864)
);

BUFx4f_ASAP7_75t_SL g865 ( 
.A(n_805),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_835),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_814),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_838),
.Y(n_868)
);

CKINVDCx11_ASAP7_75t_R g869 ( 
.A(n_805),
.Y(n_869)
);

BUFx2_ASAP7_75t_SL g870 ( 
.A(n_857),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_825),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_813),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_814),
.Y(n_875)
);

CKINVDCx11_ASAP7_75t_R g876 ( 
.A(n_826),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_819),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_829),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_823),
.A2(n_738),
.B(n_755),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_847),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_832),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_839),
.A2(n_818),
.B(n_773),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_847),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_810),
.A2(n_801),
.B1(n_779),
.B2(n_774),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_808),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_838),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_806),
.B(n_775),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_849),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_856),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_856),
.Y(n_892)
);

INVx6_ASAP7_75t_L g893 ( 
.A(n_814),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_812),
.Y(n_894)
);

OAI22xp33_ASAP7_75t_L g895 ( 
.A1(n_804),
.A2(n_784),
.B1(n_790),
.B2(n_746),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_828),
.A2(n_746),
.B1(n_776),
.B2(n_752),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_842),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_853),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_819),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_850),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_822),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_827),
.A2(n_752),
.B1(n_802),
.B2(n_783),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_852),
.A2(n_755),
.B(n_771),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_810),
.A2(n_749),
.B1(n_785),
.B2(n_762),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_848),
.B(n_845),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_848),
.A2(n_785),
.B1(n_738),
.B2(n_790),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_845),
.B(n_790),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_806),
.B(n_759),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_851),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_834),
.A2(n_790),
.B1(n_768),
.B2(n_759),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_807),
.B(n_759),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_815),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_809),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_815),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_846),
.B(n_759),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_866),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_889),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_911),
.B(n_846),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_881),
.A2(n_843),
.B(n_840),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_889),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_889),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_905),
.A2(n_844),
.B1(n_841),
.B2(n_855),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_880),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_911),
.B(n_837),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_915),
.B(n_817),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_895),
.A2(n_854),
.B(n_855),
.Y(n_930)
);

AOI21x1_ASAP7_75t_L g931 ( 
.A1(n_884),
.A2(n_809),
.B(n_833),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_866),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_866),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_881),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_912),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_908),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_868),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_912),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_908),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_907),
.B(n_809),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_872),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_884),
.A2(n_833),
.B(n_857),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_872),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_882),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_872),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_914),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_915),
.B(n_908),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_882),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_880),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_888),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_888),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_903),
.B(n_814),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_919),
.B(n_900),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_948),
.B(n_908),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_944),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_918),
.B(n_903),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_948),
.B(n_882),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_924),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_951),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_900),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_925),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_940),
.B(n_929),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_925),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_951),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_948),
.B(n_892),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_925),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_922),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_940),
.B(n_894),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_925),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_951),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_952),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_940),
.B(n_892),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_952),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_933),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_944),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_949),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_922),
.B(n_918),
.Y(n_979)
);

INVx4_ASAP7_75t_R g980 ( 
.A(n_928),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_929),
.B(n_892),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_952),
.Y(n_982)
);

NAND2x1_ASAP7_75t_L g983 ( 
.A(n_922),
.B(n_901),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_941),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_933),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_941),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_933),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_937),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_943),
.Y(n_989)
);

OAI221xp5_ASAP7_75t_L g990 ( 
.A1(n_970),
.A2(n_923),
.B1(n_860),
.B2(n_909),
.C(n_887),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_958),
.B(n_936),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_958),
.B(n_936),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_SL g993 ( 
.A1(n_970),
.A2(n_923),
.B(n_905),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_966),
.B(n_936),
.Y(n_994)
);

AOI221xp5_ASAP7_75t_L g995 ( 
.A1(n_954),
.A2(n_919),
.B1(n_897),
.B2(n_929),
.C(n_928),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_955),
.B(n_936),
.Y(n_996)
);

AOI221xp5_ASAP7_75t_L g997 ( 
.A1(n_954),
.A2(n_897),
.B1(n_928),
.B2(n_930),
.C(n_909),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_966),
.B(n_955),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_961),
.B(n_949),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_961),
.B(n_950),
.Y(n_1000)
);

AOI211xp5_ASAP7_75t_SL g1001 ( 
.A1(n_988),
.A2(n_922),
.B(n_939),
.C(n_936),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_963),
.B(n_950),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_963),
.B(n_950),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_981),
.B(n_950),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_981),
.B(n_916),
.Y(n_1005)
);

AOI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_988),
.A2(n_930),
.B1(n_858),
.B2(n_879),
.C(n_896),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_974),
.B(n_930),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_974),
.B(n_916),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_977),
.B(n_932),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_957),
.B(n_860),
.C(n_886),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_977),
.B(n_932),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_979),
.B(n_939),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_956),
.B(n_926),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_957),
.B(n_902),
.C(n_927),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_998),
.B(n_979),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_1013),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_1007),
.B(n_869),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_998),
.B(n_979),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1002),
.B(n_956),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_1012),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1003),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1007),
.B(n_978),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_991),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1008),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1009),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_999),
.B(n_978),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_991),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_992),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_992),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_1005),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_993),
.B(n_927),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_994),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_994),
.Y(n_1033)
);

NAND2x1_ASAP7_75t_L g1034 ( 
.A(n_1012),
.B(n_980),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1004),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1020),
.B(n_996),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1020),
.B(n_1001),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1034),
.B(n_979),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_1034),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1015),
.B(n_957),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1019),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1022),
.B(n_1000),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1019),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1026),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1024),
.B(n_995),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1015),
.B(n_957),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1023),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1044),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_1045),
.B(n_865),
.Y(n_1049)
);

BUFx2_ASAP7_75t_SL g1050 ( 
.A(n_1039),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_L g1051 ( 
.A(n_1039),
.B(n_1017),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1044),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1037),
.B(n_1018),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1047),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_1048),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_1051),
.B(n_1006),
.C(n_1010),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1051),
.A2(n_1049),
.B1(n_1014),
.B2(n_1053),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_876),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_1058),
.B(n_1050),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1057),
.A2(n_1052),
.B1(n_1050),
.B2(n_1041),
.C(n_1043),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_1055),
.B(n_990),
.C(n_1054),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1056),
.B(n_997),
.C(n_1054),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1055),
.B(n_1041),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1058),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1055),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_1055),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1055),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1066),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1065),
.B(n_1043),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1067),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_1060),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1059),
.B(n_1037),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1069),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1068),
.B(n_1047),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1064),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1062),
.B(n_1047),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1063),
.B(n_870),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_L g1080 ( 
.A(n_1064),
.B(n_1038),
.Y(n_1080)
);

OAI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1061),
.A2(n_1031),
.B1(n_1042),
.B2(n_1038),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1059),
.B(n_1040),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1068),
.B(n_1042),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1066),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1068),
.B(n_1040),
.Y(n_1085)
);

AOI211x1_ASAP7_75t_L g1086 ( 
.A1(n_1081),
.A2(n_1046),
.B(n_1025),
.C(n_1024),
.Y(n_1086)
);

AOI211xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1070),
.A2(n_890),
.B(n_1038),
.C(n_870),
.Y(n_1087)
);

NOR4xp25_ASAP7_75t_L g1088 ( 
.A(n_1073),
.B(n_1025),
.C(n_1030),
.D(n_1046),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_1078),
.A2(n_1038),
.B(n_1036),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1077),
.B(n_1036),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1079),
.A2(n_930),
.B(n_1016),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_R g1092 ( 
.A(n_1072),
.B(n_26),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1075),
.B(n_1021),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1084),
.B(n_874),
.C(n_871),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1078),
.A2(n_930),
.B(n_874),
.C(n_871),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1071),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1074),
.B(n_1021),
.Y(n_1097)
);

OAI221xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1083),
.A2(n_1085),
.B1(n_1076),
.B2(n_1082),
.C(n_1080),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1083),
.A2(n_1026),
.B(n_874),
.C(n_871),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1073),
.A2(n_1035),
.B(n_913),
.C(n_983),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1073),
.B(n_1018),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_1079),
.Y(n_1102)
);

OAI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1073),
.A2(n_957),
.B1(n_983),
.B2(n_1035),
.C1(n_953),
.C2(n_1028),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_1081),
.A2(n_931),
.B(n_942),
.C(n_1011),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1090),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1098),
.B(n_1023),
.Y(n_1106)
);

NOR3x1_ASAP7_75t_L g1107 ( 
.A(n_1096),
.B(n_879),
.C(n_921),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1092),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1094),
.B(n_27),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_1102),
.B(n_28),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1086),
.B(n_28),
.C(n_29),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1097),
.B(n_1027),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1093),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1091),
.A2(n_901),
.B(n_864),
.Y(n_1114)
);

NAND4xp25_ASAP7_75t_L g1115 ( 
.A(n_1087),
.B(n_910),
.C(n_901),
.D(n_906),
.Y(n_1115)
);

NOR3x1_ASAP7_75t_L g1116 ( 
.A(n_1101),
.B(n_918),
.C(n_921),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_1089),
.B(n_867),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1100),
.B(n_1027),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1088),
.B(n_1028),
.Y(n_1119)
);

NOR4xp25_ASAP7_75t_L g1120 ( 
.A(n_1095),
.B(n_30),
.C(n_32),
.D(n_33),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1104),
.B(n_1029),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_1099),
.B1(n_1103),
.B2(n_1089),
.C(n_1033),
.Y(n_1122)
);

OAI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1108),
.A2(n_1033),
.B1(n_1032),
.B2(n_1029),
.C(n_957),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1105),
.B(n_1032),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1110),
.B(n_30),
.Y(n_1125)
);

NOR4xp25_ASAP7_75t_L g1126 ( 
.A(n_1113),
.B(n_32),
.C(n_34),
.D(n_35),
.Y(n_1126)
);

OR3x1_ASAP7_75t_L g1127 ( 
.A(n_1106),
.B(n_34),
.C(n_36),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1109),
.B(n_36),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_SL g1129 ( 
.A1(n_1111),
.A2(n_37),
.B(n_38),
.Y(n_1129)
);

NAND4xp25_ASAP7_75t_SL g1130 ( 
.A(n_1111),
.B(n_37),
.C(n_39),
.D(n_40),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_L g1131 ( 
.A(n_1119),
.B(n_39),
.C(n_42),
.D(n_45),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1112),
.B(n_42),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_L g1133 ( 
.A(n_1118),
.B(n_931),
.C(n_867),
.Y(n_1133)
);

NOR3x1_ASAP7_75t_L g1134 ( 
.A(n_1121),
.B(n_921),
.C(n_937),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1107),
.B(n_1116),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_1114),
.B(n_1115),
.Y(n_1136)
);

AOI211xp5_ASAP7_75t_L g1137 ( 
.A1(n_1117),
.A2(n_875),
.B(n_873),
.C(n_885),
.Y(n_1137)
);

NAND4xp75_ASAP7_75t_L g1138 ( 
.A(n_1110),
.B(n_891),
.C(n_873),
.D(n_861),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_SL g1139 ( 
.A(n_1108),
.B(n_867),
.C(n_878),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_SL g1140 ( 
.A(n_1106),
.B(n_861),
.C(n_863),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_SL g1141 ( 
.A(n_1106),
.B(n_859),
.C(n_863),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_L g1142 ( 
.A(n_1108),
.B(n_867),
.C(n_942),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1117),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_L g1144 ( 
.A(n_1110),
.B(n_875),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1108),
.B(n_87),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1129),
.B(n_989),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1145),
.B(n_1126),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1130),
.A2(n_893),
.B1(n_922),
.B2(n_891),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1131),
.A2(n_878),
.B(n_953),
.C(n_898),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1131),
.B(n_893),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1125),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1127),
.A2(n_893),
.B1(n_953),
.B2(n_969),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1144),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1128),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1138),
.Y(n_1155)
);

OAI211xp5_ASAP7_75t_L g1156 ( 
.A1(n_1143),
.A2(n_875),
.B(n_878),
.C(n_904),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1132),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1139),
.B(n_875),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1124),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_1136),
.B(n_899),
.C(n_877),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1140),
.B(n_989),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1135),
.B(n_893),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1141),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1134),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1123),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1142),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_1137),
.B(n_92),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1133),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1122),
.A2(n_893),
.B1(n_953),
.B2(n_969),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1169),
.A2(n_953),
.B1(n_969),
.B2(n_984),
.Y(n_1170)
);

OAI21xp33_ASAP7_75t_L g1171 ( 
.A1(n_1162),
.A2(n_953),
.B(n_969),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1147),
.B(n_904),
.C(n_898),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1153),
.A2(n_898),
.B(n_862),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_L g1174 ( 
.A(n_1154),
.B(n_1151),
.Y(n_1174)
);

NAND4xp25_ASAP7_75t_L g1175 ( 
.A(n_1165),
.B(n_859),
.C(n_862),
.D(n_877),
.Y(n_1175)
);

NAND4xp75_ASAP7_75t_L g1176 ( 
.A(n_1157),
.B(n_984),
.C(n_986),
.D(n_982),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1159),
.B(n_986),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1150),
.Y(n_1178)
);

AOI211xp5_ASAP7_75t_L g1179 ( 
.A1(n_1155),
.A2(n_875),
.B(n_927),
.C(n_982),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1163),
.Y(n_1180)
);

OR5x1_ASAP7_75t_L g1181 ( 
.A(n_1156),
.B(n_980),
.C(n_875),
.D(n_953),
.E(n_103),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1166),
.B(n_899),
.C(n_877),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1168),
.B(n_973),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1152),
.A2(n_927),
.B1(n_973),
.B2(n_975),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1164),
.B(n_93),
.Y(n_1185)
);

NOR4xp75_ASAP7_75t_SL g1186 ( 
.A(n_1146),
.B(n_97),
.C(n_100),
.D(n_110),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1148),
.B(n_877),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1158),
.A2(n_1161),
.B1(n_1167),
.B2(n_1160),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1167),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1149),
.A2(n_927),
.B1(n_899),
.B2(n_975),
.C(n_960),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1153),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1180),
.B(n_972),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1174),
.B(n_899),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1189),
.A2(n_920),
.B(n_943),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1191),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1178),
.B(n_927),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_L g1197 ( 
.A(n_1185),
.B(n_927),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1173),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1182),
.B(n_939),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1183),
.B(n_972),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1188),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_L g1202 ( 
.A(n_1175),
.B(n_946),
.C(n_926),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1183),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1177),
.B(n_967),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1173),
.Y(n_1205)
);

XNOR2xp5_ASAP7_75t_L g1206 ( 
.A(n_1181),
.B(n_926),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1195),
.B(n_1187),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1203),
.A2(n_1172),
.B1(n_1184),
.B2(n_1186),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1193),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1201),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_1198),
.B(n_1170),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1205),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1193),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1206),
.A2(n_1179),
.B1(n_1171),
.B2(n_1190),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1197),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1206),
.A2(n_1176),
.B1(n_927),
.B2(n_917),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1192),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1196),
.B(n_917),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1200),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1199),
.Y(n_1220)
);

XNOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1204),
.B(n_939),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1209),
.A2(n_1202),
.B(n_1194),
.C(n_935),
.Y(n_1222)
);

NOR4xp25_ASAP7_75t_L g1223 ( 
.A(n_1212),
.B(n_960),
.C(n_965),
.D(n_967),
.Y(n_1223)
);

OR3x1_ASAP7_75t_L g1224 ( 
.A(n_1217),
.B(n_965),
.C(n_946),
.Y(n_1224)
);

XNOR2x2_ASAP7_75t_SL g1225 ( 
.A(n_1213),
.B(n_920),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1210),
.B(n_947),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1207),
.B(n_947),
.C(n_945),
.Y(n_1227)
);

OAI222xp33_ASAP7_75t_L g1228 ( 
.A1(n_1214),
.A2(n_947),
.B1(n_935),
.B2(n_938),
.C1(n_945),
.C2(n_939),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1216),
.A2(n_945),
.B1(n_947),
.B2(n_935),
.C(n_938),
.Y(n_1229)
);

AOI222xp33_ASAP7_75t_L g1230 ( 
.A1(n_1211),
.A2(n_959),
.B1(n_971),
.B2(n_968),
.C1(n_964),
.C2(n_962),
.Y(n_1230)
);

NOR2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1220),
.B(n_935),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1226),
.A2(n_1215),
.B(n_1219),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1231),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1230),
.A2(n_1221),
.B(n_1208),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1224),
.A2(n_1208),
.B1(n_1218),
.B2(n_938),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1222),
.Y(n_1236)
);

OAI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1225),
.A2(n_987),
.B1(n_985),
.B2(n_976),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1233),
.B(n_1229),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1232),
.A2(n_1228),
.B(n_1227),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1234),
.A2(n_1223),
.B(n_920),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1236),
.A2(n_945),
.B(n_938),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1238),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1242),
.B(n_1239),
.Y(n_1243)
);

AOI222xp33_ASAP7_75t_L g1244 ( 
.A1(n_1243),
.A2(n_1235),
.B1(n_1237),
.B2(n_1241),
.C1(n_1240),
.C2(n_934),
.Y(n_1244)
);

OAI221xp5_ASAP7_75t_R g1245 ( 
.A1(n_1244),
.A2(n_920),
.B1(n_987),
.B2(n_985),
.C(n_976),
.Y(n_1245)
);

AOI211xp5_ASAP7_75t_L g1246 ( 
.A1(n_1245),
.A2(n_987),
.B(n_985),
.C(n_976),
.Y(n_1246)
);


endmodule