module fake_jpeg_3336_n_452 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_25),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_58),
.B(n_74),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_89),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_83),
.Y(n_125)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_79),
.B(n_115),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_10),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_94),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_32),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_9),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_99),
.B(n_102),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_11),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_46),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_27),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_104),
.B(n_107),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_106),
.A2(n_50),
.B(n_3),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_21),
.B(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_26),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_26),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_30),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_114),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_30),
.B(n_7),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_52),
.B1(n_24),
.B2(n_23),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_117),
.A2(n_122),
.B1(n_129),
.B2(n_131),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_91),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_121),
.A2(n_139),
.B1(n_151),
.B2(n_159),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_58),
.B1(n_74),
.B2(n_69),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_84),
.B(n_23),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_52),
.B1(n_24),
.B2(n_43),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_54),
.B1(n_43),
.B2(n_22),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_134),
.A2(n_170),
.B1(n_129),
.B2(n_158),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_146),
.B1(n_158),
.B2(n_81),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_86),
.A2(n_54),
.B1(n_19),
.B2(n_22),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_79),
.A2(n_39),
.B1(n_31),
.B2(n_28),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_19),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_150),
.B(n_164),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_50),
.B1(n_12),
.B2(n_14),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_67),
.A2(n_72),
.B(n_115),
.Y(n_155)
);

BUFx12f_ASAP7_75t_SL g201 ( 
.A(n_155),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_88),
.A2(n_50),
.B1(n_3),
.B2(n_5),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_63),
.B(n_14),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_50),
.B1(n_14),
.B2(n_16),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_186),
.B1(n_139),
.B2(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_71),
.B(n_2),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_172),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_60),
.A2(n_50),
.B1(n_3),
.B2(n_5),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_71),
.B(n_2),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_85),
.B(n_87),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_65),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_146),
.B(n_182),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_193),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_189),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_73),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_212),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_192),
.A2(n_208),
.B(n_216),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_105),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_182),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g251 ( 
.A(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_203),
.Y(n_254)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_152),
.Y(n_197)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_205),
.B1(n_215),
.B2(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_105),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_134),
.A2(n_64),
.B1(n_131),
.B2(n_117),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_64),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_218),
.Y(n_268)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_210),
.B(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_126),
.B(n_133),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_145),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_122),
.B(n_135),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_227),
.B(n_230),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_143),
.A2(n_171),
.B1(n_156),
.B2(n_137),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_125),
.B(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_223),
.Y(n_275)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_141),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_116),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_118),
.B(n_127),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_240),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_148),
.B(n_142),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_118),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_229),
.A2(n_242),
.B1(n_207),
.B2(n_215),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_154),
.A2(n_147),
.B(n_161),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_132),
.B(n_128),
.C(n_130),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_132),
.A2(n_169),
.B1(n_183),
.B2(n_161),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_234),
.A2(n_236),
.B1(n_194),
.B2(n_204),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_157),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_183),
.B1(n_185),
.B2(n_157),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_173),
.A2(n_134),
.B1(n_129),
.B2(n_119),
.Y(n_237)
);

AO22x1_ASAP7_75t_L g238 ( 
.A1(n_173),
.A2(n_182),
.B1(n_181),
.B2(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_241),
.Y(n_261)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_124),
.B(n_181),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_144),
.A2(n_187),
.B(n_182),
.C(n_140),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_151),
.A2(n_165),
.B1(n_159),
.B2(n_139),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_120),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_248),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_152),
.Y(n_245)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_124),
.B(n_181),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_200),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_256),
.B(n_257),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_270),
.B(n_278),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_197),
.B1(n_245),
.B2(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_247),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_287),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_242),
.A2(n_207),
.B1(n_208),
.B2(n_201),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_214),
.B1(n_246),
.B2(n_189),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_228),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_286),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_212),
.B(n_238),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_204),
.A2(n_191),
.B(n_201),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_196),
.B(n_199),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_226),
.B(n_232),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_202),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_213),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_304),
.B(n_306),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_216),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_300),
.B(n_321),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_263),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_303),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_255),
.A2(n_206),
.B(n_241),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_271),
.A2(n_230),
.B1(n_239),
.B2(n_198),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_310),
.B1(n_313),
.B2(n_319),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_233),
.A3(n_221),
.B1(n_209),
.B2(n_197),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_285),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_231),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_315),
.B(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_318),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_245),
.B1(n_248),
.B2(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_281),
.B1(n_250),
.B2(n_255),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_316),
.B1(n_251),
.B2(n_291),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_276),
.A2(n_261),
.B(n_273),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_266),
.B1(n_289),
.B2(n_260),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_261),
.B(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_266),
.A2(n_250),
.B1(n_257),
.B2(n_260),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_268),
.A2(n_276),
.B1(n_251),
.B2(n_277),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_291),
.B1(n_283),
.B2(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_263),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_249),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_325),
.Y(n_332)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_324),
.B(n_328),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_262),
.B(n_265),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_265),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_329),
.Y(n_348)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_252),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_330),
.B(n_309),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_339),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_251),
.C(n_259),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_349),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_341),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_322),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_283),
.B1(n_293),
.B2(n_294),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_344),
.A2(n_350),
.B1(n_355),
.B2(n_329),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_267),
.C(n_253),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_314),
.A2(n_267),
.B1(n_279),
.B2(n_253),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_258),
.B(n_264),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_351),
.A2(n_354),
.B(n_306),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_258),
.C(n_264),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_357),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_326),
.A2(n_274),
.B(n_252),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_279),
.B1(n_274),
.B2(n_285),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_320),
.B1(n_302),
.B2(n_299),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_296),
.B(n_317),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_346),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_371),
.Y(n_388)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_307),
.B1(n_297),
.B2(n_323),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_367),
.B1(n_372),
.B2(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_325),
.Y(n_369)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_313),
.B(n_305),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_296),
.B1(n_304),
.B2(n_307),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_379),
.Y(n_392)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_302),
.B1(n_303),
.B2(n_321),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_380),
.A2(n_336),
.B1(n_344),
.B2(n_358),
.Y(n_397)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_336),
.B1(n_356),
.B2(n_350),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_384),
.A2(n_387),
.B1(n_397),
.B2(n_359),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_337),
.C(n_357),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_331),
.C(n_349),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_360),
.A2(n_341),
.B1(n_380),
.B2(n_361),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_332),
.C(n_331),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_370),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_360),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_395),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_369),
.Y(n_402)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_378),
.B1(n_361),
.B2(n_375),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_410),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_398),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_408),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_370),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_407),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_353),
.Y(n_406)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_372),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_390),
.C(n_338),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_332),
.B1(n_377),
.B2(n_362),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_411),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_412),
.B(n_382),
.Y(n_414)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_416),
.B(n_409),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_403),
.A2(n_388),
.B1(n_396),
.B2(n_393),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_422),
.B1(n_383),
.B2(n_381),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_400),
.A2(n_396),
.B1(n_393),
.B2(n_385),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_428),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_419),
.A2(n_394),
.B(n_368),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_426),
.B(n_432),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_423),
.A2(n_400),
.B(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_427),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_353),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_431),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_399),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_345),
.B(n_381),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_426),
.A2(n_416),
.B(n_418),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_435),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_429),
.B(n_413),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_417),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_427),
.A2(n_414),
.B(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_439),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_405),
.C(n_415),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_441),
.Y(n_447)
);

XOR2x2_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_432),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_414),
.B(n_385),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_434),
.C(n_433),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.C(n_440),
.Y(n_449)
);

O2A1O1Ixp33_ASAP7_75t_SL g448 ( 
.A1(n_447),
.A2(n_444),
.B(n_442),
.C(n_383),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_449),
.C(n_399),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_450),
.B(n_342),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_364),
.Y(n_452)
);


endmodule