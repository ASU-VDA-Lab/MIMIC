module fake_jpeg_23541_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_15),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_17),
.B1(n_14),
.B2(n_25),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.C(n_38),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_10),
.C(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_13),
.B1(n_12),
.B2(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_16),
.B1(n_23),
.B2(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_15),
.A3(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_44),
.B1(n_42),
.B2(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_46),
.B1(n_57),
.B2(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_22),
.C(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_64),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_67),
.B2(n_4),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_73),
.B1(n_5),
.B2(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_3),
.Y(n_76)
);


endmodule