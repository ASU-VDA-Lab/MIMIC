module fake_ibex_751_n_1129 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1129);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1129;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_947;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_412;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_449;
wire n_547;
wire n_727;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_671;
wire n_228;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_591;
wire n_453;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_325;
wire n_496;
wire n_301;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_943;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1082;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_1028;
wire n_1012;
wire n_993;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_721;
wire n_365;
wire n_581;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_1057;
wire n_1049;
wire n_1086;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_921;
wire n_874;
wire n_890;
wire n_1058;
wire n_1105;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_984;
wire n_1000;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_178),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_127),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_117),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_64),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_145),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_122),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_105),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_72),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_188),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_14),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_135),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_67),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_93),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_89),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_108),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_37),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_174),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_58),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_119),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_109),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_90),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_47),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_39),
.B(n_170),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_31),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_184),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_10),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_87),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_204),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_111),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_121),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_141),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_25),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_107),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_216),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_47),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_182),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_125),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_26),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_192),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_196),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_29),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_106),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_60),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_183),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_74),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_186),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_16),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_98),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_65),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_68),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_153),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_202),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_142),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_114),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_7),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_214),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_76),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_92),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_88),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_101),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_133),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_95),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_129),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_62),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_71),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_57),
.B(n_172),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_137),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_11),
.Y(n_321)
);

INVx4_ASAP7_75t_R g322 ( 
.A(n_166),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_63),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_49),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_171),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_118),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_51),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_97),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_61),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_45),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_143),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_29),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_66),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_116),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_99),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_86),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_211),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_134),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_9),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_165),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_160),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_30),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_45),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_181),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_53),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_4),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_158),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_17),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_50),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_206),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_51),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_124),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_149),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_96),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_163),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_85),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_189),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_150),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_167),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_123),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_36),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_146),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_81),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_130),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_173),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_79),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_94),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_91),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_194),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_217),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_2),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_83),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_112),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_198),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_50),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_10),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_103),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_191),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_46),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_23),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_295),
.B(n_59),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_280),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_378),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_290),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g391 ( 
.A1(n_236),
.A2(n_77),
.B(n_220),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_267),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_270),
.B(n_1),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_295),
.B(n_1),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_267),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_280),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_236),
.A2(n_78),
.B(n_215),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_254),
.A2(n_75),
.B(n_213),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_280),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_289),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_2),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_254),
.A2(n_73),
.B(n_209),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_280),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_297),
.B(n_3),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_289),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_378),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_278),
.A2(n_308),
.B(n_302),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_297),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_5),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_366),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_245),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_270),
.B(n_6),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_335),
.B(n_7),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_227),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_278),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_302),
.A2(n_80),
.B(n_205),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_229),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_258),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_288),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_258),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_353),
.B(n_8),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_355),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_226),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_240),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_240),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_434)
);

OA21x2_ASAP7_75t_L g435 ( 
.A1(n_308),
.A2(n_82),
.B(n_203),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_232),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_242),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_243),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_315),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_246),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_225),
.B(n_13),
.Y(n_441)
);

BUFx12f_ASAP7_75t_L g442 ( 
.A(n_231),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_304),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_279),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_315),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_307),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_279),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_251),
.B(n_13),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_247),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_252),
.B(n_253),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_317),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_317),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_256),
.A2(n_84),
.B(n_201),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_341),
.B(n_354),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_259),
.B(n_15),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_260),
.B(n_15),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_261),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_271),
.A2(n_273),
.B(n_272),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_223),
.B(n_16),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_376),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_327),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_226),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_226),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_276),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_283),
.B(n_18),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_327),
.Y(n_468)
);

BUFx8_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_309),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_389),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_402),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_459),
.B(n_298),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_446),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_326),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

CKINVDCx6p67_ASAP7_75t_R g482 ( 
.A(n_442),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_428),
.B(n_347),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_349),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_431),
.B(n_379),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_405),
.B(n_226),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_428),
.B(n_331),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_394),
.B(n_352),
.C(n_264),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_423),
.B(n_306),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_352),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_262),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_402),
.B(n_417),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_233),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_409),
.B(n_275),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_383),
.B1(n_382),
.B2(n_282),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_233),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_234),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_423),
.B(n_310),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_426),
.B(n_311),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_414),
.B(n_312),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_426),
.B(n_314),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_387),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_442),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_436),
.B(n_368),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_433),
.Y(n_519)
);

AO22x2_ASAP7_75t_L g520 ( 
.A1(n_448),
.A2(n_344),
.B1(n_374),
.B2(n_299),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_436),
.B(n_316),
.Y(n_522)
);

BUFx4f_ASAP7_75t_L g523 ( 
.A(n_430),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_466),
.A2(n_340),
.B1(n_286),
.B2(n_321),
.Y(n_524)
);

NOR3xp33_ASAP7_75t_L g525 ( 
.A(n_409),
.B(n_330),
.C(n_324),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_387),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_418),
.B(n_346),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_437),
.B(n_319),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_320),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_468),
.A2(n_284),
.B1(n_235),
.B2(n_237),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_379),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_469),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_469),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_388),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_447),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

INVx4_ASAP7_75t_SL g540 ( 
.A(n_429),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_438),
.B(n_323),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_440),
.B(n_239),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_469),
.B(n_235),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_385),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_440),
.B(n_241),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

BUFx6f_ASAP7_75t_SL g547 ( 
.A(n_449),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_449),
.B(n_325),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_450),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_429),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_448),
.A2(n_300),
.B1(n_237),
.B2(n_303),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_401),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_385),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_466),
.B(n_386),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_392),
.B(n_328),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_386),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_386),
.B(n_244),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_410),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_392),
.B(n_395),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_460),
.B(n_350),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_469),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_410),
.A2(n_287),
.B1(n_337),
.B2(n_377),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_451),
.B(n_329),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_400),
.B(n_248),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_434),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g570 ( 
.A(n_441),
.B(n_284),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_439),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_441),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_422),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_400),
.B(n_406),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_439),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_406),
.B(n_334),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_407),
.B(n_248),
.Y(n_578)
);

AND3x1_ASAP7_75t_L g579 ( 
.A(n_434),
.B(n_263),
.C(n_336),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_407),
.B(n_342),
.Y(n_580)
);

OAI22x1_ASAP7_75t_L g581 ( 
.A1(n_463),
.A2(n_230),
.B1(n_285),
.B2(n_265),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_461),
.B(n_348),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_412),
.B(n_249),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_455),
.B(n_269),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_445),
.A2(n_356),
.B1(n_351),
.B2(n_360),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_391),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_398),
.A2(n_370),
.B(n_362),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_461),
.B(n_359),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_460),
.B(n_318),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_462),
.B(n_364),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_444),
.B(n_250),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_444),
.B(n_250),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_444),
.B(n_369),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_393),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_467),
.C(n_456),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_569),
.A2(n_463),
.B1(n_300),
.B2(n_292),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_535),
.B(n_536),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_421),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_560),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_479),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_572),
.B(n_277),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_553),
.A2(n_303),
.B1(n_292),
.B2(n_384),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_492),
.B(n_277),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_545),
.B(n_281),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_565),
.B(n_281),
.Y(n_612)
);

NAND2x1_ASAP7_75t_L g613 ( 
.A(n_508),
.B(n_322),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_485),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_508),
.A2(n_397),
.B1(n_391),
.B2(n_425),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_542),
.B(n_313),
.Y(n_618)
);

BUFx6f_ASAP7_75t_SL g619 ( 
.A(n_500),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_483),
.B(n_313),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_484),
.B(n_333),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_493),
.A2(n_338),
.B1(n_357),
.B2(n_361),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_338),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_517),
.B(n_398),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_480),
.B(n_357),
.Y(n_626)
);

AND2x4_ASAP7_75t_SL g627 ( 
.A(n_482),
.B(n_371),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_515),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_488),
.B(n_361),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_552),
.B(n_222),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_486),
.B(n_452),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_552),
.B(n_228),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_534),
.B(n_452),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_487),
.B(n_255),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_488),
.B(n_257),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_504),
.A2(n_425),
.B1(n_435),
.B2(n_373),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_487),
.B(n_266),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_584),
.B(n_268),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_554),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_521),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_547),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_493),
.A2(n_367),
.B1(n_358),
.B2(n_274),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_510),
.A2(n_548),
.B(n_529),
.C(n_471),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_537),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_481),
.B(n_523),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_493),
.A2(n_296),
.B1(n_305),
.B2(n_365),
.Y(n_650)
);

AND2x6_ASAP7_75t_SL g651 ( 
.A(n_497),
.B(n_20),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_496),
.B(n_291),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_562),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_499),
.B(n_375),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_503),
.B(n_380),
.Y(n_655)
);

INVxp33_ASAP7_75t_L g656 ( 
.A(n_530),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_523),
.B(n_224),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_531),
.A2(n_435),
.B1(n_403),
.B2(n_453),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_474),
.A2(n_453),
.B1(n_464),
.B2(n_432),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_598),
.B(n_238),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_474),
.A2(n_453),
.B1(n_464),
.B2(n_432),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_554),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_518),
.B(n_294),
.Y(n_663)
);

NOR2x2_ASAP7_75t_L g664 ( 
.A(n_497),
.B(n_21),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_571),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_518),
.B(n_301),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_568),
.B(n_381),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_432),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_489),
.B(n_432),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_563),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_527),
.B(n_464),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_566),
.B(n_387),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_578),
.B(n_404),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_583),
.B(n_404),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_495),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_549),
.B(n_404),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_527),
.B(n_477),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_SL g680 ( 
.A(n_566),
.B(n_408),
.C(n_411),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_551),
.B(n_22),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_571),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_491),
.B(n_408),
.Y(n_683)
);

OAI221xp5_ASAP7_75t_L g684 ( 
.A1(n_498),
.A2(n_420),
.B1(n_415),
.B2(n_411),
.C(n_465),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_576),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_491),
.B(n_411),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_494),
.B(n_465),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_576),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_505),
.B(n_387),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_520),
.B(n_22),
.Y(n_690)
);

AND2x6_ASAP7_75t_SL g691 ( 
.A(n_497),
.B(n_24),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_501),
.B(n_415),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_502),
.B(n_396),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_494),
.B(n_396),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_490),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_529),
.B(n_396),
.Y(n_697)
);

AND2x6_ASAP7_75t_SL g698 ( 
.A(n_537),
.B(n_28),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_558),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_593),
.A2(n_399),
.B(n_30),
.C(n_31),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_564),
.B(n_490),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_475),
.B(n_506),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_561),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_399),
.Y(n_704)
);

AND2x6_ASAP7_75t_SL g705 ( 
.A(n_592),
.B(n_28),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_525),
.B(n_32),
.C(n_33),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_500),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_475),
.B(n_32),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_506),
.B(n_33),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_533),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_520),
.B(n_34),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_507),
.B(n_34),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_507),
.B(n_35),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_562),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_538),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_520),
.B(n_36),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_509),
.B(n_37),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_38),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_587),
.B(n_126),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_38),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_522),
.B(n_39),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_522),
.B(n_128),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_607),
.B(n_543),
.Y(n_723)
);

O2A1O1Ixp5_ASAP7_75t_SL g724 ( 
.A1(n_689),
.A2(n_567),
.B(n_589),
.C(n_478),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_642),
.Y(n_725)
);

INVx3_ASAP7_75t_SL g726 ( 
.A(n_707),
.Y(n_726)
);

OAI22x1_ASAP7_75t_L g727 ( 
.A1(n_720),
.A2(n_570),
.B1(n_569),
.B2(n_579),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_604),
.A2(n_614),
.B1(n_701),
.B2(n_690),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_647),
.A2(n_605),
.B(n_681),
.C(n_671),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_604),
.A2(n_593),
.B(n_586),
.C(n_577),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_574),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_616),
.B(n_498),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_608),
.B(n_677),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_649),
.B(n_574),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_609),
.A2(n_585),
.B1(n_524),
.B2(n_541),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_643),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_602),
.A2(n_476),
.B1(n_592),
.B2(n_580),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_626),
.B(n_528),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_642),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_597),
.B(n_594),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_667),
.A2(n_541),
.B(n_528),
.C(n_567),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_625),
.A2(n_596),
.B(n_589),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_656),
.B(n_524),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_662),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_620),
.B(n_557),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_620),
.B(n_557),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_621),
.B(n_577),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_648),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_711),
.A2(n_580),
.B1(n_582),
.B2(n_590),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_645),
.B(n_582),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_600),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_716),
.A2(n_588),
.B1(n_573),
.B2(n_470),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_644),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_645),
.B(n_540),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_720),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_662),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_675),
.Y(n_758)
);

AND2x2_ASAP7_75t_SL g759 ( 
.A(n_675),
.B(n_595),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_639),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_610),
.B(n_514),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_619),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_622),
.B(n_40),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_646),
.B(n_650),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_617),
.A2(n_638),
.B(n_702),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_641),
.B(n_40),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_601),
.A2(n_706),
.B1(n_718),
.B2(n_680),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_539),
.C(n_546),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_679),
.B(n_41),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_664),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_611),
.B(n_42),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_601),
.A2(n_680),
.B1(n_704),
.B2(n_670),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_658),
.A2(n_661),
.B(n_659),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_627),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_719),
.A2(n_550),
.B(n_540),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_663),
.B(n_42),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_666),
.B(n_43),
.Y(n_777)
);

AO21x1_ASAP7_75t_L g778 ( 
.A1(n_697),
.A2(n_599),
.B(n_532),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_657),
.B(n_43),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_618),
.B(n_44),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_659),
.A2(n_559),
.B(n_526),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_670),
.A2(n_709),
.B1(n_721),
.B2(n_712),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_713),
.A2(n_559),
.B1(n_526),
.B2(n_512),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_653),
.Y(n_784)
);

AO22x1_ASAP7_75t_L g785 ( 
.A1(n_619),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_624),
.B(n_630),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_615),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_672),
.B(n_54),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_54),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_669),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_668),
.B(n_55),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_714),
.A2(n_655),
.B(n_654),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_698),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_714),
.A2(n_56),
.B1(n_511),
.B2(n_70),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_603),
.B(n_56),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_714),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_665),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_612),
.B(n_100),
.Y(n_799)
);

BUFx12f_ASAP7_75t_L g800 ( 
.A(n_705),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_636),
.B(n_640),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_652),
.A2(n_102),
.B(n_110),
.Y(n_802)
);

OAI21xp33_ASAP7_75t_L g803 ( 
.A1(n_717),
.A2(n_113),
.B(n_115),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_688),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_693),
.A2(n_138),
.B(n_139),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_637),
.B(n_140),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_651),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_703),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.Y(n_808)
);

AND2x2_ASAP7_75t_SL g809 ( 
.A(n_691),
.B(n_154),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_674),
.A2(n_159),
.B(n_161),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_678),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_660),
.B(n_162),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_676),
.A2(n_168),
.B(n_169),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_694),
.A2(n_180),
.B(n_185),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_623),
.A2(n_628),
.B(n_632),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_660),
.B(n_193),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_692),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_629),
.A2(n_199),
.B(n_200),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_631),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_722),
.A2(n_699),
.B(n_696),
.C(n_686),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_682),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_SL g822 ( 
.A(n_700),
.B(n_684),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_685),
.A2(n_708),
.B1(n_710),
.B2(n_715),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_634),
.B(n_687),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_683),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_683),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_695),
.B(n_686),
.Y(n_827)
);

AOI21xp33_ASAP7_75t_L g828 ( 
.A1(n_734),
.A2(n_733),
.B(n_729),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_766),
.B(n_777),
.C(n_776),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_726),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_730),
.A2(n_748),
.B(n_746),
.C(n_747),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_744),
.A2(n_727),
.B1(n_737),
.B2(n_764),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_728),
.A2(n_750),
.B1(n_753),
.B2(n_732),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_SL g834 ( 
.A(n_758),
.B(n_756),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_731),
.B(n_728),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_792),
.A2(n_742),
.B(n_740),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_SL g837 ( 
.A(n_800),
.B(n_774),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_811),
.B(n_723),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_822),
.B(n_820),
.C(n_771),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_754),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_SL g841 ( 
.A(n_807),
.B(n_767),
.C(n_770),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_749),
.B(n_763),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_762),
.B(n_767),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_735),
.A2(n_817),
.B1(n_796),
.B2(n_738),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_796),
.A2(n_794),
.B1(n_790),
.B2(n_791),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_759),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_793),
.B(n_809),
.Y(n_847)
);

AO31x2_ASAP7_75t_L g848 ( 
.A1(n_823),
.A2(n_795),
.A3(n_808),
.B(n_802),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_789),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_782),
.A2(n_741),
.B(n_812),
.C(n_772),
.Y(n_850)
);

AND2x6_ASAP7_75t_SL g851 ( 
.A(n_789),
.B(n_779),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_825),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_769),
.A2(n_750),
.B1(n_801),
.B2(n_788),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_751),
.B(n_819),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_826),
.B(n_821),
.Y(n_855)
);

AO31x2_ASAP7_75t_L g856 ( 
.A1(n_810),
.A2(n_813),
.A3(n_806),
.B(n_805),
.Y(n_856)
);

AO31x2_ASAP7_75t_L g857 ( 
.A1(n_818),
.A2(n_814),
.A3(n_780),
.B(n_815),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_827),
.A2(n_824),
.B1(n_789),
.B2(n_816),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_799),
.A2(n_804),
.B1(n_798),
.B2(n_755),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_787),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_797),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_768),
.A2(n_783),
.B(n_761),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_725),
.A2(n_739),
.B1(n_745),
.B2(n_757),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_798),
.B(n_785),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_752),
.A2(n_551),
.B1(n_530),
.B2(n_543),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_760),
.A2(n_730),
.B(n_729),
.C(n_746),
.Y(n_866)
);

AOI221x1_ASAP7_75t_L g867 ( 
.A1(n_784),
.A2(n_773),
.B1(n_765),
.B2(n_781),
.C(n_803),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_743),
.B(n_600),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_726),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_730),
.A2(n_765),
.B(n_724),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_766),
.B(n_777),
.C(n_776),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_726),
.Y(n_872)
);

AO31x2_ASAP7_75t_L g873 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_726),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_730),
.A2(n_765),
.B(n_724),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_730),
.A2(n_765),
.B(n_724),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_744),
.B(n_572),
.Y(n_877)
);

CKINVDCx12_ASAP7_75t_R g878 ( 
.A(n_789),
.Y(n_878)
);

CKINVDCx11_ASAP7_75t_R g879 ( 
.A(n_726),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_726),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_744),
.B(n_572),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_730),
.A2(n_765),
.B(n_724),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_726),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_734),
.B(n_656),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_726),
.Y(n_885)
);

AO31x2_ASAP7_75t_L g886 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_886)
);

AO31x2_ASAP7_75t_L g887 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_737),
.B(n_607),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_736),
.Y(n_889)
);

AO31x2_ASAP7_75t_L g890 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_744),
.B(n_572),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_744),
.B(n_572),
.Y(n_892)
);

AO31x2_ASAP7_75t_L g893 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_893)
);

AO31x2_ASAP7_75t_L g894 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_729),
.A2(n_786),
.B(n_746),
.C(n_748),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_729),
.A2(n_786),
.B(n_746),
.C(n_748),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_734),
.B(n_656),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_729),
.A2(n_786),
.B(n_746),
.C(n_748),
.Y(n_898)
);

AO31x2_ASAP7_75t_L g899 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_734),
.B(n_656),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_817),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_817),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_726),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

NAND3x1_ASAP7_75t_L g906 ( 
.A(n_809),
.B(n_525),
.C(n_706),
.Y(n_906)
);

OAI22x1_ASAP7_75t_L g907 ( 
.A1(n_770),
.A2(n_607),
.B1(n_609),
.B2(n_720),
.Y(n_907)
);

OAI22x1_ASAP7_75t_L g908 ( 
.A1(n_770),
.A2(n_607),
.B1(n_609),
.B2(n_720),
.Y(n_908)
);

AO21x2_ASAP7_75t_L g909 ( 
.A1(n_773),
.A2(n_781),
.B(n_765),
.Y(n_909)
);

BUFx4_ASAP7_75t_SL g910 ( 
.A(n_774),
.Y(n_910)
);

AO31x2_ASAP7_75t_L g911 ( 
.A1(n_775),
.A2(n_765),
.A3(n_730),
.B(n_778),
.Y(n_911)
);

AOI221xp5_ASAP7_75t_L g912 ( 
.A1(n_727),
.A2(n_579),
.B1(n_581),
.B2(n_656),
.C(n_520),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_734),
.B(n_656),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_726),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_726),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_744),
.B(n_572),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_765),
.B(n_724),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_734),
.B(n_656),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_723),
.B(n_645),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_726),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_729),
.A2(n_786),
.B(n_746),
.C(n_748),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_830),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_840),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_879),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_852),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_SL g926 ( 
.A1(n_895),
.A2(n_898),
.B(n_896),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_889),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_860),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_897),
.B(n_901),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_854),
.B(n_900),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_913),
.B(n_918),
.Y(n_931)
);

OA21x2_ASAP7_75t_L g932 ( 
.A1(n_876),
.A2(n_917),
.B(n_882),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_828),
.A2(n_912),
.B1(n_832),
.B2(n_865),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_845),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_874),
.Y(n_935)
);

CKINVDCx11_ASAP7_75t_R g936 ( 
.A(n_914),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_880),
.Y(n_937)
);

AO31x2_ASAP7_75t_L g938 ( 
.A1(n_862),
.A2(n_850),
.A3(n_833),
.B(n_836),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_855),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_900),
.Y(n_940)
);

OAI222xp33_ASAP7_75t_L g941 ( 
.A1(n_849),
.A2(n_846),
.B1(n_844),
.B2(n_853),
.C1(n_842),
.C2(n_888),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_861),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_878),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_839),
.A2(n_877),
.B(n_916),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_883),
.Y(n_945)
);

BUFx2_ASAP7_75t_R g946 ( 
.A(n_905),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_881),
.A2(n_892),
.B(n_891),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_910),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_858),
.B(n_866),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_859),
.B(n_843),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_914),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_869),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_873),
.A2(n_886),
.B(n_899),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_864),
.A2(n_847),
.B(n_834),
.C(n_903),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_904),
.B(n_915),
.Y(n_955)
);

BUFx4f_ASAP7_75t_SL g956 ( 
.A(n_920),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_902),
.A2(n_863),
.B(n_841),
.C(n_838),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_872),
.Y(n_958)
);

AO31x2_ASAP7_75t_L g959 ( 
.A1(n_873),
.A2(n_886),
.A3(n_911),
.B(n_899),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_906),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_908),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_909),
.A2(n_868),
.B(n_907),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_887),
.A2(n_899),
.B(n_894),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_851),
.B(n_885),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_837),
.B(n_887),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_890),
.A2(n_893),
.B(n_911),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_848),
.B(n_857),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_893),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_848),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_856),
.B(n_835),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_870),
.A2(n_876),
.B(n_875),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_829),
.B(n_871),
.C(n_839),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_835),
.A2(n_828),
.B1(n_912),
.B2(n_832),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_861),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_880),
.B(n_607),
.Y(n_975)
);

OA21x2_ASAP7_75t_L g976 ( 
.A1(n_867),
.A2(n_875),
.B(n_870),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_884),
.B(n_656),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_835),
.B(n_744),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_895),
.A2(n_898),
.B(n_896),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_879),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_840),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_870),
.A2(n_876),
.B(n_875),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_840),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_858),
.B(n_839),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_831),
.A2(n_921),
.B(n_895),
.C(n_898),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_928),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_970),
.B(n_978),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_954),
.B(n_950),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_SL g989 ( 
.A1(n_960),
.A2(n_951),
.B1(n_934),
.B2(n_939),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_925),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_979),
.B(n_985),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_926),
.B(n_973),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_944),
.A2(n_972),
.B(n_947),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_973),
.B(n_984),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_971),
.B(n_982),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_940),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_923),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_971),
.B(n_982),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_932),
.B(n_938),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_932),
.B(n_938),
.Y(n_1000)
);

BUFx5_ASAP7_75t_L g1001 ( 
.A(n_930),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_927),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_981),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_983),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_940),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_932),
.B(n_938),
.Y(n_1006)
);

AO31x2_ASAP7_75t_L g1007 ( 
.A1(n_967),
.A2(n_969),
.A3(n_968),
.B(n_962),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_938),
.B(n_963),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_963),
.B(n_953),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_996),
.B(n_965),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_1001),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_1001),
.Y(n_1013)
);

OAI211xp5_ASAP7_75t_SL g1014 ( 
.A1(n_989),
.A2(n_931),
.B(n_929),
.C(n_964),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_991),
.B(n_949),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_992),
.A2(n_933),
.B1(n_977),
.B2(n_950),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_967),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_990),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1009),
.B(n_953),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_1001),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_999),
.B(n_1000),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_987),
.B(n_959),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_1005),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_989),
.A2(n_933),
.B1(n_954),
.B2(n_957),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_987),
.B(n_959),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_996),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_986),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_999),
.B(n_966),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_1006),
.B(n_959),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_995),
.B(n_976),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_1029),
.B(n_1028),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1015),
.B(n_997),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1022),
.B(n_995),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1010),
.B(n_998),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1027),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1023),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_1018),
.B(n_996),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_987),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_1026),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1021),
.B(n_1002),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1010),
.B(n_1007),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_1012),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_1039),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1036),
.B(n_1014),
.C(n_1024),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1035),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1035),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_1011),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1038),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1040),
.B(n_1042),
.Y(n_1051)
);

NAND2x1_ASAP7_75t_SL g1052 ( 
.A(n_1031),
.B(n_980),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1034),
.B(n_1021),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1034),
.B(n_1021),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1043),
.B(n_1017),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_1032),
.B(n_1014),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1043),
.B(n_1019),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1031),
.B(n_1011),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1033),
.B(n_1025),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1057),
.B(n_1031),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1052),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_1046),
.B(n_1024),
.C(n_993),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1053),
.B(n_1037),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1057),
.B(n_1031),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1047),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1048),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1053),
.B(n_1030),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_1045),
.A2(n_948),
.B(n_951),
.C(n_1056),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_1049),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1058),
.B(n_924),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1050),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1056),
.B(n_980),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1054),
.B(n_1041),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_1059),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1071),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_1069),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1061),
.B(n_946),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1074),
.B(n_1054),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1071),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1071),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1061),
.A2(n_1058),
.B1(n_1049),
.B2(n_1020),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1060),
.B(n_1058),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1065),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_1051),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1065),
.Y(n_1086)
);

INVxp33_ASAP7_75t_L g1087 ( 
.A(n_1070),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1068),
.A2(n_1049),
.B(n_1044),
.Y(n_1088)
);

OAI221xp5_ASAP7_75t_L g1089 ( 
.A1(n_1077),
.A2(n_1062),
.B1(n_1072),
.B2(n_1069),
.C(n_1073),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_1088),
.B(n_924),
.C(n_935),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1081),
.A2(n_1049),
.B(n_1063),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1087),
.A2(n_1029),
.B1(n_991),
.B2(n_1028),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1083),
.Y(n_1093)
);

AOI221x1_ASAP7_75t_L g1094 ( 
.A1(n_1076),
.A2(n_993),
.B1(n_1066),
.B2(n_1004),
.C(n_1003),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1076),
.A2(n_1067),
.B(n_1055),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1076),
.A2(n_1059),
.B1(n_1013),
.B2(n_1012),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_1094),
.B(n_1089),
.C(n_1092),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1096),
.A2(n_1076),
.B(n_955),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1090),
.A2(n_1083),
.B1(n_1086),
.B2(n_1078),
.C(n_1085),
.Y(n_1099)
);

OAI211xp5_ASAP7_75t_L g1100 ( 
.A1(n_1091),
.A2(n_936),
.B(n_1016),
.C(n_992),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_1095),
.B(n_936),
.C(n_943),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_1086),
.B1(n_1079),
.B2(n_1080),
.C(n_961),
.Y(n_1102)
);

AOI221x1_ASAP7_75t_L g1103 ( 
.A1(n_1090),
.A2(n_1079),
.B1(n_1080),
.B2(n_957),
.C(n_1066),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_1089),
.A2(n_1016),
.B1(n_1082),
.B2(n_1075),
.C(n_988),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_SL g1105 ( 
.A1(n_1100),
.A2(n_941),
.B(n_955),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1099),
.B(n_1101),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1102),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1103),
.B(n_1085),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1097),
.A2(n_991),
.B(n_942),
.Y(n_1109)
);

NAND4xp75_ASAP7_75t_L g1110 ( 
.A(n_1104),
.B(n_988),
.C(n_1082),
.D(n_994),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1106),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_1084),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1108),
.A2(n_1106),
.B1(n_1110),
.B2(n_1105),
.Y(n_1113)
);

XNOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1107),
.B(n_937),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_1109),
.B(n_1098),
.C(n_935),
.Y(n_1115)
);

NOR3x1_ASAP7_75t_L g1116 ( 
.A(n_1109),
.B(n_922),
.C(n_952),
.Y(n_1116)
);

XNOR2xp5_ASAP7_75t_L g1117 ( 
.A(n_1114),
.B(n_975),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_L g1118 ( 
.A(n_1115),
.B(n_974),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1113),
.A2(n_1064),
.B1(n_1084),
.B2(n_945),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1111),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1116),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1120),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1121),
.Y(n_1123)
);

AOI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_1123),
.B1(n_1117),
.B2(n_945),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1124),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1125),
.B(n_1123),
.Y(n_1126)
);

AOI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1126),
.A2(n_1118),
.B(n_1119),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1128),
.A2(n_1112),
.B1(n_956),
.B2(n_958),
.Y(n_1129)
);


endmodule