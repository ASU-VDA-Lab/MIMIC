module fake_aes_176_n_669 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_669);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_27), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_76), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_0), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_54), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_77), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_38), .Y(n_84) );
CKINVDCx14_ASAP7_75t_R g85 ( .A(n_7), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_30), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_57), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_5), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_8), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_36), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_14), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_4), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_28), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_75), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_2), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_74), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_33), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_24), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_73), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_6), .Y(n_110) );
BUFx5_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_55), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_69), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_23), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_42), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_9), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_24), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_37), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_91), .B(n_1), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_85), .B(n_1), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_98), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_122), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
NAND2xp33_ASAP7_75t_R g139 ( .A(n_79), .B(n_2), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_108), .B(n_29), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_111), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_108), .B(n_26), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_120), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_103), .B(n_3), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_97), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_91), .B(n_4), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_123), .B(n_5), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_88), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_79), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_111), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_86), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_86), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_88), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_88), .Y(n_166) );
NOR2xp33_ASAP7_75t_R g167 ( .A(n_94), .B(n_34), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_111), .B(n_6), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_127), .A2(n_124), .B(n_123), .C(n_106), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_127), .B(n_82), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_132), .B(n_116), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g172 ( .A(n_154), .B(n_116), .C(n_96), .Y(n_172) );
AO22x2_ASAP7_75t_L g173 ( .A1(n_130), .A2(n_124), .B1(n_105), .B2(n_112), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_132), .B(n_114), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_130), .A2(n_119), .B1(n_80), .B2(n_118), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_134), .A2(n_119), .B1(n_115), .B2(n_100), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_134), .B(n_102), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_129), .B(n_102), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_130), .B(n_121), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_148), .B(n_156), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_154), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_159), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_129), .B(n_117), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_135), .B(n_114), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_148), .B(n_113), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
AO22x2_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_83), .B1(n_84), .B2(n_109), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_153), .B(n_94), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_135), .B(n_107), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_137), .B(n_99), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_142), .B(n_104), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_142), .B(n_101), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_150), .B(n_111), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g208 ( .A(n_128), .B(n_151), .C(n_168), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_152), .B(n_111), .Y(n_209) );
NOR2x1p5_ASAP7_75t_L g210 ( .A(n_131), .B(n_95), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_157), .B(n_88), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_160), .B(n_8), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_160), .B(n_40), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_161), .B(n_35), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_126), .B(n_9), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_128), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_161), .B(n_10), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_165), .B(n_10), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
INVx6_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_168), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_154), .B(n_45), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_143), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_133), .B(n_12), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_162), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_141), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_165), .B(n_49), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_139), .B(n_16), .C(n_17), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_165), .B(n_17), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_136), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_222), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_222), .Y(n_235) );
NOR3xp33_ASAP7_75t_SL g236 ( .A(n_184), .B(n_177), .C(n_171), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_217), .B(n_147), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_219), .B(n_126), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_179), .B(n_126), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_188), .B(n_140), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_178), .B(n_140), .Y(n_242) );
NOR2xp33_ASAP7_75t_R g243 ( .A(n_184), .B(n_149), .Y(n_243) );
BUFx4f_ASAP7_75t_L g244 ( .A(n_180), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_183), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_183), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_193), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_220), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_186), .B(n_195), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_232), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_186), .B(n_140), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_175), .B(n_144), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_186), .B(n_167), .Y(n_254) );
BUFx8_ASAP7_75t_L g255 ( .A(n_226), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_187), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_195), .B(n_167), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_182), .B(n_141), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_187), .Y(n_259) );
AND3x1_ASAP7_75t_SL g260 ( .A(n_210), .B(n_18), .C(n_19), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_176), .Y(n_262) );
OAI221xp5_ASAP7_75t_L g263 ( .A1(n_169), .A2(n_158), .B1(n_146), .B2(n_144), .C(n_162), .Y(n_263) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
NOR2xp33_ASAP7_75t_R g265 ( .A(n_182), .B(n_141), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_190), .B(n_144), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_190), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_190), .B(n_158), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_185), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_191), .B(n_158), .Y(n_273) );
NOR2xp33_ASAP7_75t_R g274 ( .A(n_199), .B(n_141), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_190), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
NOR3xp33_ASAP7_75t_SL g277 ( .A(n_169), .B(n_18), .C(n_19), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_208), .B(n_146), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_192), .A2(n_145), .B1(n_141), .B2(n_146), .Y(n_280) );
OR2x6_ASAP7_75t_SL g281 ( .A(n_230), .B(n_20), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_195), .B(n_145), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_173), .B(n_20), .Y(n_283) );
INVx6_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
BUFx4f_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_231), .Y(n_286) );
BUFx12f_ASAP7_75t_L g287 ( .A(n_213), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_170), .A2(n_162), .B(n_164), .C(n_166), .Y(n_288) );
NOR3xp33_ASAP7_75t_SL g289 ( .A(n_170), .B(n_21), .C(n_22), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_197), .B(n_145), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_218), .B(n_231), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_176), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_198), .B(n_145), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_202), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_173), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_218), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_200), .B(n_141), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_203), .B(n_166), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_278), .A2(n_206), .B(n_211), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_269), .A2(n_173), .B1(n_192), .B2(n_223), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_243), .Y(n_304) );
BUFx4_ASAP7_75t_SL g305 ( .A(n_251), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_272), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_245), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_269), .B(n_192), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_247), .B(n_172), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_296), .A2(n_194), .B(n_201), .C(n_209), .Y(n_310) );
OAI21x1_ASAP7_75t_SL g311 ( .A1(n_280), .A2(n_228), .B(n_204), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_291), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_250), .B(n_202), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_224), .B(n_216), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_292), .A2(n_223), .B1(n_228), .B2(n_224), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_287), .Y(n_317) );
INVx5_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_294), .B(n_221), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_238), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_291), .B(n_225), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_287), .A2(n_223), .B1(n_207), .B2(n_225), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_248), .B(n_214), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_243), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_291), .B(n_225), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_271), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_285), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_285), .B(n_214), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_239), .A2(n_212), .B(n_229), .C(n_215), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_282), .A2(n_229), .B(n_215), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_270), .B(n_145), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_251), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_237), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_244), .B(n_22), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_270), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_252), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_284), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_245), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
AND2x6_ASAP7_75t_L g344 ( .A(n_295), .B(n_141), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_275), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_253), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_267), .B(n_145), .Y(n_347) );
BUFx12f_ASAP7_75t_L g348 ( .A(n_255), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_244), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_256), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_284), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_284), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_331), .A2(n_266), .B(n_249), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_326), .Y(n_354) );
AND2x6_ASAP7_75t_L g355 ( .A(n_332), .B(n_295), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_308), .B(n_264), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_320), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_339), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_308), .A2(n_286), .B1(n_261), .B2(n_295), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_315), .A2(n_261), .B(n_286), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_308), .A2(n_264), .B1(n_283), .B2(n_255), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_313), .B(n_236), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_318), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_346), .B(n_257), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_303), .A2(n_255), .B1(n_242), .B2(n_254), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g366 ( .A1(n_334), .A2(n_242), .B(n_253), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_343), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_333), .B(n_246), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_301), .A2(n_290), .B(n_293), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_329), .A2(n_298), .B(n_273), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_308), .A2(n_281), .B1(n_246), .B2(n_234), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_345), .B(n_273), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_307), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_310), .A2(n_300), .B(n_240), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_309), .A2(n_241), .B(n_263), .Y(n_375) );
CKINVDCx6p67_ASAP7_75t_R g376 ( .A(n_348), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_302), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_306), .A2(n_259), .B1(n_279), .B2(n_268), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_348), .A2(n_304), .B1(n_324), .B2(n_335), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_312), .A2(n_259), .B1(n_279), .B2(n_268), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_327), .B(n_234), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_325), .B(n_276), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_345), .B(n_276), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_365), .A2(n_322), .B(n_289), .C(n_316), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_361), .A2(n_323), .B1(n_304), .B2(n_324), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_325), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_319), .B(n_277), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_371), .B(n_330), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_380), .B(n_317), .C(n_260), .D(n_288), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_337), .B1(n_336), .B2(n_338), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_383), .B(n_312), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
NAND2x1_ASAP7_75t_L g394 ( .A(n_373), .B(n_307), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_372), .A2(n_352), .B1(n_327), .B2(n_311), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_372), .B(n_317), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_328), .B1(n_349), .B2(n_327), .C(n_351), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_332), .B1(n_321), .B2(n_352), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_383), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_354), .A2(n_305), .B1(n_340), .B2(n_318), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_370), .B(n_353), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_377), .A2(n_311), .B1(n_340), .B2(n_332), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_378), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_384), .A2(n_288), .B1(n_298), .B2(n_342), .C(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_356), .B(n_314), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_384), .A2(n_347), .B1(n_350), .B2(n_314), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_354), .A2(n_318), .B1(n_234), .B2(n_342), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_356), .B(n_342), .Y(n_412) );
NAND2xp33_ASAP7_75t_R g413 ( .A(n_399), .B(n_377), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_393), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_395), .B(n_355), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_397), .B(n_355), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_355), .B1(n_375), .B2(n_368), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_385), .A2(n_376), .B1(n_379), .B2(n_381), .C(n_363), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_393), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_355), .B1(n_376), .B2(n_347), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_408), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_408), .B(n_363), .Y(n_425) );
AOI211xp5_ASAP7_75t_SL g426 ( .A1(n_403), .A2(n_382), .B(n_347), .C(n_330), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_396), .A2(n_355), .B1(n_382), .B2(n_374), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_405), .A2(n_355), .B1(n_382), .B2(n_344), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_402), .B(n_373), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_404), .B(n_164), .C(n_166), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
INVx5_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_398), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_386), .B(n_23), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_391), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_406), .A2(n_373), .B1(n_318), .B2(n_330), .Y(n_440) );
AND2x6_ASAP7_75t_SL g441 ( .A(n_406), .B(n_344), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
AOI33xp33_ASAP7_75t_L g443 ( .A1(n_398), .A2(n_189), .A3(n_227), .B1(n_205), .B2(n_164), .B3(n_166), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_387), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_392), .B(n_373), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_410), .A2(n_374), .B1(n_318), .B2(n_344), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_412), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_445), .B(n_389), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_424), .B(n_401), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_444), .B(n_400), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_419), .B(n_369), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_437), .B(n_407), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_440), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_431), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_444), .B(n_411), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_440), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_431), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_424), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_445), .B(n_166), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_437), .B(n_369), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_446), .B(n_341), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_307), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_446), .B(n_166), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_427), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_422), .B(n_25), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_166), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_448), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_442), .B(n_164), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_439), .B(n_341), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_436), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_442), .B(n_164), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_427), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_442), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_436), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_414), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_439), .Y(n_485) );
NOR2x1p5_ASAP7_75t_L g486 ( .A(n_430), .B(n_341), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_414), .B(n_164), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_419), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_421), .B(n_164), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_421), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_415), .B(n_341), .Y(n_492) );
NAND4xp25_ASAP7_75t_SL g493 ( .A(n_423), .B(n_31), .C(n_43), .D(n_46), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_438), .A2(n_300), .B1(n_155), .B2(n_307), .C(n_341), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_436), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_421), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_420), .B(n_155), .C(n_307), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_436), .B(n_155), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_461), .B(n_435), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_456), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_488), .B(n_419), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_474), .B(n_436), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_456), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_449), .B(n_435), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
AND2x4_ASAP7_75t_SL g506 ( .A(n_477), .B(n_425), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_488), .B(n_419), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_449), .B(n_436), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_461), .B(n_433), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_485), .B(n_433), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_455), .B(n_436), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_452), .B(n_415), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_481), .B(n_417), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_472), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_454), .B(n_417), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_454), .B(n_425), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_458), .B(n_428), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_450), .B(n_428), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_460), .B(n_420), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_462), .B(n_447), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_471), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_483), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_450), .B(n_426), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_497), .A2(n_413), .B1(n_418), .B2(n_429), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_484), .B(n_426), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_478), .B(n_447), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_478), .B(n_155), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_497), .A2(n_434), .B1(n_145), .B2(n_141), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_479), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_482), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_484), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_489), .B(n_443), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_471), .B(n_155), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_489), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_486), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_491), .B(n_155), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_457), .B(n_434), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_496), .B(n_441), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_479), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_477), .B(n_344), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_496), .B(n_141), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_463), .B(n_47), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_468), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_463), .B(n_50), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_468), .B(n_145), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_505), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_517), .A2(n_494), .B(n_476), .C(n_455), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_512), .A2(n_459), .B(n_493), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_523), .B(n_453), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_512), .B(n_477), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_529), .A2(n_459), .B1(n_457), .B2(n_464), .C(n_495), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_514), .B(n_465), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_506), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_502), .A2(n_498), .B(n_495), .Y(n_564) );
NOR3xp33_ASAP7_75t_SL g565 ( .A(n_528), .B(n_465), .C(n_466), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_506), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_519), .B(n_483), .Y(n_567) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_543), .B(n_486), .Y(n_568) );
OAI22xp33_ASAP7_75t_SL g569 ( .A1(n_543), .A2(n_477), .B1(n_488), .B2(n_467), .Y(n_569) );
OAI322xp33_ASAP7_75t_L g570 ( .A1(n_522), .A2(n_467), .A3(n_492), .B1(n_473), .B2(n_475), .C1(n_480), .C2(n_498), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_513), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_521), .A2(n_473), .B1(n_480), .B2(n_475), .C1(n_453), .C2(n_487), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_518), .B(n_492), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_504), .B(n_453), .Y(n_575) );
OAI322xp33_ASAP7_75t_L g576 ( .A1(n_522), .A2(n_490), .A3(n_487), .B1(n_196), .B2(n_205), .C1(n_227), .C2(n_189), .Y(n_576) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_537), .A2(n_490), .A3(n_453), .B1(n_235), .B2(n_60), .Y(n_577) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_548), .Y(n_578) );
OA211x2_ASAP7_75t_L g579 ( .A1(n_549), .A2(n_52), .B(n_53), .C(n_56), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_501), .B(n_274), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_540), .B(n_196), .C(n_234), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_504), .B(n_61), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_509), .B(n_62), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_526), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_526), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_545), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_520), .A2(n_145), .B1(n_344), .B2(n_274), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_499), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_552), .B(n_63), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_530), .A2(n_344), .B1(n_196), .B2(n_258), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_547), .A2(n_235), .B1(n_233), .B2(n_67), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_511), .B(n_64), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_515), .B(n_66), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_511), .B(n_71), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_531), .Y(n_595) );
AOI33xp33_ASAP7_75t_L g596 ( .A1(n_523), .A2(n_196), .A3(n_233), .B1(n_258), .B2(n_265), .B3(n_532), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_500), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_536), .Y(n_598) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_551), .B(n_233), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_588), .B(n_532), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g602 ( .A1(n_586), .A2(n_556), .A3(n_566), .B1(n_563), .B2(n_578), .C1(n_559), .C2(n_568), .Y(n_602) );
XNOR2xp5_ASAP7_75t_L g603 ( .A(n_599), .B(n_515), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_559), .B(n_501), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g606 ( .A1(n_561), .A2(n_538), .B1(n_539), .B2(n_542), .C1(n_546), .C2(n_551), .Y(n_606) );
AOI322xp5_ASAP7_75t_L g607 ( .A1(n_568), .A2(n_525), .A3(n_553), .B1(n_508), .B2(n_533), .C1(n_544), .C2(n_535), .Y(n_607) );
NAND2xp33_ASAP7_75t_L g608 ( .A(n_565), .B(n_545), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_562), .B(n_510), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g610 ( .A(n_558), .B(n_554), .C(n_550), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_598), .Y(n_611) );
NOR3xp33_ASAP7_75t_SL g612 ( .A(n_570), .B(n_508), .C(n_499), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_574), .B(n_510), .Y(n_613) );
NOR2xp33_ASAP7_75t_R g614 ( .A(n_593), .B(n_553), .Y(n_614) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_557), .A2(n_535), .B(n_533), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_575), .B(n_527), .Y(n_616) );
AOI222xp33_ASAP7_75t_SL g617 ( .A1(n_595), .A2(n_535), .B1(n_503), .B2(n_516), .C1(n_524), .C2(n_534), .Y(n_617) );
NAND2xp33_ASAP7_75t_R g618 ( .A(n_593), .B(n_544), .Y(n_618) );
AOI31xp33_ASAP7_75t_L g619 ( .A1(n_560), .A2(n_503), .A3(n_516), .B(n_524), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_571), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
NAND3xp33_ASAP7_75t_SL g622 ( .A(n_560), .B(n_541), .C(n_233), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_573), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_584), .B(n_541), .Y(n_624) );
NOR4xp25_ASAP7_75t_SL g625 ( .A(n_580), .B(n_585), .C(n_599), .D(n_569), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_567), .B(n_592), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_564), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_589), .Y(n_628) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_597), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_612), .B(n_583), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_623), .B(n_594), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_602), .B(n_596), .C(n_582), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_627), .B(n_596), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_605), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_609), .B(n_581), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_608), .B(n_591), .C(n_577), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_603), .B(n_579), .Y(n_638) );
OAI211xp5_ASAP7_75t_SL g639 ( .A1(n_606), .A2(n_590), .B(n_580), .C(n_587), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_608), .A2(n_576), .B1(n_590), .B2(n_587), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_616), .B(n_604), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_607), .A2(n_600), .B1(n_626), .B2(n_613), .C(n_625), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_619), .A2(n_622), .B(n_615), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_611), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_626), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_631), .A2(n_610), .B(n_620), .C(n_621), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_618), .B1(n_617), .B2(n_628), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_643), .A2(n_618), .B1(n_629), .B2(n_628), .Y(n_648) );
INVx5_ASAP7_75t_L g649 ( .A(n_630), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_635), .Y(n_650) );
OAI31xp33_ASAP7_75t_L g651 ( .A1(n_642), .A2(n_624), .A3(n_614), .B(n_628), .Y(n_651) );
OAI221xp5_ASAP7_75t_SL g652 ( .A1(n_637), .A2(n_640), .B1(n_645), .B2(n_632), .C(n_636), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_640), .B(n_639), .C(n_630), .Y(n_653) );
OAI321xp33_ASAP7_75t_L g654 ( .A1(n_634), .A2(n_642), .A3(n_623), .B1(n_632), .B2(n_635), .C(n_633), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_644), .A2(n_637), .B(n_642), .Y(n_655) );
AO211x2_ASAP7_75t_L g656 ( .A1(n_641), .A2(n_632), .B(n_637), .C(n_633), .Y(n_656) );
AOI21xp33_ASAP7_75t_SL g657 ( .A1(n_642), .A2(n_637), .B(n_638), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_649), .B(n_651), .Y(n_658) );
NOR3x1_ASAP7_75t_L g659 ( .A(n_653), .B(n_655), .C(n_656), .Y(n_659) );
OR3x2_ASAP7_75t_L g660 ( .A(n_657), .B(n_652), .C(n_654), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_650), .Y(n_661) );
OR3x1_ASAP7_75t_L g662 ( .A(n_660), .B(n_646), .C(n_652), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_661), .B(n_649), .C(n_647), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_659), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_664), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_662), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_666), .B1(n_663), .B2(n_658), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_648), .B(n_649), .Y(n_669) );
endmodule