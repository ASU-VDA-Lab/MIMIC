module fake_jpeg_7758_n_88 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_62),
.B1(n_51),
.B2(n_52),
.Y(n_73)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_6),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_53),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_75),
.B(n_71),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_78),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_70),
.C(n_42),
.Y(n_81)
);

OAI322xp33_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_45),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_9),
.B(n_18),
.C(n_19),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_21),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.C1(n_26),
.C2(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_36),
.C(n_31),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_29),
.C(n_32),
.Y(n_88)
);


endmodule