module fake_jpeg_17024_n_144 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_25),
.B1(n_8),
.B2(n_10),
.Y(n_51)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_18),
.A2(n_1),
.B1(n_13),
.B2(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_24),
.B1(n_20),
.B2(n_28),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_24),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_45),
.B(n_51),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_26),
.B(n_15),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_32),
.C(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_31),
.B(n_30),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_58),
.C(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_68),
.Y(n_83)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_30),
.C(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_50),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_37),
.B(n_35),
.C(n_33),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_29),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_37),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_58),
.B1(n_69),
.B2(n_54),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_93),
.B1(n_101),
.B2(n_82),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_60),
.B1(n_55),
.B2(n_71),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_53),
.C(n_21),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_23),
.C(n_27),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_23),
.B(n_27),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_14),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_61),
.B1(n_66),
.B2(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_82),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_6),
.B(n_8),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_108),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_94),
.C(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_119),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_103),
.B1(n_104),
.B2(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_121),
.B(n_110),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_126),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_112),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_132),
.B(n_133),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_119),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_120),
.B(n_108),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_99),
.B(n_106),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_136),
.B(n_137),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_12),
.B(n_81),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_139),
.C(n_78),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_78),
.Y(n_144)
);


endmodule