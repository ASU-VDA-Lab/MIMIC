module fake_jpeg_9972_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_40),
.Y(n_57)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_24),
.Y(n_90)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_62),
.Y(n_84)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_41),
.B1(n_34),
.B2(n_29),
.Y(n_64)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_64),
.B(n_76),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_69),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_28),
.B2(n_16),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_82),
.B1(n_59),
.B2(n_55),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_40),
.C(n_37),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_20),
.C(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_30),
.B1(n_26),
.B2(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_88),
.B1(n_58),
.B2(n_46),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_11),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_115),
.B1(n_65),
.B2(n_79),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_118),
.C(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_90),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_75),
.B1(n_66),
.B2(n_77),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_89),
.B1(n_88),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_55),
.B1(n_47),
.B2(n_37),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_64),
.B(n_20),
.CI(n_32),
.CON(n_117),
.SN(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_90),
.B(n_20),
.C(n_32),
.D(n_21),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_22),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_17),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_96),
.B1(n_2),
.B2(n_3),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_139),
.B1(n_9),
.B2(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_136),
.C(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_146),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_80),
.B1(n_92),
.B2(n_86),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_135),
.B1(n_108),
.B2(n_105),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_80),
.B1(n_86),
.B2(n_66),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_75),
.C(n_72),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_77),
.B1(n_52),
.B2(n_27),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_27),
.B(n_20),
.C(n_32),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_128),
.B(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_95),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_98),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_93),
.B1(n_107),
.B2(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_17),
.C(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_119),
.B1(n_117),
.B2(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_158),
.B1(n_175),
.B2(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_117),
.B1(n_120),
.B2(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_160),
.B(n_168),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_165),
.B(n_157),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_116),
.B(n_118),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_172),
.B(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_180),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_116),
.C(n_109),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_174),
.C(n_179),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_96),
.C(n_17),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_96),
.B1(n_21),
.B2(n_20),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_176),
.A2(n_178),
.B1(n_11),
.B2(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_1),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_125),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_145),
.C(n_144),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_10),
.Y(n_192)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_182),
.C(n_167),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_194),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_204),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_141),
.B(n_3),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_207),
.B1(n_209),
.B2(n_162),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_211),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_141),
.B1(n_3),
.B2(n_5),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_141),
.B(n_5),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_11),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_152),
.B1(n_158),
.B2(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_186),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_152),
.B1(n_160),
.B2(n_181),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_164),
.B1(n_159),
.B2(n_151),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_179),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_187),
.C(n_193),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_163),
.C(n_177),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_232),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_174),
.B1(n_6),
.B2(n_2),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_7),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_227),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_202),
.B(n_186),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_251),
.B1(n_253),
.B2(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_187),
.C(n_184),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_255),
.C(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_254),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_210),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_220),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_197),
.B1(n_207),
.B2(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_197),
.B1(n_209),
.B2(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_6),
.C(n_7),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_10),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.C(n_268),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_254),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_237),
.B1(n_250),
.B2(n_240),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_214),
.C(n_213),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_244),
.B(n_253),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_212),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_271),
.Y(n_275)
);

FAx1_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_269),
.CI(n_270),
.CON(n_286),
.SN(n_286)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_242),
.B(n_238),
.C(n_247),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_243),
.C(n_245),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_282),
.B(n_262),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_237),
.B1(n_239),
.B2(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_255),
.C(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_263),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_12),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_221),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_267),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_289),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_273),
.C(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_293),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_274),
.B1(n_14),
.B2(n_15),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_278),
.B(n_12),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_272),
.B(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_300),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_280),
.C(n_274),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_308),
.B(n_302),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_274),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_285),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_307),
.B(n_300),
.CI(n_298),
.CON(n_310),
.SN(n_310)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_305),
.B1(n_311),
.B2(n_307),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_6),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);


endmodule