module fake_jpeg_14648_n_334 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_40),
.B(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_46),
.B(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_24),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_58),
.Y(n_77)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_66),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_18),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_87),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_83),
.B(n_84),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_37),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_31),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_85),
.B(n_3),
.C(n_4),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_93),
.B1(n_106),
.B2(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_38),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_103),
.Y(n_135)
);

INVx2_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_17),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_39),
.B(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_41),
.A2(n_30),
.B1(n_14),
.B2(n_27),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_14),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_63),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_27),
.B1(n_17),
.B2(n_20),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_44),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_43),
.B(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_1),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_121),
.Y(n_159)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_31),
.B1(n_25),
.B2(n_16),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_61),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_45),
.B(n_2),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_57),
.B1(n_56),
.B2(n_31),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_124),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_31),
.B1(n_10),
.B2(n_8),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_143),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_132),
.B(n_157),
.Y(n_195)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

OR2x4_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_52),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_148),
.Y(n_182)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_95),
.B1(n_72),
.B2(n_76),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_10),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_63),
.B(n_3),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_9),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_149),
.Y(n_185)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_9),
.B1(n_16),
.B2(n_25),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_9),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_25),
.B1(n_52),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_113),
.B1(n_88),
.B2(n_104),
.Y(n_168)
);

OR2x4_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_52),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_94),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_45),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_50),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_153),
.Y(n_175)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_2),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_3),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_91),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_96),
.A2(n_69),
.B(n_48),
.C(n_6),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_77),
.B(n_71),
.Y(n_173)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_164),
.Y(n_190)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_173),
.B(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_175),
.B(n_201),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_109),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_201),
.B(n_203),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_118),
.B1(n_102),
.B2(n_112),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_191),
.B1(n_196),
.B2(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_102),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_192),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_111),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_3),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_6),
.B(n_7),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_188),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_144),
.B1(n_129),
.B2(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_76),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_82),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_199),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_122),
.A2(n_72),
.B1(n_95),
.B2(n_78),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_138),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_82),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_126),
.B(n_4),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_73),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_135),
.B(n_4),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_166),
.C(n_159),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_205),
.B(n_207),
.C(n_214),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_206),
.B(n_208),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_135),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_156),
.Y(n_208)
);

INVx6_ASAP7_75t_SL g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_215),
.Y(n_236)
);

HAxp5_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_127),
.CON(n_210),
.SN(n_210)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_229),
.B(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_179),
.B(n_170),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_135),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_130),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_155),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_130),
.C(n_141),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_133),
.B1(n_161),
.B2(n_139),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_188),
.B1(n_196),
.B2(n_136),
.Y(n_260)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_183),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_180),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_163),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_207),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g273 ( 
.A1(n_235),
.A2(n_218),
.A3(n_195),
.B1(n_185),
.B2(n_222),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_237),
.B(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_239),
.B(n_240),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_186),
.B(n_182),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_186),
.B(n_182),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_184),
.B(n_177),
.Y(n_246)
);

AO21x2_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_196),
.B(n_173),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_257),
.B1(n_260),
.B2(n_230),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_254),
.C(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_175),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_178),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_212),
.A2(n_177),
.B(n_179),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_259),
.B(n_195),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_168),
.B1(n_177),
.B2(n_173),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_184),
.B(n_173),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_234),
.B1(n_220),
.B2(n_204),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_267),
.B1(n_270),
.B2(n_275),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_215),
.B1(n_231),
.B2(n_216),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_214),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_219),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_238),
.B(n_249),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_232),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_277),
.C(n_256),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_185),
.C(n_223),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_226),
.C(n_211),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_196),
.B(n_224),
.C(n_206),
.D(n_189),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_259),
.B(n_246),
.C(n_242),
.D(n_260),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_237),
.B(n_209),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_247),
.B(n_244),
.C(n_245),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_248),
.B(n_272),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_292),
.C(n_278),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_282),
.B(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_283),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_250),
.C(n_252),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_243),
.B(n_235),
.C(n_241),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_269),
.B(n_279),
.C(n_261),
.D(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_286),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_307),
.C(n_310),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_263),
.B1(n_248),
.B2(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_308),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_282),
.B1(n_295),
.B2(n_288),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_277),
.C(n_274),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_251),
.B1(n_198),
.B2(n_193),
.Y(n_308)
);

AOI22x1_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_198),
.B1(n_172),
.B2(n_193),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_291),
.B1(n_285),
.B2(n_172),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_171),
.C(n_134),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_315),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_294),
.C(n_297),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_306),
.B(n_309),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_320),
.B(n_301),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_147),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_310),
.B(n_302),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_312),
.A3(n_318),
.B1(n_301),
.B2(n_314),
.C1(n_320),
.C2(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_317),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_327),
.A3(n_322),
.B1(n_317),
.B2(n_165),
.C1(n_134),
.C2(n_78),
.Y(n_332)
);

AOI311xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_330),
.A3(n_99),
.B(n_164),
.C(n_6),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_99),
.Y(n_334)
);


endmodule