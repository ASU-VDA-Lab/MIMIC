module fake_jpeg_9297_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_59),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_18),
.B1(n_29),
.B2(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_16),
.B1(n_20),
.B2(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_32),
.Y(n_63)
);

OAI21x1_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_30),
.B(n_28),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_40),
.C(n_23),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_86),
.C(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_84),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_81),
.B(n_19),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_88),
.B1(n_61),
.B2(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_79),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_108),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_110),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_107),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_76),
.C(n_64),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_28),
.B(n_21),
.C(n_60),
.D(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_40),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_72),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_102),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_45),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_120),
.B(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_124),
.C(n_128),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_119),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_2),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_43),
.B(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_126),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_56),
.B(n_43),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_128),
.B(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_58),
.B1(n_72),
.B2(n_85),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_106),
.B1(n_91),
.B2(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_56),
.B(n_53),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_53),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_138),
.B(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_145),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_143),
.B(n_154),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_105),
.B1(n_98),
.B2(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_94),
.B1(n_111),
.B2(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_161),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_R g152 ( 
.A(n_115),
.B(n_92),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_117),
.A3(n_116),
.B1(n_134),
.B2(n_10),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_157),
.B1(n_167),
.B2(n_130),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_53),
.B(n_4),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_3),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_159),
.C(n_129),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_5),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_6),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_130),
.C(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_189),
.B(n_7),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_159),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_179),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_114),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_187),
.B1(n_172),
.B2(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_133),
.C(n_119),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_143),
.C(n_160),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_165),
.B1(n_162),
.B2(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_149),
.B1(n_153),
.B2(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_141),
.B(n_154),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_212),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_166),
.B1(n_148),
.B2(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_148),
.B1(n_116),
.B2(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_205),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_176),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_157),
.B1(n_117),
.B2(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_191),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_132),
.B1(n_131),
.B2(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_177),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_218),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_183),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_191),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_227),
.C(n_215),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_212),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_201),
.B1(n_198),
.B2(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_197),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_173),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_236),
.Y(n_244)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_242),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_214),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_196),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_169),
.B1(n_200),
.B2(n_194),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_169),
.B1(n_179),
.B2(n_9),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_226),
.B(n_224),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_7),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_222),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_246),
.B(n_252),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_236),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_216),
.B(n_221),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_255),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_242),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_10),
.B(n_11),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_241),
.C(n_229),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_261),
.B(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_259),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_8),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_10),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_256),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_265),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_15),
.B(n_13),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_253),
.B1(n_255),
.B2(n_14),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_12),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_270),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_12),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_14),
.C(n_15),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_269),
.B1(n_263),
.B2(n_273),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_15),
.Y(n_277)
);


endmodule