module fake_jpeg_3521_n_218 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_218);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_62),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_79),
.B1(n_67),
.B2(n_68),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_79),
.B1(n_67),
.B2(n_68),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_55),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_70),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_74),
.B1(n_73),
.B2(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_61),
.B1(n_71),
.B2(n_70),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_81),
.B1(n_82),
.B2(n_93),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_84),
.Y(n_103)
);

OAI221xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_112),
.B1(n_116),
.B2(n_0),
.C(n_3),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_72),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_81),
.B1(n_83),
.B2(n_58),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_63),
.B(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR4xp25_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_28),
.C(n_51),
.D(n_48),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_83),
.B1(n_58),
.B2(n_62),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_110),
.B1(n_56),
.B2(n_5),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_63),
.B1(n_96),
.B2(n_76),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_101),
.Y(n_147)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_45),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_77),
.B1(n_64),
.B2(n_60),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_131),
.B1(n_139),
.B2(n_110),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_77),
.B1(n_57),
.B2(n_54),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_140),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_56),
.C(n_47),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_8),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_152),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_163),
.B1(n_122),
.B2(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_156),
.B(n_157),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_46),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_153),
.B(n_13),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_0),
.B(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_6),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

OR2x6_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_44),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_164),
.B(n_138),
.Y(n_171)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_6),
.CON(n_160),
.SN(n_160)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_14),
.C(n_15),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_171),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_138),
.B(n_21),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_175),
.B1(n_160),
.B2(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_23),
.B(n_40),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_182),
.B(n_165),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_22),
.B(n_38),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_162),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_144),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_166),
.A3(n_179),
.B1(n_169),
.B2(n_174),
.C1(n_181),
.C2(n_168),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_191),
.A3(n_188),
.B1(n_185),
.B2(n_16),
.C1(n_19),
.C2(n_18),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_182),
.B1(n_180),
.B2(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_198),
.B1(n_201),
.B2(n_18),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_172),
.B1(n_183),
.B2(n_17),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_207),
.B1(n_202),
.B2(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_27),
.C(n_34),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_210),
.B(n_206),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_209),
.B(n_196),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_207),
.C(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_201),
.B1(n_204),
.B2(n_35),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_43),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_205),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_217),
.Y(n_218)
);


endmodule