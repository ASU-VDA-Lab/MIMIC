module fake_jpeg_15677_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_72),
.Y(n_108)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_61),
.Y(n_110)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_51),
.B1(n_76),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_76),
.B1(n_70),
.B2(n_65),
.Y(n_119)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_55),
.B(n_71),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_102),
.B(n_58),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_74),
.B(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_59),
.B1(n_77),
.B2(n_63),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_119),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_59),
.B1(n_56),
.B2(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_68),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_61),
.B1(n_77),
.B2(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_2),
.Y(n_130)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_130),
.B(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_2),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_116),
.B(n_115),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_139),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_132),
.B(n_129),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_131),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_147),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_114),
.B1(n_124),
.B2(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_127),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_147),
.B1(n_34),
.B2(n_36),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_30),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_155),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_158),
.C(n_157),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_29),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_37),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_28),
.B(n_47),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_23),
.B1(n_49),
.B2(n_48),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_21),
.B(n_46),
.C(n_43),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_18),
.B(n_20),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_17),
.A3(n_42),
.B1(n_41),
.B2(n_38),
.C1(n_7),
.C2(n_14),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_16),
.B(n_120),
.Y(n_174)
);


endmodule