module real_aes_8149_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g492 ( .A(n_1), .Y(n_492) );
INVx1_ASAP7_75t_L g263 ( .A(n_2), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_3), .A2(n_36), .B1(n_182), .B2(n_520), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g170 ( .A1(n_4), .A2(n_171), .B(n_172), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_5), .B(n_169), .Y(n_469) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_239), .B(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_37), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g179 ( .A(n_9), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_10), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
INVx1_ASAP7_75t_L g488 ( .A(n_12), .Y(n_488) );
INVx1_ASAP7_75t_L g245 ( .A(n_13), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_14), .B(n_147), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_15), .B(n_137), .Y(n_497) );
AO32x2_ASAP7_75t_L g517 ( .A1(n_16), .A2(n_136), .A3(n_169), .B1(n_480), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_17), .B(n_182), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_18), .B(n_190), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_19), .B(n_137), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_20), .A2(n_49), .B1(n_182), .B2(n_520), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_21), .B(n_171), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_22), .A2(n_74), .B1(n_147), .B2(n_182), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_23), .B(n_182), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_24), .B(n_167), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_25), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_26), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_27), .B(n_184), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_28), .B(n_177), .Y(n_264) );
INVx1_ASAP7_75t_L g155 ( .A(n_29), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_30), .B(n_184), .Y(n_514) );
INVx2_ASAP7_75t_L g149 ( .A(n_31), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_32), .B(n_182), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_33), .B(n_184), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_34), .A2(n_41), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_34), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_35), .A2(n_144), .B(n_156), .C(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g153 ( .A(n_38), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_39), .A2(n_102), .B1(n_111), .B2(n_745), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_40), .B(n_177), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_41), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_42), .B(n_182), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_43), .A2(n_87), .B1(n_207), .B2(n_520), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_44), .B(n_182), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_45), .B(n_182), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_46), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_47), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_48), .B(n_171), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_50), .A2(n_59), .B1(n_147), .B2(n_182), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_51), .A2(n_147), .B1(n_150), .B2(n_156), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_52), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_53), .B(n_182), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_54), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_55), .B(n_182), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_56), .A2(n_176), .B(n_178), .C(n_181), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_57), .Y(n_220) );
INVx1_ASAP7_75t_L g173 ( .A(n_58), .Y(n_173) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_61), .B(n_182), .Y(n_493) );
INVx1_ASAP7_75t_L g140 ( .A(n_62), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_63), .Y(n_116) );
AO32x2_ASAP7_75t_L g537 ( .A1(n_64), .A2(n_169), .A3(n_225), .B1(n_480), .B2(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g477 ( .A(n_65), .Y(n_477) );
INVx1_ASAP7_75t_L g509 ( .A(n_66), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_SL g189 ( .A1(n_67), .A2(n_181), .B(n_190), .C(n_191), .Y(n_189) );
INVxp67_ASAP7_75t_L g192 ( .A(n_68), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_69), .B(n_147), .Y(n_510) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_71), .Y(n_164) );
INVx1_ASAP7_75t_L g213 ( .A(n_72), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_73), .A2(n_99), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_73), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_75), .A2(n_144), .B(n_156), .C(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_76), .B(n_520), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_77), .B(n_147), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_78), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_80), .B(n_190), .Y(n_204) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_81), .A2(n_447), .B1(n_735), .B2(n_738), .C1(n_739), .C2(n_741), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_82), .B(n_147), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_83), .A2(n_144), .B(n_156), .C(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g107 ( .A(n_84), .Y(n_107) );
OR2x2_ASAP7_75t_L g119 ( .A(n_84), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g450 ( .A(n_84), .B(n_121), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_85), .B(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_86), .A2(n_100), .B1(n_147), .B2(n_148), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_89), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_90), .A2(n_144), .B(n_156), .C(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_91), .Y(n_235) );
INVx1_ASAP7_75t_L g188 ( .A(n_92), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_93), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_94), .B(n_203), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_95), .B(n_147), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_96), .B(n_169), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_98), .A2(n_171), .B(n_187), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g737 ( .A(n_99), .Y(n_737) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g746 ( .A(n_103), .Y(n_746) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g734 ( .A(n_107), .B(n_121), .Y(n_734) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_107), .B(n_120), .Y(n_743) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_445), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g744 ( .A(n_116), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_442), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g444 ( .A(n_119), .Y(n_444) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_441), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g441 ( .A(n_129), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_129), .A2(n_448), .B1(n_451), .B2(n_732), .Y(n_447) );
AND3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_366), .C(n_415), .Y(n_129) );
NOR3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_273), .C(n_311), .Y(n_130) );
OAI222xp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_194), .B1(n_248), .B2(n_254), .C1(n_268), .C2(n_271), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_165), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_133), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_133), .B(n_316), .Y(n_407) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g284 ( .A(n_134), .B(n_185), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_134), .B(n_166), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_134), .B(n_304), .Y(n_327) );
OR2x2_ASAP7_75t_L g351 ( .A(n_134), .B(n_166), .Y(n_351) );
OR2x2_ASAP7_75t_L g359 ( .A(n_134), .B(n_258), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_134), .B(n_185), .Y(n_362) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g256 ( .A(n_135), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g270 ( .A(n_135), .B(n_185), .Y(n_270) );
AND2x2_ASAP7_75t_L g320 ( .A(n_135), .B(n_258), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_135), .B(n_166), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_135), .B(n_419), .Y(n_440) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_163), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_136), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_136), .A2(n_259), .B(n_266), .Y(n_258) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_138), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI22xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B1(n_159), .B2(n_160), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_143), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_143), .A2(n_174), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_143), .A2(n_174), .B(n_241), .C(n_242), .Y(n_240) );
INVx4_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g160 ( .A(n_144), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g171 ( .A(n_144), .B(n_161), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_144), .A2(n_461), .B(n_464), .Y(n_460) );
BUFx3_ASAP7_75t_L g480 ( .A(n_144), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_144), .A2(n_487), .B(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_144), .A2(n_508), .B(n_511), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_144), .A2(n_524), .B(n_528), .Y(n_523) );
INVx2_ASAP7_75t_L g265 ( .A(n_147), .Y(n_265) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx1_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_150) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx4_ASAP7_75t_L g243 ( .A(n_151), .Y(n_243) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
AND2x2_ASAP7_75t_L g161 ( .A(n_152), .B(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx3_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx5_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
BUFx3_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
INVx1_ASAP7_75t_L g520 ( .A(n_157), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_160), .A2(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g467 ( .A(n_162), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_165), .A2(n_359), .B(n_360), .C(n_363), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_165), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_165), .B(n_303), .Y(n_425) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_185), .Y(n_165) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_166), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g283 ( .A(n_166), .Y(n_283) );
AND2x2_ASAP7_75t_L g310 ( .A(n_166), .B(n_304), .Y(n_310) );
INVx1_ASAP7_75t_SL g318 ( .A(n_166), .Y(n_318) );
AND2x2_ASAP7_75t_L g341 ( .A(n_166), .B(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g419 ( .A(n_166), .Y(n_419) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_183), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g209 ( .A(n_168), .B(n_210), .Y(n_209) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_168), .B(n_480), .C(n_499), .Y(n_498) );
AO21x1_ASAP7_75t_L g543 ( .A1(n_168), .A2(n_499), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_169), .A2(n_186), .B(n_193), .Y(n_185) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_169), .A2(n_460), .B(n_469), .Y(n_459) );
BUFx2_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
O2A1O1Ixp5_ASAP7_75t_L g476 ( .A1(n_176), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_176), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_177), .A2(n_468), .B1(n_500), .B2(n_501), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_177), .A2(n_468), .B1(n_519), .B2(n_521), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_177), .A2(n_180), .B1(n_539), .B2(n_540), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_180), .B(n_192), .Y(n_191) );
INVx5_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
O2A1O1Ixp5_ASAP7_75t_SL g508 ( .A1(n_181), .A2(n_203), .B(n_509), .C(n_510), .Y(n_508) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
INVx2_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_184), .A2(n_238), .B(n_247), .Y(n_237) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_184), .A2(n_507), .B(n_514), .Y(n_506) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_184), .A2(n_523), .B(n_531), .Y(n_522) );
BUFx2_ASAP7_75t_L g255 ( .A(n_185), .Y(n_255) );
INVx1_ASAP7_75t_L g317 ( .A(n_185), .Y(n_317) );
INVx3_ASAP7_75t_L g342 ( .A(n_185), .Y(n_342) );
INVx1_ASAP7_75t_L g527 ( .A(n_190), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_194), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_222), .Y(n_194) );
INVx1_ASAP7_75t_L g338 ( .A(n_195), .Y(n_338) );
OAI32xp33_ASAP7_75t_L g344 ( .A1(n_195), .A2(n_283), .A3(n_345), .B1(n_346), .B2(n_347), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_195), .A2(n_349), .B1(n_352), .B2(n_357), .Y(n_348) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g286 ( .A(n_196), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g364 ( .A(n_196), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g434 ( .A(n_196), .B(n_380), .Y(n_434) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
AND2x2_ASAP7_75t_L g249 ( .A(n_197), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
INVx1_ASAP7_75t_L g298 ( .A(n_197), .Y(n_298) );
OR2x2_ASAP7_75t_L g306 ( .A(n_197), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g313 ( .A(n_197), .B(n_287), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_197), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_197), .B(n_252), .Y(n_334) );
INVx3_ASAP7_75t_L g356 ( .A(n_197), .Y(n_356) );
AND2x2_ASAP7_75t_L g381 ( .A(n_197), .B(n_253), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_197), .B(n_346), .Y(n_429) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
AOI21xp5_ASAP7_75t_SL g198 ( .A1(n_199), .A2(n_200), .B(n_208), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_205), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_203), .A2(n_263), .B(n_264), .C(n_265), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_203), .A2(n_462), .B(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g468 ( .A(n_203), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_203), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_205), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g218 ( .A(n_208), .Y(n_218) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_208), .A2(n_472), .B(n_481), .Y(n_471) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_208), .A2(n_486), .B(n_494), .Y(n_485) );
INVx2_ASAP7_75t_L g253 ( .A(n_211), .Y(n_253) );
AND2x2_ASAP7_75t_L g385 ( .A(n_211), .B(n_223), .Y(n_385) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_221), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_221), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g427 ( .A(n_222), .Y(n_427) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
AND2x2_ASAP7_75t_L g299 ( .A(n_223), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_223), .B(n_253), .Y(n_307) );
AND2x2_ASAP7_75t_L g365 ( .A(n_223), .B(n_288), .Y(n_365) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
AND2x2_ASAP7_75t_L g278 ( .A(n_224), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_224), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_224), .B(n_253), .Y(n_353) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_232), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_236), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_236), .B(n_253), .Y(n_346) );
AND2x2_ASAP7_75t_L g355 ( .A(n_236), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g380 ( .A(n_236), .Y(n_380) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g288 ( .A(n_237), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_243), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g490 ( .A(n_243), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_243), .A2(n_512), .B(n_513), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_248), .A2(n_258), .B1(n_417), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_250), .A2(n_361), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_251), .B(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g398 ( .A(n_251), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_252), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g325 ( .A(n_252), .B(n_278), .Y(n_325) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
INVx1_ASAP7_75t_L g331 ( .A(n_253), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_406), .B1(n_423), .B2(n_426), .C(n_428), .Y(n_422) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g293 ( .A(n_255), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_255), .B(n_304), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_256), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g347 ( .A(n_256), .B(n_293), .Y(n_347) );
INVx3_ASAP7_75t_SL g388 ( .A(n_256), .Y(n_388) );
AND2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_257), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_257), .B(n_270), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_257), .B(n_316), .Y(n_402) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
OAI322xp33_ASAP7_75t_L g399 ( .A1(n_258), .A2(n_330), .A3(n_352), .B1(n_400), .B2(n_402), .C1(n_403), .C2(n_404), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_265), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_269), .A2(n_272), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_270), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g371 ( .A(n_270), .B(n_283), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_270), .B(n_310), .Y(n_386) );
INVxp67_ASAP7_75t_L g337 ( .A(n_272), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_272), .A2(n_344), .B(n_348), .C(n_358), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_282), .B1(n_285), .B2(n_289), .C(n_294), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g297 ( .A(n_281), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g414 ( .A(n_281), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_282), .A2(n_431), .B1(n_436), .B2(n_437), .C(n_439), .Y(n_430) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_283), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g330 ( .A(n_283), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_283), .B(n_361), .Y(n_368) );
AND2x2_ASAP7_75t_L g410 ( .A(n_283), .B(n_388), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_284), .A2(n_296), .B1(n_406), .B2(n_407), .Y(n_405) );
OR2x2_ASAP7_75t_L g436 ( .A(n_284), .B(n_304), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g413 ( .A(n_287), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_287), .B(n_381), .Y(n_438) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_292), .B(n_303), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_301), .B1(n_305), .B2(n_308), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g369 ( .A(n_297), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_297), .B(n_337), .Y(n_404) );
AOI322xp5_ASAP7_75t_L g328 ( .A1(n_299), .A2(n_329), .A3(n_331), .B1(n_332), .B2(n_334), .C1(n_335), .C2(n_339), .Y(n_328) );
INVxp67_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_302), .A2(n_307), .B1(n_324), .B2(n_326), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_303), .B(n_316), .Y(n_403) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_304), .B(n_342), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_304), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g400 ( .A(n_306), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND3xp33_ASAP7_75t_SL g311 ( .A(n_312), .B(n_328), .C(n_343), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_319), .B2(n_321), .C(n_323), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_315), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g329 ( .A(n_320), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_322), .Y(n_401) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_327), .B(n_341), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_330), .B(n_388), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_331), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g406 ( .A(n_334), .Y(n_406) );
AND2x2_ASAP7_75t_L g421 ( .A(n_334), .B(n_398), .Y(n_421) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_345), .A2(n_416), .B(n_422), .C(n_430), .Y(n_415) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g384 ( .A(n_355), .B(n_385), .Y(n_384) );
NAND2x1_ASAP7_75t_SL g426 ( .A(n_356), .B(n_427), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_359), .Y(n_396) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
AND2x2_ASAP7_75t_L g395 ( .A(n_365), .B(n_381), .Y(n_395) );
NOR5xp2_ASAP7_75t_L g366 ( .A(n_367), .B(n_382), .C(n_399), .D(n_405), .E(n_408), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B1(n_370), .B2(n_372), .C(n_374), .Y(n_367) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_371), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g397 ( .A(n_381), .B(n_398), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_386), .B1(n_387), .B2(n_389), .C(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B1(n_396), .B2(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
AOI211xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_411), .B(n_413), .C(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_441), .A2(n_448), .B1(n_452), .B2(n_740), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_442), .B(n_446), .C(n_744), .Y(n_445) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_656), .Y(n_452) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_454), .B(n_614), .Y(n_453) );
NOR4xp25_ASAP7_75t_L g454 ( .A(n_455), .B(n_554), .C(n_590), .D(n_604), .Y(n_454) );
OAI221xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_502), .B1(n_532), .B2(n_541), .C(n_545), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_456), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_482), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
AND2x2_ASAP7_75t_L g551 ( .A(n_459), .B(n_471), .Y(n_551) );
INVx3_ASAP7_75t_L g559 ( .A(n_459), .Y(n_559) );
AND2x2_ASAP7_75t_L g613 ( .A(n_459), .B(n_485), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_459), .B(n_484), .Y(n_649) );
AND2x2_ASAP7_75t_L g707 ( .A(n_459), .B(n_569), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_468), .Y(n_464) );
INVx2_ASAP7_75t_L g478 ( .A(n_467), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_468), .A2(n_478), .B(n_492), .C(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g542 ( .A(n_470), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g556 ( .A(n_470), .B(n_485), .Y(n_556) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_471), .B(n_485), .Y(n_571) );
AND2x2_ASAP7_75t_L g583 ( .A(n_471), .B(n_559), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_471), .B(n_543), .Y(n_585) );
AND2x2_ASAP7_75t_L g620 ( .A(n_471), .B(n_543), .Y(n_620) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_471), .Y(n_665) );
INVx1_ASAP7_75t_L g673 ( .A(n_471), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_476), .B(n_480), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_482), .A2(n_591), .B1(n_595), .B2(n_599), .C(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g550 ( .A(n_483), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_495), .Y(n_483) );
INVx2_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
AND2x2_ASAP7_75t_L g602 ( .A(n_484), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g621 ( .A(n_484), .B(n_559), .Y(n_621) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g684 ( .A(n_485), .B(n_559), .Y(n_684) );
AND2x2_ASAP7_75t_L g606 ( .A(n_495), .B(n_551), .Y(n_606) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_495), .A2(n_630), .A3(n_675), .B1(n_677), .B2(n_680), .C1(n_682), .C2(n_686), .Y(n_674) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_496), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
AND2x2_ASAP7_75t_L g679 ( .A(n_496), .B(n_559), .Y(n_679) );
AND2x2_ASAP7_75t_L g711 ( .A(n_496), .B(n_583), .Y(n_711) );
OR2x2_ASAP7_75t_L g714 ( .A(n_496), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g544 ( .A(n_497), .Y(n_544) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
INVx1_ASAP7_75t_L g727 ( .A(n_504), .Y(n_727) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g534 ( .A(n_505), .B(n_522), .Y(n_534) );
INVx2_ASAP7_75t_L g567 ( .A(n_505), .Y(n_567) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g589 ( .A(n_506), .Y(n_589) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_506), .Y(n_597) );
OR2x2_ASAP7_75t_L g721 ( .A(n_506), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g638 ( .A(n_515), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
AND2x2_ASAP7_75t_L g535 ( .A(n_516), .B(n_536), .Y(n_535) );
NOR2xp67_ASAP7_75t_L g593 ( .A(n_516), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g647 ( .A(n_516), .B(n_537), .Y(n_647) );
OR2x2_ASAP7_75t_L g655 ( .A(n_516), .B(n_589), .Y(n_655) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_517), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g598 ( .A(n_517), .B(n_522), .Y(n_598) );
AND2x2_ASAP7_75t_L g662 ( .A(n_517), .B(n_537), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_522), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g575 ( .A(n_522), .Y(n_575) );
INVx1_ASAP7_75t_L g580 ( .A(n_522), .Y(n_580) );
AND2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_522), .Y(n_670) );
INVx1_ASAP7_75t_L g722 ( .A(n_522), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_527), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g699 ( .A(n_533), .B(n_608), .Y(n_699) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g626 ( .A(n_535), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g725 ( .A(n_535), .B(n_660), .Y(n_725) );
INVx1_ASAP7_75t_L g547 ( .A(n_536), .Y(n_547) );
AND2x2_ASAP7_75t_L g573 ( .A(n_536), .B(n_567), .Y(n_573) );
BUFx2_ASAP7_75t_L g632 ( .A(n_536), .Y(n_632) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_537), .Y(n_553) );
INVx1_ASAP7_75t_L g563 ( .A(n_537), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g701 ( .A(n_541), .B(n_548), .Y(n_701) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI32xp33_ASAP7_75t_L g545 ( .A1(n_542), .A2(n_546), .A3(n_548), .B1(n_550), .B2(n_552), .Y(n_545) );
AND2x2_ASAP7_75t_L g685 ( .A(n_542), .B(n_558), .Y(n_685) );
AND2x2_ASAP7_75t_L g723 ( .A(n_542), .B(n_621), .Y(n_723) );
INVx1_ASAP7_75t_L g603 ( .A(n_543), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_547), .B(n_609), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_548), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_548), .B(n_551), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_548), .B(n_620), .Y(n_702) );
OR2x2_ASAP7_75t_L g716 ( .A(n_548), .B(n_585), .Y(n_716) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g643 ( .A(n_549), .B(n_551), .Y(n_643) );
OR2x2_ASAP7_75t_L g652 ( .A(n_549), .B(n_639), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_551), .B(n_602), .Y(n_624) );
INVx2_ASAP7_75t_L g639 ( .A(n_553), .Y(n_639) );
OR2x2_ASAP7_75t_L g654 ( .A(n_553), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_553), .B(n_670), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_553), .A2(n_646), .B(n_727), .C(n_728), .Y(n_726) );
OAI321xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_560), .A3(n_565), .B1(n_568), .B2(n_572), .C(n_576), .Y(n_554) );
INVx1_ASAP7_75t_L g667 ( .A(n_555), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g678 ( .A(n_556), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g630 ( .A(n_558), .Y(n_630) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_559), .B(n_673), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_560), .A2(n_698), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_697) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AND2x2_ASAP7_75t_L g635 ( .A(n_562), .B(n_609), .Y(n_635) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_563), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g608 ( .A(n_564), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_565), .A2(n_606), .B(n_651), .C(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g617 ( .A(n_567), .B(n_574), .Y(n_617) );
BUFx2_ASAP7_75t_L g627 ( .A(n_567), .Y(n_627) );
INVx1_ASAP7_75t_L g642 ( .A(n_567), .Y(n_642) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OR2x2_ASAP7_75t_L g648 ( .A(n_570), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g731 ( .A(n_570), .Y(n_731) );
INVx1_ASAP7_75t_L g724 ( .A(n_571), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g577 ( .A(n_573), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g681 ( .A(n_573), .B(n_598), .Y(n_681) );
INVx1_ASAP7_75t_L g610 ( .A(n_574), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B1(n_584), .B2(n_586), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_578), .B(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g646 ( .A(n_579), .B(n_647), .Y(n_646) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_580), .B(n_589), .Y(n_609) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g601 ( .A(n_583), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g611 ( .A(n_585), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_588), .A2(n_706), .B1(n_708), .B2(n_709), .C(n_710), .Y(n_705) );
INVx1_ASAP7_75t_L g594 ( .A(n_589), .Y(n_594) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_589), .Y(n_660) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_592), .B(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_593), .A2(n_598), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_596), .B(n_606), .Y(n_703) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g672 ( .A(n_597), .Y(n_672) );
AND2x2_ASAP7_75t_L g631 ( .A(n_598), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g720 ( .A(n_598), .Y(n_720) );
INVx1_ASAP7_75t_L g636 ( .A(n_601), .Y(n_636) );
INVx1_ASAP7_75t_L g691 ( .A(n_602), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B1(n_610), .B2(n_611), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_608), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g676 ( .A(n_609), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_609), .B(n_647), .Y(n_713) );
OR2x2_ASAP7_75t_L g686 ( .A(n_610), .B(n_639), .Y(n_686) );
INVx1_ASAP7_75t_L g625 ( .A(n_611), .Y(n_625) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_613), .B(n_664), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_633), .C(n_644), .Y(n_614) );
OAI211xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_622), .C(n_628), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_617), .A2(n_688), .B1(n_692), .B2(n_695), .C(n_697), .Y(n_687) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g629 ( .A(n_620), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g683 ( .A(n_620), .B(n_684), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_621), .A2(n_669), .B(n_671), .C(n_673), .Y(n_668) );
INVx2_ASAP7_75t_L g715 ( .A(n_621), .Y(n_715) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_625), .B(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g694 ( .A(n_627), .B(n_647), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_636), .B(n_637), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_643), .B(n_730), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B(n_650), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g671 ( .A(n_647), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND4x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_687), .C(n_704), .D(n_726), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_674), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_663), .B(n_666), .C(n_668), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_662), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_673), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g708 ( .A(n_683), .Y(n_708) );
INVx2_ASAP7_75t_SL g696 ( .A(n_684), .Y(n_696) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g709 ( .A(n_694), .Y(n_709) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_712), .Y(n_704) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B1(n_716), .B2(n_717), .C(n_718), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g740 ( .A(n_733), .Y(n_740) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_735), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
endmodule