module fake_jpeg_4678_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_29),
.Y(n_49)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_26),
.B1(n_19),
.B2(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_26),
.B1(n_19),
.B2(n_15),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_57),
.B1(n_61),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_65),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_31),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_36),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_17),
.B(n_28),
.C(n_32),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_41),
.B(n_23),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_41),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_81),
.B1(n_53),
.B2(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_83),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_35),
.C(n_32),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_22),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_46),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_58),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_34),
.B1(n_19),
.B2(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_89),
.B1(n_104),
.B2(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_59),
.B1(n_50),
.B2(n_64),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_50),
.A3(n_65),
.B1(n_35),
.B2(n_37),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_32),
.B(n_53),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_99),
.B(n_78),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_58),
.B1(n_42),
.B2(n_68),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_54),
.B1(n_34),
.B2(n_43),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_68),
.B1(n_81),
.B2(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_58),
.B1(n_42),
.B2(n_60),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_69),
.A3(n_75),
.B1(n_74),
.B2(n_78),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_118),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_103),
.B(n_76),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_119),
.B1(n_73),
.B2(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_71),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_81),
.C(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_134),
.C(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_138),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_92),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_132),
.B(n_135),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_88),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_76),
.B(n_67),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_106),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_73),
.B1(n_99),
.B2(n_100),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_125),
.B1(n_108),
.B2(n_114),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_121),
.B1(n_112),
.B2(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_73),
.B(n_95),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_107),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_115),
.CI(n_119),
.CON(n_169),
.SN(n_169)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_151),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_113),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_166),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_117),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_150),
.B1(n_169),
.B2(n_146),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_117),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_165),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_111),
.B1(n_87),
.B2(n_84),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_145),
.B1(n_127),
.B2(n_138),
.Y(n_176)
);

NOR2x1_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_130),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_175),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_134),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_188),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_177),
.B1(n_18),
.B2(n_25),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_129),
.B1(n_127),
.B2(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_87),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_156),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_28),
.B1(n_20),
.B2(n_23),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_35),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_77),
.B1(n_34),
.B2(n_25),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_24),
.C(n_13),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_56),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_170),
.C(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_199),
.C(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_161),
.C(n_169),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_56),
.C(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_40),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_206),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_21),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_178),
.B(n_25),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_40),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_35),
.C(n_40),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_184),
.C(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_182),
.B1(n_180),
.B2(n_173),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_210),
.B1(n_207),
.B2(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_216),
.C(n_219),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_172),
.C(n_187),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_224),
.B(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_188),
.C(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_21),
.B1(n_16),
.B2(n_24),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_24),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_219),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_13),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_21),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_0),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_239),
.B1(n_214),
.B2(n_1),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_212),
.C(n_209),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_234),
.C(n_242),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_201),
.C(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_0),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_13),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_6),
.B(n_1),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_6),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_217),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_0),
.C(n_1),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_254),
.C(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_3),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_253),
.B(n_4),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_3),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_3),
.C(n_4),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_256),
.B(n_259),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_228),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_264),
.B(n_7),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_233),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_270),
.B(n_271),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_256),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_268),
.B(n_8),
.Y(n_274)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_252),
.B(n_251),
.C(n_254),
.D(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_8),
.C(n_9),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_7),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_12),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_8),
.B(n_9),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_274),
.B(n_10),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_8),
.C(n_9),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_10),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_11),
.B(n_12),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_278),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_11),
.Y(n_284)
);


endmodule