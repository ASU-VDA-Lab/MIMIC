module fake_jpeg_714_n_234 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_234);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx10_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_34),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_72),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_84),
.B1(n_81),
.B2(n_78),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_84),
.B1(n_81),
.B2(n_58),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_59),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_68),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_74),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_64),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_116),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_65),
.C(n_55),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_115),
.C(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_71),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_63),
.B(n_75),
.C(n_66),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_64),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_137),
.B1(n_102),
.B2(n_99),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_73),
.C(n_60),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_141),
.Y(n_148)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_82),
.B(n_62),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_82),
.B(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_23),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_77),
.C(n_74),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_153),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_67),
.B(n_77),
.C(n_25),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_150),
.B(n_32),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_67),
.B1(n_24),
.B2(n_26),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_0),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_0),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_159),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_2),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_165),
.Y(n_166)
);

AO21x2_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_28),
.B(n_50),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_163),
.B1(n_131),
.B2(n_128),
.Y(n_170)
);

NAND2xp67_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_4),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_5),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_122),
.B1(n_131),
.B2(n_139),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_184),
.B1(n_22),
.B2(n_49),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_148),
.Y(n_169)
);

OAI31xp33_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_160),
.A3(n_163),
.B(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_29),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_177),
.Y(n_200)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_129),
.C(n_30),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_12),
.C(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_162),
.B1(n_150),
.B2(n_11),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_12),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_35),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_36),
.C(n_48),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_171),
.C(n_166),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_207),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_171),
.B(n_184),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_170),
.B1(n_168),
.B2(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_166),
.B1(n_185),
.B2(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_195),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_176),
.B1(n_37),
.B2(n_41),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_200),
.C(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_203),
.C(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_14),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_18),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_203),
.B1(n_18),
.B2(n_17),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_223),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_224),
.B1(n_215),
.B2(n_218),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_43),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_214),
.Y(n_227)
);

AOI31xp67_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_221),
.A3(n_217),
.B(n_223),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_217),
.B(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_20),
.B(n_21),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_33),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_45),
.B(n_46),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_47),
.Y(n_234)
);


endmodule