module fake_jpeg_19615_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_5),
.A2(n_6),
.B1(n_4),
.B2(n_1),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_0),
.B(n_2),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_22),
.B(n_10),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_2),
.B1(n_5),
.B2(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_12),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_21),
.B(n_11),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_15),
.A2(n_11),
.B1(n_14),
.B2(n_17),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_14),
.C(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_26),
.C(n_27),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_26),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_28),
.B(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_41)
);


endmodule