module fake_jpeg_903_n_650 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_3),
.B(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_61),
.Y(n_184)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_20),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g219 ( 
.A(n_63),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_75),
.Y(n_142)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g185 ( 
.A(n_66),
.Y(n_185)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_72),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_24),
.A2(n_19),
.B(n_18),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_56),
.B(n_55),
.Y(n_135)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_76),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_30),
.Y(n_77)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx2_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_87),
.Y(n_143)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_83),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_1),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_84),
.B(n_37),
.Y(n_178)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_30),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_88),
.Y(n_224)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_91),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_29),
.B(n_4),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_94),
.Y(n_223)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_100),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_33),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_29),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_115),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_110),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_35),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_23),
.B1(n_46),
.B2(n_48),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_38),
.B(n_18),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_36),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_122),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_36),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_5),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_38),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_39),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_130),
.Y(n_183)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_27),
.B1(n_42),
.B2(n_45),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_133),
.A2(n_141),
.B1(n_152),
.B2(n_155),
.Y(n_266)
);

OR2x2_ASAP7_75t_SL g237 ( 
.A(n_135),
.B(n_61),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_53),
.B1(n_47),
.B2(n_51),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_136),
.A2(n_167),
.B1(n_189),
.B2(n_191),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_78),
.B(n_39),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_151),
.B(n_160),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_27),
.B1(n_42),
.B2(n_45),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_50),
.B1(n_23),
.B2(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_156),
.B(n_112),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_50),
.B1(n_46),
.B2(n_53),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_157),
.A2(n_161),
.B1(n_163),
.B2(n_179),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_49),
.B1(n_47),
.B2(n_51),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_72),
.A2(n_56),
.B1(n_55),
.B2(n_26),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_84),
.A2(n_49),
.B1(n_37),
.B2(n_26),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_166),
.A2(n_181),
.B1(n_199),
.B2(n_88),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_84),
.A2(n_37),
.B1(n_26),
.B2(n_21),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_178),
.B(n_215),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_116),
.A2(n_21),
.B1(n_43),
.B2(n_25),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_62),
.A2(n_68),
.B1(n_64),
.B2(n_124),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_77),
.B(n_21),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_196),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_200),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_70),
.A2(n_54),
.B1(n_8),
.B2(n_9),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_197),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_85),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_89),
.B(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_193),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_81),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_63),
.B(n_10),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_129),
.A2(n_90),
.B1(n_123),
.B2(n_117),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_80),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_66),
.B(n_17),
.C(n_14),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_91),
.B(n_12),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_206),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_93),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_204),
.A2(n_217),
.B1(n_162),
.B2(n_172),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_205),
.A2(n_216),
.B1(n_220),
.B2(n_103),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_91),
.B(n_15),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_63),
.B(n_15),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_211),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_58),
.B(n_111),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_94),
.A2(n_99),
.B1(n_74),
.B2(n_125),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_95),
.A2(n_71),
.B1(n_96),
.B2(n_98),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_61),
.A2(n_98),
.B1(n_96),
.B2(n_83),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_101),
.B(n_107),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_61),
.B(n_101),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_69),
.B(n_76),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_112),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_142),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_229),
.B(n_237),
.C(n_245),
.Y(n_324)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_131),
.Y(n_231)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_232),
.B(n_250),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_234),
.Y(n_332)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_139),
.B(n_178),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_236),
.B(n_246),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_238),
.B(n_241),
.Y(n_358)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_239),
.Y(n_361)
);

HB1xp67_ASAP7_75t_SL g327 ( 
.A(n_240),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_134),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g243 ( 
.A(n_215),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g364 ( 
.A(n_243),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_143),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_178),
.B(n_107),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_253),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_254),
.A2(n_290),
.B1(n_313),
.B2(n_184),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_179),
.A2(n_163),
.B(n_194),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_255),
.A2(n_311),
.B(n_184),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_148),
.B(n_195),
.C(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_291),
.C(n_293),
.Y(n_343)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_258),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_158),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_263),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_260),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_193),
.B(n_211),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_261),
.Y(n_366)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_262),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_166),
.B(n_156),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_154),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_159),
.B(n_174),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_267),
.Y(n_360)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_170),
.B(n_171),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_131),
.Y(n_271)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_228),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_272),
.Y(n_329)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_273),
.Y(n_334)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_154),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_275),
.B(n_285),
.Y(n_348)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_277),
.Y(n_333)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_165),
.Y(n_278)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_279),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_136),
.B(n_167),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_287),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_185),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_281),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_144),
.A2(n_181),
.B1(n_175),
.B2(n_180),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_282),
.A2(n_304),
.B1(n_305),
.B2(n_310),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_309),
.B1(n_164),
.B2(n_218),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_185),
.B(n_215),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_284),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_176),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_286),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_169),
.B(n_177),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_183),
.B(n_189),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_299),
.Y(n_349)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_216),
.A2(n_199),
.B1(n_141),
.B2(n_190),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_180),
.C(n_183),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_150),
.B(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_297),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_198),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_150),
.B(n_225),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_303),
.C(n_285),
.Y(n_369)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_145),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_301),
.Y(n_359)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_145),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_306),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_198),
.B(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_147),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_138),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_207),
.B(n_147),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_182),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_176),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_308),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_149),
.A2(n_153),
.B1(n_212),
.B2(n_162),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_207),
.A2(n_202),
.B1(n_218),
.B2(n_168),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_138),
.A2(n_184),
.B(n_153),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_172),
.B1(n_202),
.B2(n_182),
.Y(n_325)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_168),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_244),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_325),
.A2(n_365),
.B1(n_309),
.B2(n_311),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_345),
.A2(n_351),
.B1(n_355),
.B2(n_370),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_288),
.A2(n_149),
.B1(n_212),
.B2(n_164),
.Y(n_355)
);

NAND2x1_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_303),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_SL g362 ( 
.A(n_259),
.B(n_227),
.C(n_261),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_237),
.C(n_246),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_263),
.A2(n_227),
.B1(n_280),
.B2(n_232),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_283),
.A2(n_268),
.B1(n_266),
.B2(n_296),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_244),
.A2(n_255),
.B(n_285),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_300),
.B(n_293),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_329),
.B(n_236),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_374),
.B(n_388),
.Y(n_456)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_378),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_370),
.A2(n_261),
.B1(n_252),
.B2(n_242),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_377),
.A2(n_386),
.B1(n_398),
.B2(n_409),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_395),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_364),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_380),
.B(n_391),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_256),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_381),
.Y(n_443)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_344),
.C(n_343),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_397),
.C(n_411),
.Y(n_422)
);

BUFx12_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_385),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_317),
.A2(n_252),
.B1(n_248),
.B2(n_307),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_326),
.B(n_292),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_251),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_403),
.B(n_419),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_291),
.B1(n_287),
.B2(n_230),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_394),
.B1(n_323),
.B2(n_340),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_317),
.A2(n_257),
.B1(n_305),
.B2(n_233),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_344),
.B(n_303),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_319),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_293),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_351),
.A2(n_301),
.B1(n_302),
.B2(n_271),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_400),
.B(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_368),
.B(n_262),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_405),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_403),
.A2(n_407),
.B(n_418),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_316),
.B(n_269),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_414),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_243),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_357),
.B(n_277),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_406),
.B(n_408),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_358),
.A2(n_234),
.B1(n_313),
.B2(n_300),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_341),
.B(n_273),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_349),
.A2(n_231),
.B1(n_235),
.B2(n_239),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_410),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_343),
.B(n_279),
.C(n_298),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_267),
.C(n_278),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_419),
.C(n_348),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_363),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_340),
.B(n_234),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_415),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_348),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_416),
.B(n_417),
.Y(n_449)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_327),
.A2(n_294),
.B1(n_299),
.B2(n_276),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_274),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_353),
.B(n_258),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_420),
.B(n_421),
.Y(n_458)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_321),
.Y(n_421)
);

AOI22x1_ASAP7_75t_L g425 ( 
.A1(n_412),
.A2(n_356),
.B1(n_349),
.B2(n_340),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_425),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_426),
.B(n_411),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_428),
.A2(n_430),
.B1(n_433),
.B2(n_377),
.Y(n_468)
);

OAI22x1_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_345),
.B1(n_234),
.B2(n_347),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_431),
.A2(n_439),
.B(n_447),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_393),
.A2(n_359),
.B1(n_324),
.B2(n_369),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_320),
.B1(n_338),
.B2(n_367),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_434),
.A2(n_342),
.B1(n_336),
.B2(n_371),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_333),
.C(n_354),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_440),
.C(n_413),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_350),
.B(n_332),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_334),
.C(n_319),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_400),
.A2(n_320),
.B1(n_367),
.B2(n_342),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_445),
.A2(n_379),
.B1(n_375),
.B2(n_382),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_392),
.A2(n_332),
.B(n_334),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_448),
.B(n_457),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_322),
.B(n_275),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_454),
.B(n_460),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_346),
.B(n_360),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_339),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_378),
.A2(n_339),
.B(n_337),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_414),
.A2(n_322),
.B(n_314),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_456),
.B(n_374),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_463),
.B(n_465),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_448),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_456),
.B(n_386),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_468),
.A2(n_474),
.B1(n_487),
.B2(n_492),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_394),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_469),
.B(n_475),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_496),
.B1(n_439),
.B2(n_430),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_398),
.B1(n_404),
.B2(n_397),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_427),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_459),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_477),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_438),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_490),
.C(n_495),
.Y(n_502)
);

OAI32xp33_ASAP7_75t_L g480 ( 
.A1(n_435),
.A2(n_389),
.A3(n_387),
.B1(n_417),
.B2(n_376),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_480),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_435),
.A2(n_396),
.B1(n_409),
.B2(n_391),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_481),
.A2(n_442),
.B1(n_260),
.B2(n_297),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_449),
.Y(n_482)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_482),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_421),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_483),
.Y(n_505)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_443),
.B(n_372),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_485),
.B(n_486),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_446),
.B(n_337),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_424),
.Y(n_488)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_488),
.Y(n_506)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_336),
.C(n_371),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_430),
.A2(n_410),
.B1(n_383),
.B2(n_314),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_360),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_499),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_361),
.Y(n_494)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_457),
.C(n_423),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_425),
.A2(n_295),
.B1(n_289),
.B2(n_321),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_434),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_497),
.B(n_498),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_449),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_361),
.C(n_330),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_426),
.C(n_436),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_468),
.A2(n_437),
.B1(n_431),
.B2(n_425),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_503),
.A2(n_519),
.B1(n_521),
.B2(n_479),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_471),
.A2(n_444),
.B(n_454),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_504),
.A2(n_483),
.B(n_496),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_472),
.A2(n_444),
.B(n_447),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_507),
.A2(n_470),
.B(n_471),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_508),
.A2(n_515),
.B1(n_534),
.B2(n_535),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_512),
.C(n_513),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_440),
.C(n_460),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_494),
.Y(n_514)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_499),
.C(n_467),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_428),
.B1(n_437),
.B2(n_433),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_453),
.C(n_461),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_517),
.C(n_530),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_453),
.C(n_461),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_458),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_491),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_479),
.A2(n_477),
.B1(n_474),
.B2(n_492),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_479),
.A2(n_458),
.B1(n_462),
.B2(n_445),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_464),
.B(n_455),
.C(n_451),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_472),
.A2(n_451),
.B(n_452),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_532),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_473),
.A2(n_452),
.B1(n_442),
.B2(n_321),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_501),
.B(n_488),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_SL g568 ( 
.A(n_536),
.B(n_548),
.C(n_557),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_529),
.B(n_465),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_537),
.B(n_543),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_538),
.A2(n_547),
.B(n_555),
.Y(n_577)
);

OAI21xp33_ASAP7_75t_L g539 ( 
.A1(n_516),
.A2(n_470),
.B(n_500),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_539),
.B(n_551),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_542),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_476),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_544),
.B(n_554),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_552),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_504),
.A2(n_483),
.B(n_498),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_501),
.Y(n_549)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_526),
.Y(n_550)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_550),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_482),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_520),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_502),
.B(n_481),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_533),
.A2(n_487),
.B1(n_480),
.B2(n_484),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_489),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_556),
.B(n_561),
.Y(n_584)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_510),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_505),
.B(n_466),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_558),
.B(n_559),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_531),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_512),
.B(n_330),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_528),
.A2(n_335),
.B1(n_385),
.B2(n_306),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_562),
.A2(n_563),
.B1(n_521),
.B2(n_510),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_531),
.B(n_506),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_533),
.B(n_507),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_565),
.A2(n_524),
.B(n_522),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_556),
.B(n_509),
.C(n_517),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_567),
.B(n_569),
.Y(n_598)
);

AO221x1_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_534),
.B1(n_508),
.B2(n_535),
.C(n_515),
.Y(n_569)
);

INVx13_ASAP7_75t_L g570 ( 
.A(n_552),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_570),
.B(n_574),
.Y(n_605)
);

BUFx12_ASAP7_75t_L g571 ( 
.A(n_547),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_571),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_575),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_538),
.B(n_545),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_576),
.A2(n_582),
.B(n_536),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_541),
.B(n_513),
.C(n_532),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_247),
.C(n_249),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_560),
.A2(n_503),
.B1(n_563),
.B2(n_558),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_580),
.A2(n_562),
.B1(n_520),
.B2(n_385),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_558),
.A2(n_506),
.B(n_527),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_544),
.B(n_518),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_541),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_587),
.B(n_593),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_582),
.Y(n_588)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_588),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_589),
.A2(n_592),
.B(n_594),
.Y(n_606)
);

A2O1A1O1Ixp25_ASAP7_75t_L g592 ( 
.A1(n_565),
.A2(n_511),
.B(n_553),
.C(n_555),
.D(n_523),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_561),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_576),
.A2(n_523),
.B(n_554),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_595),
.A2(n_599),
.B1(n_575),
.B2(n_579),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_553),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_596),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_597),
.A2(n_590),
.B1(n_605),
.B2(n_591),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_566),
.A2(n_335),
.B1(n_385),
.B2(n_264),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_601),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_585),
.B(n_573),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_603),
.Y(n_609)
);

OAI221xp5_ASAP7_75t_L g603 ( 
.A1(n_564),
.A2(n_574),
.B1(n_579),
.B2(n_567),
.C(n_566),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_572),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_577),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_581),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_584),
.C(n_583),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_608),
.B(n_616),
.Y(n_631)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_612),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_572),
.B1(n_580),
.B2(n_568),
.Y(n_614)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_614),
.Y(n_622)
);

OAI21x1_ASAP7_75t_SL g630 ( 
.A1(n_615),
.A2(n_620),
.B(n_619),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_598),
.B(n_584),
.C(n_583),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_586),
.C(n_569),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_617),
.B(n_587),
.Y(n_623)
);

OAI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_618),
.A2(n_619),
.B1(n_597),
.B2(n_607),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_589),
.A2(n_571),
.B1(n_581),
.B2(n_570),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_620),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_627),
.Y(n_635)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_625),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_609),
.A2(n_592),
.B1(n_571),
.B2(n_601),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_626),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_613),
.B(n_599),
.C(n_571),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_609),
.A2(n_570),
.B(n_606),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_628),
.A2(n_630),
.B(n_620),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_611),
.B(n_606),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_629),
.B(n_610),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_617),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_633),
.B(n_634),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_616),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_636),
.B(n_638),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g639 ( 
.A(n_622),
.B(n_608),
.Y(n_639)
);

AOI321xp33_ASAP7_75t_L g641 ( 
.A1(n_639),
.A2(n_626),
.A3(n_624),
.B1(n_627),
.B2(n_625),
.C(n_618),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_641),
.A2(n_643),
.B(n_635),
.Y(n_646)
);

BUFx24_ASAP7_75t_SL g642 ( 
.A(n_637),
.Y(n_642)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_642),
.Y(n_645)
);

BUFx24_ASAP7_75t_SL g643 ( 
.A(n_637),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_644),
.C(n_640),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_645),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_632),
.B(n_624),
.Y(n_650)
);


endmodule