module fake_jpeg_30093_n_64 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

INVx1_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

XNOR2x1_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_27),
.B1(n_24),
.B2(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_2),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_14),
.B(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_37),
.B1(n_8),
.B2(n_9),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_5),
.C(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_42),
.B1(n_11),
.B2(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_42),
.B1(n_13),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_22),
.B(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_53),
.C(n_59),
.Y(n_63)
);

NOR4xp25_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_56),
.C(n_20),
.D(n_61),
.Y(n_64)
);


endmodule