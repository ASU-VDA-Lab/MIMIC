module real_jpeg_28463_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_0),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_8),
.B1(n_22),
.B2(n_26),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_26),
.B1(n_45),
.B2(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_7),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_8),
.B1(n_22),
.B2(n_29),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_8),
.B(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_19),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_9),
.B(n_38),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_7),
.A2(n_42),
.B(n_46),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_7),
.B(n_51),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_9),
.B1(n_22),
.B2(n_52),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_29),
.B(n_114),
.C(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_108),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_106),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_82),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_15),
.B(n_82),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_60),
.C(n_72),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_16)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_33),
.C(n_49),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_27),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_19),
.A2(n_28),
.B1(n_30),
.B2(n_86),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_20),
.A2(n_25),
.B(n_29),
.C(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_29),
.A2(n_38),
.B(n_43),
.C(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_29),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_29),
.B(n_44),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_36),
.B(n_40),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_36),
.A2(n_40),
.B1(n_44),
.B2(n_98),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_45),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_96),
.C(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_48),
.A2(n_49),
.B1(n_95),
.B2(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_54),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_53),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_72),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_64),
.A2(n_65),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_129),
.C(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_71),
.B(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_88),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_76),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_96),
.B1(n_136),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_164),
.B(n_168),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_132),
.B(n_163),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_111),
.B(n_120),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_119),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_129),
.C(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_158),
.B(n_162),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_143),
.B(n_157),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B(n_156),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_153),
.B(n_155),
.Y(n_147)
);

INVx5_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.Y(n_168)
);


endmodule