module fake_jpeg_10868_n_367 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_367);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_367;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_48),
.Y(n_85)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_72),
.Y(n_96)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_55),
.Y(n_90)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_52),
.Y(n_88)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g107 ( 
.A(n_54),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_56),
.Y(n_121)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_11),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_27),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_38),
.B1(n_27),
.B2(n_14),
.Y(n_79)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

BUFx2_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_79),
.A2(n_82),
.B1(n_89),
.B2(n_94),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_83),
.B(n_103),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_24),
.B1(n_29),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_106),
.B1(n_117),
.B2(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_104),
.B(n_87),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_38),
.B1(n_21),
.B2(n_14),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_41),
.A2(n_21),
.B1(n_14),
.B2(n_38),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_56),
.B1(n_63),
.B2(n_65),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_64),
.B1(n_51),
.B2(n_47),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_19),
.B1(n_36),
.B2(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_62),
.B1(n_71),
.B2(n_44),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_124),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_45),
.A2(n_21),
.B1(n_31),
.B2(n_29),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_127),
.B1(n_69),
.B2(n_68),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_39),
.B1(n_28),
.B2(n_26),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_58),
.A2(n_39),
.B1(n_28),
.B2(n_26),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_128),
.B(n_135),
.Y(n_206)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_54),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_4),
.Y(n_135)
);

NAND2x1p5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_74),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_139),
.B(n_143),
.Y(n_176)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_154),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_140),
.B(n_142),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_65),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_68),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_161),
.B1(n_154),
.B2(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_100),
.B1(n_120),
.B2(n_102),
.Y(n_183)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_10),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_10),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_108),
.A2(n_80),
.B1(n_119),
.B2(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_93),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_165),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_78),
.B1(n_92),
.B2(n_100),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_105),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_89),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_87),
.B(n_92),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_102),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_180),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_117),
.B1(n_78),
.B2(n_99),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_179),
.A2(n_183),
.B1(n_130),
.B2(n_152),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_111),
.C(n_107),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_111),
.C(n_97),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_184),
.B(n_150),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_133),
.B(n_114),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_196),
.B(n_205),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_126),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_159),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_134),
.B(n_145),
.C(n_162),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_203),
.A2(n_190),
.B(n_183),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_143),
.B(n_112),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_172),
.B1(n_131),
.B2(n_120),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_174),
.B1(n_146),
.B2(n_137),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_112),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_167),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_138),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_222),
.Y(n_266)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_229),
.Y(n_261)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_167),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_226),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_159),
.B1(n_171),
.B2(n_166),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_213),
.B1(n_204),
.B2(n_200),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_236),
.B(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_237),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_129),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_235),
.B(n_212),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_176),
.A2(n_155),
.B1(n_156),
.B2(n_126),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_191),
.A2(n_164),
.B1(n_151),
.B2(n_132),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_247),
.B(n_248),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_146),
.B1(n_151),
.B2(n_188),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_206),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_191),
.B1(n_190),
.B2(n_205),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_179),
.B1(n_189),
.B2(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_184),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_187),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_186),
.B(n_178),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_197),
.C(n_186),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_178),
.C(n_204),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_260),
.B(n_232),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_210),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_264),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_210),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_274),
.B1(n_265),
.B2(n_261),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_182),
.B(n_213),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_260),
.B(n_259),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_227),
.A2(n_182),
.B1(n_236),
.B2(n_240),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_240),
.A2(n_247),
.B1(n_215),
.B2(n_231),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_228),
.B1(n_225),
.B2(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

OA21x2_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_225),
.B(n_218),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_275),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_249),
.B(n_237),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_282),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_285),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_259),
.A2(n_225),
.B(n_224),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_288),
.B1(n_294),
.B2(n_295),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_248),
.C(n_245),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_297),
.C(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_229),
.B(n_219),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_221),
.B(n_226),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_255),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_241),
.B1(n_233),
.B2(n_216),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_268),
.B1(n_276),
.B2(n_258),
.Y(n_318)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_296),
.A2(n_299),
.B1(n_269),
.B2(n_255),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_239),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_239),
.C(n_252),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_308),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_279),
.B1(n_290),
.B2(n_261),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_309),
.B1(n_316),
.B2(n_293),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_304),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_252),
.C(n_257),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_311),
.C(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_257),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_280),
.A2(n_269),
.B1(n_265),
.B2(n_273),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_256),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_256),
.C(n_254),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_274),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_284),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_286),
.B1(n_281),
.B2(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_320),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_302),
.B1(n_313),
.B2(n_307),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_327),
.B1(n_330),
.B2(n_332),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_297),
.C(n_254),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_324),
.C(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_285),
.C(n_284),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_278),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_282),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_267),
.B1(n_281),
.B2(n_266),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_305),
.B1(n_306),
.B2(n_300),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_308),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_315),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_301),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_299),
.C(n_267),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_336),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_335),
.B(n_340),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_304),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_314),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_272),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_322),
.A2(n_294),
.B1(n_295),
.B2(n_276),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_258),
.C(n_282),
.Y(n_344)
);

OA21x2_ASAP7_75t_SL g351 ( 
.A1(n_345),
.A2(n_341),
.B(n_344),
.Y(n_351)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_350),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_338),
.A2(n_327),
.B1(n_326),
.B2(n_329),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_353),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_339),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_337),
.B1(n_319),
.B2(n_331),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_355),
.A2(n_358),
.B1(n_352),
.B2(n_334),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_347),
.A2(n_337),
.B(n_340),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_356),
.A2(n_346),
.B(n_348),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_331),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_357),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_361),
.Y(n_363)
);

AOI322xp5_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_263),
.A3(n_352),
.B1(n_354),
.B2(n_355),
.C1(n_358),
.C2(n_363),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_364),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_365),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_263),
.Y(n_367)
);


endmodule