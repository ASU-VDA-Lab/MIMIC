module fake_jpeg_11380_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_52),
.B(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_58),
.B(n_67),
.Y(n_134)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_61),
.B(n_64),
.Y(n_144)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_0),
.CON(n_66),
.SN(n_66)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_13),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_91),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_23),
.B1(n_46),
.B2(n_21),
.Y(n_102)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_98),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_97),
.Y(n_131)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_40),
.B1(n_36),
.B2(n_48),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_28),
.B1(n_36),
.B2(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_106),
.A2(n_136),
.B1(n_30),
.B2(n_54),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_109),
.B(n_114),
.Y(n_160)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_118),
.B(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_121),
.B(n_138),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_3),
.Y(n_180)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_48),
.B1(n_36),
.B2(n_34),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_41),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_34),
.B1(n_30),
.B2(n_42),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_89),
.B1(n_81),
.B2(n_77),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_21),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_41),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_31),
.B(n_24),
.C(n_71),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_154),
.A2(n_191),
.B(n_201),
.C(n_198),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_155),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_31),
.B(n_40),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_191),
.B(n_112),
.Y(n_212)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_93),
.B1(n_92),
.B2(n_90),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_159),
.A2(n_188),
.B1(n_199),
.B2(n_206),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_172),
.B1(n_179),
.B2(n_126),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_193),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_166),
.A2(n_182),
.B1(n_192),
.B2(n_108),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_48),
.B1(n_144),
.B2(n_146),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_170),
.B(n_176),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_1),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_34),
.B1(n_30),
.B2(n_73),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_202),
.Y(n_225)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_146),
.B1(n_128),
.B2(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_34),
.B1(n_30),
.B2(n_65),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_7),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_181),
.B(n_101),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_76),
.B1(n_74),
.B2(n_51),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_113),
.A2(n_19),
.B1(n_27),
.B2(n_70),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_19),
.C(n_12),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_195),
.Y(n_217)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_19),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_27),
.C(n_4),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_100),
.B(n_3),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_203),
.Y(n_231)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_128),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_5),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_122),
.B1(n_147),
.B2(n_125),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_115),
.B1(n_152),
.B2(n_153),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_150),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_209),
.A2(n_9),
.B1(n_10),
.B2(n_233),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_212),
.A2(n_253),
.B(n_206),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_218),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_241),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_147),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_101),
.C(n_151),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_250),
.C(n_200),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_159),
.A2(n_119),
.B1(n_143),
.B2(n_137),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_229),
.B1(n_201),
.B2(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_119),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_234),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_199),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_176),
.B1(n_161),
.B2(n_167),
.Y(n_229)
);

BUFx4f_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_236),
.B1(n_247),
.B2(n_248),
.Y(n_265)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_156),
.B(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_126),
.B1(n_143),
.B2(n_137),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_129),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_240),
.B(n_252),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_162),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_180),
.A2(n_154),
.B1(n_195),
.B2(n_189),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_157),
.A2(n_129),
.B1(n_103),
.B2(n_127),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_160),
.B(n_101),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_170),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_103),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_191),
.B(n_198),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_255),
.A2(n_282),
.B(n_296),
.Y(n_325)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_220),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_259),
.B(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_184),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_267),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_177),
.C(n_194),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_213),
.C(n_219),
.Y(n_327)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_178),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_268),
.B(n_269),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_272),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_163),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_273),
.A2(n_291),
.B1(n_297),
.B2(n_286),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_228),
.A2(n_117),
.B1(n_127),
.B2(n_186),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_175),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_285),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_239),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_287),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_151),
.B(n_171),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_243),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_117),
.B1(n_197),
.B2(n_152),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_229),
.A2(n_158),
.B1(n_174),
.B2(n_187),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_286),
.A2(n_248),
.B1(n_236),
.B2(n_242),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_239),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_232),
.A2(n_108),
.B1(n_10),
.B2(n_11),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_208),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_9),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_293),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_210),
.B(n_9),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_225),
.A2(n_10),
.B1(n_227),
.B2(n_237),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_210),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_10),
.B(n_217),
.Y(n_296)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_327),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_259),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_321),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_214),
.B(n_223),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_305),
.A2(n_315),
.B(n_323),
.Y(n_359)
);

CKINVDCx12_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_308),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_214),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_258),
.C(n_278),
.Y(n_352)
);

INVx6_ASAP7_75t_SL g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_310),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_274),
.A2(n_245),
.B(n_223),
.Y(n_315)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_292),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_255),
.A2(n_246),
.B(n_238),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_333),
.B1(n_289),
.B2(n_285),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_235),
.B(n_230),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_329),
.B(n_330),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_224),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_221),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_256),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_261),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_268),
.A2(n_221),
.B(n_230),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_272),
.B(n_256),
.C(n_265),
.D(n_269),
.Y(n_343)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_344),
.B1(n_358),
.B2(n_361),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_343),
.A2(n_302),
.B(n_328),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_322),
.A2(n_298),
.B1(n_275),
.B2(n_287),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_331),
.B1(n_319),
.B2(n_313),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_348),
.B1(n_266),
.B2(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_319),
.A2(n_273),
.B1(n_284),
.B2(n_278),
.Y(n_348)
);

O2A1O1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_325),
.A2(n_302),
.B(n_313),
.C(n_312),
.Y(n_349)
);

OAI31xp33_ASAP7_75t_L g371 ( 
.A1(n_349),
.A2(n_343),
.A3(n_359),
.B(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_356),
.C(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_353),
.B(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_284),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_363),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_263),
.C(n_279),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_265),
.B1(n_268),
.B2(n_271),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_307),
.A2(n_268),
.B1(n_271),
.B2(n_294),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_321),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_293),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_260),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_368),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_307),
.A2(n_266),
.B1(n_257),
.B2(n_270),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_367),
.A2(n_370),
.B1(n_318),
.B2(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_301),
.A2(n_276),
.B1(n_288),
.B2(n_264),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_371),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_382),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_309),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_387),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_358),
.A2(n_325),
.B1(n_305),
.B2(n_328),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_383),
.B1(n_392),
.B2(n_361),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_359),
.A2(n_329),
.B(n_323),
.C(n_310),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_389),
.C(n_374),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_376),
.B(n_377),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_365),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_363),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_336),
.B(n_306),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_339),
.B(n_324),
.Y(n_388)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_263),
.C(n_266),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_338),
.B(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_355),
.B(n_320),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_348),
.Y(n_406)
);

AOI21xp33_ASAP7_75t_L g396 ( 
.A1(n_357),
.A2(n_332),
.B(n_281),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_396),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_398),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_404),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_406),
.B(n_385),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_419),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_340),
.C(n_367),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_411),
.C(n_413),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_351),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_382),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_351),
.C(n_368),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_341),
.C(n_354),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_378),
.A2(n_342),
.B1(n_350),
.B2(n_347),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_414),
.Y(n_438)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_394),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_298),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_366),
.C(n_369),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_421),
.C(n_375),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_366),
.C(n_369),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_430),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_379),
.B1(n_381),
.B2(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_415),
.B(n_390),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_426),
.B(n_428),
.Y(n_445)
);

XNOR2x1_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_371),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_435),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_381),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_399),
.A2(n_394),
.B(n_375),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_419),
.B(n_421),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_420),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_397),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_433),
.B(n_436),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_375),
.C(n_393),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_408),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_440),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_402),
.A2(n_375),
.B(n_384),
.Y(n_439)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_439),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_397),
.Y(n_440)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_438),
.A2(n_410),
.B1(n_405),
.B2(n_423),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_411),
.C(n_413),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_452),
.C(n_453),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_422),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_412),
.B(n_406),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_449),
.A2(n_422),
.B(n_430),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_393),
.C(n_384),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_304),
.C(n_337),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_304),
.C(n_337),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_308),
.C(n_337),
.Y(n_467)
);

INVx11_ASAP7_75t_L g457 ( 
.A(n_452),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_453),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_454),
.A2(n_439),
.B(n_436),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_458),
.A2(n_461),
.B(n_463),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_449),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_460),
.B(n_465),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_439),
.B(n_432),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_462),
.A2(n_468),
.B(n_445),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_450),
.A2(n_442),
.B(n_441),
.Y(n_463)
);

FAx1_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_424),
.CI(n_440),
.CON(n_466),
.SN(n_466)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_444),
.Y(n_473)
);

NAND2x1_ASAP7_75t_SL g468 ( 
.A(n_444),
.B(n_316),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_470),
.B(n_472),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_473),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_447),
.C(n_451),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_299),
.A3(n_316),
.B1(n_455),
.B2(n_362),
.C1(n_297),
.C2(n_243),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_467),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_462),
.A2(n_455),
.B(n_362),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_468),
.B(n_477),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_464),
.C(n_458),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_456),
.C(n_457),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_479),
.A2(n_481),
.B(n_464),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_463),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_483),
.A2(n_477),
.B(n_469),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_485),
.Y(n_487)
);

AOI321xp33_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_480),
.A3(n_479),
.B1(n_482),
.B2(n_466),
.C(n_459),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_480),
.C(n_461),
.Y(n_489)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_487),
.B(n_466),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_299),
.Y(n_491)
);


endmodule