module fake_jpeg_13714_n_519 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_55),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_20),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_56),
.B(n_57),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_60),
.B(n_65),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_8),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_77),
.Y(n_155)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_33),
.B(n_8),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_34),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_83),
.B(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_34),
.B(n_7),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_24),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_134),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_88),
.B1(n_81),
.B2(n_66),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_139),
.B1(n_142),
.B2(n_23),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_29),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_32),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_121),
.B(n_69),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_59),
.B(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_32),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_50),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_46),
.B1(n_16),
.B2(n_39),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_55),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_74),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_158),
.B1(n_30),
.B2(n_47),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_80),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_173),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_170),
.Y(n_235)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_167),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_110),
.A2(n_68),
.B1(n_64),
.B2(n_93),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_168),
.A2(n_192),
.B1(n_200),
.B2(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_169),
.Y(n_214)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_174),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_30),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

AND2x4_ASAP7_75t_SL g178 ( 
.A(n_107),
.B(n_24),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_178),
.Y(n_245)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_29),
.B(n_49),
.C(n_47),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_181),
.A2(n_123),
.A3(n_45),
.B1(n_40),
.B2(n_42),
.Y(n_234)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_184),
.B(n_185),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_134),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_191),
.Y(n_211)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_25),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_126),
.A2(n_96),
.B1(n_91),
.B2(n_23),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_42),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_194),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_41),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_102),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_120),
.B1(n_123),
.B2(n_42),
.Y(n_240)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_203),
.Y(n_221)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_206),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_136),
.A2(n_23),
.B1(n_38),
.B2(n_47),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_119),
.A2(n_94),
.B1(n_63),
.B2(n_53),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_115),
.B(n_23),
.Y(n_215)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_120),
.Y(n_224)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_112),
.B1(n_119),
.B2(n_147),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_167),
.B(n_206),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_178),
.B(n_122),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_108),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_234),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_166),
.A2(n_129),
.B1(n_136),
.B2(n_125),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_168),
.B1(n_192),
.B2(n_205),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_108),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_177),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_177),
.C(n_161),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_201),
.C(n_195),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_195),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_164),
.C(n_133),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_258),
.C(n_268),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_203),
.C(n_190),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_283),
.B1(n_265),
.B2(n_267),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_166),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_186),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_189),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_228),
.A2(n_207),
.B1(n_105),
.B2(n_118),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_267),
.B1(n_282),
.B2(n_283),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_235),
.A2(n_245),
.B1(n_226),
.B2(n_211),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_133),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_218),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_198),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_281),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_284),
.B(n_238),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_225),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_197),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_231),
.C(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_180),
.C(n_165),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_235),
.A2(n_182),
.B1(n_105),
.B2(n_125),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_226),
.A2(n_117),
.B1(n_118),
.B2(n_140),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_215),
.A2(n_29),
.B(n_25),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_230),
.B1(n_232),
.B2(n_200),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_296),
.B1(n_297),
.B2(n_216),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_242),
.B1(n_216),
.B2(n_238),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_286),
.A2(n_243),
.B1(n_248),
.B2(n_212),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_306),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_266),
.B1(n_275),
.B2(n_281),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_249),
.A2(n_230),
.B1(n_214),
.B2(n_117),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_249),
.A2(n_214),
.B1(n_162),
.B2(n_227),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_299),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_227),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_250),
.B(n_261),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_233),
.B1(n_237),
.B2(n_220),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_233),
.B1(n_220),
.B2(n_260),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_246),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_246),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_237),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_315),
.A2(n_216),
.B(n_210),
.Y(n_339)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_331),
.B1(n_336),
.B2(n_351),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_252),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_322),
.B(n_325),
.C(n_338),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_323),
.B(n_324),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_307),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_253),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_327),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_258),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_328),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_299),
.B(n_250),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g369 ( 
.A1(n_329),
.A2(n_347),
.B(n_349),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_305),
.A2(n_255),
.B1(n_271),
.B2(n_257),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_315),
.A2(n_256),
.B(n_210),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_334),
.A2(n_339),
.B(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_341),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_305),
.A2(n_223),
.B1(n_212),
.B2(n_280),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_343),
.B1(n_353),
.B2(n_310),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_319),
.C(n_299),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_244),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_346),
.C(n_299),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_298),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_293),
.A2(n_244),
.B(n_243),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_248),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_209),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_348),
.B(n_289),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_301),
.A2(n_241),
.B(n_225),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_310),
.A2(n_159),
.B1(n_150),
.B2(n_241),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_297),
.A2(n_296),
.B1(n_285),
.B2(n_300),
.Y(n_353)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_325),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_359),
.B(n_370),
.Y(n_411)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_384),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_367),
.B1(n_347),
.B2(n_351),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_292),
.B1(n_291),
.B2(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_368),
.C(n_355),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_337),
.A2(n_300),
.B1(n_317),
.B2(n_301),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_318),
.C(n_287),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_338),
.B(n_298),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_308),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_381),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_287),
.B1(n_290),
.B2(n_291),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_383),
.B1(n_385),
.B2(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_320),
.B(n_290),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_304),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_380),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_313),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_347),
.A2(n_295),
.B1(n_304),
.B2(n_289),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_295),
.B1(n_304),
.B2(n_302),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_377),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_346),
.C(n_328),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_396),
.C(n_398),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_327),
.Y(n_392)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_330),
.B1(n_328),
.B2(n_326),
.Y(n_395)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_366),
.C(n_368),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g397 ( 
.A(n_359),
.B(n_330),
.CI(n_334),
.CON(n_397),
.SN(n_397)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_369),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_381),
.C(n_357),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_400),
.A2(n_371),
.B1(n_378),
.B2(n_380),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_342),
.C(n_339),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_410),
.C(n_412),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_377),
.A2(n_327),
.B(n_302),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_404),
.A2(n_21),
.B(n_9),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_38),
.B1(n_49),
.B2(n_45),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_414),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_172),
.C(n_49),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_45),
.C(n_41),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_371),
.A2(n_41),
.B1(n_40),
.B2(n_25),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_40),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_383),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_420),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_387),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_439),
.B1(n_414),
.B2(n_415),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_426),
.Y(n_459)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_391),
.C(n_396),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_437),
.C(n_438),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_394),
.B(n_375),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_432),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_394),
.B(n_386),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_397),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_436),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_21),
.C(n_1),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_0),
.C(n_1),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_7),
.B1(n_13),
.B2(n_2),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_390),
.B1(n_402),
.B2(n_393),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_441),
.A2(n_446),
.B1(n_433),
.B2(n_427),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_434),
.A2(n_404),
.B(n_398),
.Y(n_442)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_411),
.C(n_395),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_444),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_411),
.C(n_410),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_425),
.A2(n_412),
.B1(n_388),
.B2(n_401),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_449),
.B(n_418),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_409),
.C(n_397),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_453),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_452),
.A2(n_427),
.B1(n_438),
.B2(n_436),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_0),
.C(n_1),
.Y(n_453)
);

FAx1_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_9),
.CI(n_2),
.CON(n_455),
.SN(n_455)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_439),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_431),
.B1(n_419),
.B2(n_428),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_460),
.A2(n_476),
.B1(n_4),
.B2(n_9),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_431),
.B(n_435),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_458),
.B(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_450),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_466),
.B(n_440),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_418),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_452),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_437),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_455),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_444),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_475),
.Y(n_490)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_459),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_474),
.B(n_458),
.Y(n_481)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_456),
.A2(n_10),
.B1(n_4),
.B2(n_6),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_465),
.A2(n_471),
.B1(n_462),
.B2(n_474),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_478),
.Y(n_498)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_440),
.C(n_453),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_476),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_488),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_469),
.A2(n_455),
.B(n_448),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_487),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_472),
.A2(n_10),
.B(n_12),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_460),
.A2(n_10),
.B(n_13),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_14),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_461),
.C(n_463),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_496),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_13),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_497),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_501),
.A2(n_0),
.B1(n_488),
.B2(n_498),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_14),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_502),
.B(n_489),
.Y(n_507)
);

O2A1O1Ixp33_ASAP7_75t_SL g504 ( 
.A1(n_500),
.A2(n_483),
.B(n_480),
.C(n_486),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_504),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_494),
.A2(n_491),
.B(n_482),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_505),
.A2(n_500),
.B(n_492),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_507),
.B(n_508),
.Y(n_511)
);

NOR3xp33_ASAP7_75t_SL g508 ( 
.A(n_493),
.B(n_478),
.C(n_485),
.Y(n_508)
);

OAI21x1_ASAP7_75t_SL g510 ( 
.A1(n_509),
.A2(n_499),
.B(n_498),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_510),
.B(n_512),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_511),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_506),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_514),
.C(n_513),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_517),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_503),
.Y(n_519)
);


endmodule