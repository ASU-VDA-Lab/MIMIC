module real_jpeg_18386_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_3),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_3),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_3),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_3),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_3),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_3),
.B(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_4),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_100),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_5),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g433 ( 
.A(n_6),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_7),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_7),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_8),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_13),
.B1(n_220),
.B2(n_223),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_8),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_8),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_8),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_8),
.B(n_194),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_8),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_8),
.B(n_439),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_9),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_9),
.B(n_200),
.Y(n_199)
);

AND2x4_ASAP7_75t_SL g243 ( 
.A(n_9),
.B(n_244),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_9),
.B(n_293),
.Y(n_292)
);

AND2x4_ASAP7_75t_SL g345 ( 
.A(n_9),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_9),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_10),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_10),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_10),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_10),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_10),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_10),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_10),
.B(n_454),
.Y(n_453)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_12),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_12),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_12),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_12),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_12),
.B(n_50),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_13),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_13),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_13),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_13),
.B(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_13),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_14),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_15),
.B(n_74),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_15),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_231),
.Y(n_230)
);

AND2x4_ASAP7_75t_SL g248 ( 
.A(n_15),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_15),
.B(n_50),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g137 ( 
.A(n_16),
.Y(n_137)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_208),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_206),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_157),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_21),
.B(n_157),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_95),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.C(n_87),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_51),
.Y(n_24)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_25),
.B(n_40),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_26),
.B(n_31),
.C(n_36),
.Y(n_152)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_28),
.Y(n_249)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_39),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_49),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_41),
.B(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_45),
.A2(n_49),
.B1(n_65),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_45),
.Y(n_166)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_48),
.Y(n_231)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_48),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_53),
.C(n_60),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_51),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_52),
.B(n_228),
.C(n_230),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_52),
.A2(n_53),
.B1(n_230),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_66),
.B1(n_103),
.B2(n_104),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_64),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_104),
.C(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_67),
.B(n_87),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.C(n_81),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_68),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.C(n_75),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_69),
.B(n_75),
.Y(n_181)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_73),
.B(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_78),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_89),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_90),
.C(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_85),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_86),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_90),
.B(n_184),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_90),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_131),
.B1(n_155),
.B2(n_156),
.Y(n_95)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_113),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_99),
.Y(n_107)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_126),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_126),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_149),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_148),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_153),
.Y(n_149)
);

XNOR2x2_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_158),
.B(n_160),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_162),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_182),
.C(n_203),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_163),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_180),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_164),
.B(n_167),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.C(n_175),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_168),
.A2(n_175),
.B1(n_176),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_168),
.Y(n_305)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_172),
.B(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_175),
.B(n_369),
.C(n_372),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_175),
.A2(n_176),
.B1(n_369),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_178),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

XNOR2x2_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_182),
.B(n_203),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.C(n_198),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_183),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_188),
.Y(n_217)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_185),
.Y(n_440)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_191),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_198),
.A2(n_199),
.B1(n_349),
.B2(n_350),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_199),
.B(n_344),
.C(n_349),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_202),
.Y(n_335)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_313),
.B(n_483),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_306),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_267),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_212),
.B(n_267),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_259),
.Y(n_212)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_213),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_232),
.C(n_255),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_227),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_216),
.B(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_218),
.A2(n_219),
.B1(n_227),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_219),
.A2(n_329),
.B(n_336),
.Y(n_328)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_222),
.Y(n_399)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_226),
.Y(n_371)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_227),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_233),
.A2(n_256),
.B1(n_257),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_247),
.C(n_250),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.C(n_243),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_235),
.A2(n_243),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_239),
.B(n_325),
.Y(n_324)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_243),
.B(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_262),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.C(n_275),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_269),
.A2(n_270),
.B1(n_273),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_299),
.C(n_303),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_277),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.C(n_287),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_279),
.B(n_378),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_282),
.B(n_287),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_283),
.B(n_286),
.Y(n_376)
);

NOR2x1_ASAP7_75t_R g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.C(n_296),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_292),
.A2(n_296),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_292),
.B(n_428),
.C(n_430),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_292),
.A2(n_366),
.B1(n_430),
.B2(n_431),
.Y(n_443)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_294),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_295),
.Y(n_449)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_303),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_306),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_307),
.B(n_309),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_379),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.C(n_356),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_316),
.B(n_320),
.Y(n_482)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_353),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_353),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.C(n_343),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_328),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_387),
.C(n_391),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_344),
.B(n_470),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_348),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_345),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_345),
.A2(n_437),
.B1(n_438),
.B2(n_451),
.Y(n_450)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_357),
.B(n_359),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.C(n_377),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_360),
.B(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_362),
.B(n_377),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.C(n_375),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_363),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_368),
.B(n_376),
.Y(n_465)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_412),
.Y(n_411)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_481),
.C(n_482),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_476),
.B(n_480),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_461),
.B(n_475),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_422),
.B(n_460),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_408),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_384),
.B(n_408),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_392),
.C(n_400),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_392),
.A2(n_393),
.B1(n_400),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_394),
.B(n_398),
.Y(n_429)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

AO22x1_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_400)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_401),
.Y(n_406)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_404),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_406),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_414),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_410),
.B(n_414),
.C(n_474),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_417),
.C(n_418),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_434),
.B(n_459),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_SL g459 ( 
.A(n_424),
.B(n_427),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_429),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_444),
.B(n_458),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_441),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_441),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_452),
.B(n_457),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_450),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_450),
.Y(n_457)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_473),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_SL g475 ( 
.A(n_462),
.B(n_473),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_468),
.C(n_472),
.Y(n_477)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_472),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_478),
.Y(n_480)
);


endmodule