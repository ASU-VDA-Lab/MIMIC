module fake_jpeg_29745_n_74 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx13_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_18),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_1),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_28),
.C(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_11),
.B(n_22),
.C(n_21),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_10),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_30),
.C(n_26),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_39),
.B1(n_8),
.B2(n_14),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.C(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_20),
.C(n_19),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.C(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_61),
.B1(n_7),
.B2(n_60),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_15),
.B1(n_16),
.B2(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_64),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);


endmodule