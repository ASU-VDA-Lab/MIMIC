module fake_jpeg_12216_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_6),
.B(n_38),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_57),
.B1(n_53),
.B2(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_60),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_5),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_66),
.B1(n_52),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_52),
.B1(n_60),
.B2(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_65),
.B1(n_51),
.B2(n_50),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_67),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_8),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_101),
.B1(n_102),
.B2(n_12),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_50),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_16),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_104),
.C(n_74),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_15),
.C(n_41),
.Y(n_99)
);

NOR2x1p5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_1),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_81),
.Y(n_107)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_9),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_10),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_81),
.B1(n_35),
.B2(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_11),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_103),
.B1(n_20),
.B2(n_21),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_123),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_128),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_37),
.C(n_26),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_33),
.C(n_36),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_123),
.C(n_122),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_130),
.B1(n_105),
.B2(n_126),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_105),
.C(n_12),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_134),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_141),
.B(n_124),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_140),
.C(n_142),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_133),
.B(n_136),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_135),
.B(n_129),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_125),
.B(n_40),
.C(n_43),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_39),
.B(n_117),
.Y(n_148)
);

OAI21x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_121),
.B(n_126),
.Y(n_149)
);


endmodule