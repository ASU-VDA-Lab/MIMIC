module real_jpeg_25888_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_32),
.B1(n_72),
.B2(n_74),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_32),
.B1(n_50),
.B2(n_51),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_2),
.A2(n_37),
.B1(n_40),
.B2(n_65),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_65),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_4),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_43),
.B1(n_72),
.B2(n_95),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_61),
.B(n_66),
.C(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_59),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_49),
.B(n_50),
.C(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_23),
.C(n_39),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_4),
.B(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_4),
.B(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_4),
.B(n_41),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_24),
.B1(n_37),
.B2(n_40),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_137),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_136),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_112),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_16),
.B(n_112),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_76),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.C(n_57),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_18),
.A2(n_19),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_33),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_27),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_21),
.A2(n_85),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_23),
.B(n_224),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_31),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_25),
.A2(n_84),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_25),
.B(n_84),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_25),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_28),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_28),
.B(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_44),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_34),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_42),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_35),
.B(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_35),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_40),
.B1(n_49),
.B2(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_37),
.B(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_40),
.A2(n_43),
.B(n_53),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_41),
.B(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_42),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_43),
.A2(n_50),
.B(n_60),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_44),
.A2(n_88),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_44),
.B(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_46),
.A2(n_57),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_46),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_55),
.Y(n_46)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_47),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_47),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_48)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_54),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_73),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_68),
.Y(n_96)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_94),
.Y(n_146)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_104),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_80),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_85),
.B(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_87),
.A2(n_110),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_87),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_89),
.B(n_196),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_124),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_102),
.B(n_153),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_105),
.A2(n_111),
.B1(n_180),
.B2(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.C(n_135),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_113),
.A2(n_114),
.B1(n_135),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_119),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_128),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_173),
.B(n_249),
.C(n_254),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_161),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_139),
.B(n_161),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_157),
.B2(n_160),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_155),
.B2(n_156),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_142),
.B(n_156),
.C(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_163),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_171),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_248),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_190),
.B(n_247),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_176),
.B(n_187),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_182),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_182),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_242),
.B(n_246),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_233),
.B(n_241),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_213),
.B(n_232),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_220),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_195),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_207),
.B2(n_212),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_206),
.C(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_231),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);


endmodule