module fake_netlist_5_1945_n_1887 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1887);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1887;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_100),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_33),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_44),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_48),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_17),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_99),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_82),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_66),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_57),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_64),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_43),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_44),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_57),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_63),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_85),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_68),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_67),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_101),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_45),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_97),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_27),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_42),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_1),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_77),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_29),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_79),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_125),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_116),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_89),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_142),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_110),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_122),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_22),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_74),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_28),
.Y(n_249)
);

CKINVDCx12_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_119),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_62),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_23),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_164),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_9),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_103),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_124),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_43),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_15),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_52),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_19),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_73),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_39),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_35),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_23),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_45),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_70),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_154),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_55),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_130),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_173),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_95),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_55),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_166),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_67),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_132),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_31),
.B(n_30),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_37),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_106),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_171),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_7),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_41),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_121),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_59),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_5),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_149),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_98),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_120),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_80),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_115),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_30),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_5),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_75),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_83),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_27),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_134),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_18),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_54),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_13),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_87),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_138),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_36),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_50),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_31),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_65),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_6),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_18),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_140),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_53),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_88),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_52),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_144),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_59),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_21),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_2),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_24),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_47),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_126),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_69),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_65),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_46),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_4),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_36),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_91),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_26),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_49),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_14),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_4),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_135),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_204),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_229),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_229),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_229),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_177),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_229),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_191),
.B(n_0),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_230),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_182),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_194),
.B(n_0),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_194),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_229),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_231),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_231),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_219),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_191),
.B(n_2),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_179),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_179),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_183),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_192),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_203),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_184),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_184),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_187),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_236),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_197),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_200),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_187),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_201),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_205),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_181),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_211),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_204),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_220),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_211),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_221),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_214),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_218),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_218),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_225),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_228),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_224),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_232),
.B(n_175),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_233),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_178),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_224),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_R g407 ( 
.A(n_238),
.B(n_137),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_240),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_265),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_178),
.B(n_6),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_181),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_242),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_265),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_270),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_244),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_257),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_270),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_274),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_305),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_274),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_275),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_275),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_266),
.B(n_7),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_284),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_266),
.B(n_10),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_203),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_259),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_278),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_284),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_282),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_186),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_213),
.B(n_12),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_213),
.B(n_12),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_285),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_285),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_283),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_180),
.B(n_16),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_288),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_288),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_356),
.B(n_243),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_356),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_357),
.B(n_286),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_354),
.B(n_243),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_412),
.B(n_208),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_362),
.A2(n_208),
.B1(n_293),
.B2(n_223),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_359),
.B(n_289),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_361),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_354),
.B(n_246),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_367),
.B(n_354),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_391),
.B(n_299),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_308),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_373),
.A2(n_327),
.B1(n_337),
.B2(n_252),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_438),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_412),
.B(n_215),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_374),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_433),
.A2(n_293),
.B1(n_258),
.B2(n_269),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_365),
.B(n_239),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_434),
.B(n_239),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_363),
.B(n_383),
.Y(n_476)
);

NAND2x1_ASAP7_75t_L g477 ( 
.A(n_365),
.B(n_309),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_420),
.B(n_309),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_368),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_368),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_432),
.B(n_360),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_369),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_375),
.B(n_311),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_380),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_370),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_382),
.B(n_315),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_246),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_370),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_372),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_382),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_386),
.B(n_346),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_372),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_317),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_371),
.A2(n_226),
.B1(n_329),
.B2(n_216),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_411),
.B(n_346),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_364),
.B(n_215),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_396),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_396),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_397),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_464),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_460),
.B(n_462),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_464),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_424),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_460),
.B(n_376),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_478),
.B(n_377),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_476),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_456),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_470),
.B(n_384),
.C(n_378),
.Y(n_541)
);

INVxp33_ASAP7_75t_SL g542 ( 
.A(n_476),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_385),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

AND2x2_ASAP7_75t_SL g547 ( 
.A(n_475),
.B(n_472),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_462),
.B(n_387),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_486),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_486),
.B(n_388),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_475),
.B(n_424),
.C(n_426),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_499),
.B(n_394),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_484),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_499),
.B(n_400),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_472),
.B(n_413),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_470),
.A2(n_508),
.B1(n_463),
.B2(n_449),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_455),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_510),
.B(n_417),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_446),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_454),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_454),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_472),
.A2(n_426),
.B1(n_351),
.B2(n_277),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_471),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_447),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_472),
.A2(n_277),
.B1(n_351),
.B2(n_347),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_466),
.B(n_428),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_446),
.B(n_180),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_441),
.B(n_456),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_446),
.B(n_185),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_452),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_486),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_509),
.A2(n_347),
.B1(n_300),
.B2(n_307),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_466),
.B(n_405),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_509),
.B(n_429),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_458),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_458),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_455),
.Y(n_594)
);

AO22x2_ASAP7_75t_L g595 ( 
.A1(n_449),
.A2(n_292),
.B1(n_296),
.B2(n_301),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_509),
.A2(n_392),
.B1(n_404),
.B2(n_401),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_463),
.A2(n_321),
.B1(n_210),
.B2(n_212),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_473),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_444),
.B(n_431),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_505),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_488),
.B(n_437),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_505),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_473),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_505),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_505),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_477),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_444),
.B(n_196),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_495),
.A2(n_501),
.B1(n_494),
.B2(n_488),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_185),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_486),
.B(n_408),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_516),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_495),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_500),
.B(n_409),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_516),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_500),
.B(n_467),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_516),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_450),
.B(n_247),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_494),
.B(n_403),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_480),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_455),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_480),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_516),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_500),
.B(n_416),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_507),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_480),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_451),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_453),
.A2(n_291),
.B1(n_290),
.B2(n_287),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_507),
.B(n_405),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_455),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_500),
.B(n_407),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_450),
.B(n_251),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_455),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_451),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_501),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_461),
.B(n_358),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_508),
.B(n_461),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_459),
.B(n_281),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_469),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_451),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_459),
.B(n_298),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_501),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_457),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_469),
.B(n_193),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_482),
.A2(n_254),
.B1(n_245),
.B2(n_345),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_482),
.B(n_330),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_457),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_489),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_490),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_459),
.B(n_323),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_490),
.B(n_190),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_457),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_492),
.B(n_493),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_459),
.B(n_193),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_492),
.B(n_402),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_493),
.A2(n_300),
.B1(n_292),
.B2(n_296),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_498),
.B(n_209),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_459),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_498),
.B(n_217),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_459),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_SL g667 ( 
.A(n_502),
.B(n_234),
.C(n_227),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_459),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_502),
.B(n_402),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_504),
.B(n_215),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_627),
.B(n_468),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_627),
.B(n_468),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_547),
.B(n_468),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_531),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_547),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_553),
.A2(n_222),
.B1(n_207),
.B2(n_206),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_538),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_519),
.B(n_468),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_547),
.B(n_468),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_592),
.B(n_468),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_584),
.B(n_504),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_562),
.B(n_249),
.C(n_235),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_565),
.A2(n_352),
.B1(n_215),
.B2(n_333),
.Y(n_685)
);

AND2x4_ASAP7_75t_SL g686 ( 
.A(n_523),
.B(n_352),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_592),
.B(n_468),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_520),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_584),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_593),
.B(n_474),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_521),
.Y(n_691)
);

BUFx5_ASAP7_75t_L g692 ( 
.A(n_581),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_580),
.B(n_253),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_593),
.B(n_474),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_602),
.B(n_474),
.Y(n_695)
);

BUFx5_ASAP7_75t_L g696 ( 
.A(n_581),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_614),
.B(n_474),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_614),
.B(n_474),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_529),
.Y(n_699)
);

OAI22x1_ASAP7_75t_SL g700 ( 
.A1(n_542),
.A2(n_271),
.B1(n_279),
.B2(n_276),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_553),
.A2(n_302),
.B1(n_198),
.B2(n_199),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_584),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_543),
.B(n_255),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_554),
.B(n_560),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_610),
.B(n_474),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_631),
.B(n_474),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_530),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_522),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_551),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_600),
.B(n_256),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_567),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_522),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_524),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_609),
.B(n_496),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_523),
.B(n_305),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_529),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_619),
.B(n_496),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_635),
.B(n_496),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_540),
.B(n_506),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_496),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_523),
.B(n_607),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_533),
.B(n_496),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_548),
.B(n_496),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_532),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_524),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_523),
.B(n_305),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_541),
.B(n_262),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_639),
.B(n_496),
.Y(n_730)
);

AO221x1_ASAP7_75t_L g731 ( 
.A1(n_595),
.A2(n_650),
.B1(n_630),
.B2(n_596),
.C(n_304),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_607),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_574),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_528),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_532),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_608),
.B(n_305),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_639),
.B(n_512),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_530),
.A2(n_195),
.B1(n_202),
.B2(n_206),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_647),
.B(n_512),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_608),
.B(n_305),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_528),
.B(n_305),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_647),
.B(n_512),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_611),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_530),
.A2(n_306),
.B1(n_207),
.B2(n_222),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_534),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_644),
.B(n_515),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_640),
.B(n_506),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_530),
.A2(n_332),
.B1(n_237),
.B2(n_248),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_534),
.B(n_334),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_661),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_661),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_644),
.B(n_653),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_561),
.B(n_263),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_597),
.B(n_340),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_581),
.B(n_202),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_546),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_620),
.A2(n_250),
.B1(n_237),
.B2(n_322),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_653),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_654),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_654),
.B(n_515),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_623),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_546),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_590),
.B(n_268),
.C(n_264),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_655),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_622),
.A2(n_248),
.B(n_260),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_597),
.B(n_260),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_511),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_655),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_623),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_669),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_611),
.B(n_511),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_611),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_659),
.B(n_515),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_669),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_556),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_556),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_649),
.B(n_513),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_557),
.B(n_261),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_611),
.B(n_513),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_557),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_530),
.A2(n_261),
.B1(n_267),
.B2(n_294),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_657),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_611),
.B(n_514),
.Y(n_783)
);

INVx8_ASAP7_75t_L g784 ( 
.A(n_581),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_663),
.B(n_665),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_558),
.Y(n_786)
);

BUFx6f_ASAP7_75t_SL g787 ( 
.A(n_649),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_558),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_564),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_649),
.B(n_517),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_597),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_564),
.Y(n_792)
);

AO221x1_ASAP7_75t_L g793 ( 
.A1(n_595),
.A2(n_341),
.B1(n_303),
.B2(n_304),
.C(n_307),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_566),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_549),
.B(n_352),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_566),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_597),
.B(n_267),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_569),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_601),
.B(n_294),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_601),
.B(n_297),
.Y(n_800)
);

AO21x2_ASAP7_75t_L g801 ( 
.A1(n_656),
.A2(n_306),
.B(n_302),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_603),
.B(n_297),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_569),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_581),
.B(n_310),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_598),
.A2(n_332),
.B1(n_322),
.B2(n_314),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_571),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_660),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_571),
.B(n_310),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_537),
.B(n_641),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_314),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_605),
.B(n_517),
.Y(n_811)
);

NOR3xp33_ASAP7_75t_L g812 ( 
.A(n_667),
.B(n_320),
.C(n_272),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_538),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_591),
.A2(n_250),
.B1(n_352),
.B2(n_491),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_605),
.B(n_481),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_518),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_518),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_606),
.B(n_481),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_531),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_581),
.A2(n_319),
.B1(n_349),
.B2(n_343),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_670),
.B(n_273),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_606),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_649),
.Y(n_823)
);

BUFx5_ASAP7_75t_L g824 ( 
.A(n_581),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_598),
.B(n_295),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_643),
.B(n_481),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_646),
.B(n_483),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_589),
.B(n_651),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_531),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_664),
.B(n_483),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_649),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_660),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_572),
.B(n_295),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_526),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_595),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_664),
.B(n_483),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_660),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_666),
.B(n_503),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_575),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_526),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_586),
.B(n_406),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_705),
.B(n_577),
.C(n_617),
.Y(n_842)
);

BUFx8_ASAP7_75t_L g843 ( 
.A(n_733),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_706),
.A2(n_666),
.B(n_578),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_782),
.B(n_559),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_710),
.B(n_588),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_785),
.B(n_586),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_671),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_704),
.B(n_586),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_680),
.A2(n_578),
.B(n_575),
.Y(n_850)
);

AND2x2_ASAP7_75t_SL g851 ( 
.A(n_677),
.B(n_301),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_671),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_550),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_678),
.A2(n_634),
.B(n_587),
.C(n_582),
.Y(n_854)
);

CKINVDCx10_ASAP7_75t_R g855 ( 
.A(n_679),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_693),
.B(n_586),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_674),
.A2(n_587),
.B(n_582),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_688),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_688),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_695),
.A2(n_535),
.B(n_531),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_711),
.B(n_586),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_712),
.B(n_767),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_674),
.A2(n_535),
.B(n_531),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_809),
.A2(n_586),
.B1(n_615),
.B2(n_612),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_681),
.A2(n_555),
.B(n_535),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_709),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_713),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_721),
.B(n_588),
.Y(n_869)
);

AO21x1_ASAP7_75t_L g870 ( 
.A1(n_744),
.A2(n_616),
.B(n_613),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_777),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_707),
.B(n_758),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_683),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_759),
.B(n_586),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_764),
.B(n_536),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_768),
.B(n_536),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_681),
.A2(n_544),
.B(n_536),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_675),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_675),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_682),
.A2(n_555),
.B(n_535),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_687),
.A2(n_555),
.B(n_535),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_724),
.A2(n_563),
.B(n_555),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_770),
.B(n_595),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_776),
.B(n_544),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_725),
.A2(n_563),
.B(n_555),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_697),
.A2(n_616),
.B(n_613),
.Y(n_886)
);

CKINVDCx10_ASAP7_75t_R g887 ( 
.A(n_679),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_713),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_702),
.A2(n_626),
.B(n_629),
.C(n_637),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_780),
.B(n_544),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_828),
.A2(n_662),
.B(n_325),
.C(n_319),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_675),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_719),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_685),
.B(n_312),
.C(n_280),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_835),
.B(n_542),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_675),
.Y(n_896)
);

AOI33xp33_ASAP7_75t_L g897 ( 
.A1(n_774),
.A2(n_406),
.A3(n_410),
.B1(n_414),
.B2(n_415),
.B3(n_418),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_722),
.A2(n_570),
.B(n_563),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_786),
.B(n_552),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_738),
.A2(n_668),
.B1(n_552),
.B2(n_579),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_691),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_788),
.B(n_552),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_792),
.B(n_579),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_672),
.A2(n_570),
.B(n_563),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_673),
.A2(n_570),
.B(n_563),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_794),
.B(n_579),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_714),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_683),
.B(n_410),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_714),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

NOR2x1_ASAP7_75t_L g911 ( 
.A(n_723),
.B(n_618),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_826),
.A2(n_594),
.B(n_570),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_715),
.A2(n_594),
.B(n_570),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_718),
.A2(n_594),
.B(n_633),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_796),
.B(n_633),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_798),
.B(n_633),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_692),
.B(n_660),
.Y(n_917)
);

OR2x6_ASAP7_75t_SL g918 ( 
.A(n_813),
.B(n_313),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_720),
.A2(n_594),
.B(n_636),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_813),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_691),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_803),
.B(n_636),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_806),
.B(n_636),
.Y(n_923)
);

BUFx4_ASAP7_75t_SL g924 ( 
.A(n_763),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_690),
.A2(n_594),
.B(n_668),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_732),
.B(n_668),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_734),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_747),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_732),
.B(n_527),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_694),
.A2(n_525),
.B(n_618),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_692),
.B(n_625),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_752),
.B(n_527),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_734),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_756),
.B(n_539),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_716),
.A2(n_728),
.B(n_827),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_762),
.B(n_545),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_795),
.B(n_295),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_762),
.B(n_545),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_691),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_775),
.B(n_568),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_819),
.A2(n_525),
.B(n_625),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_748),
.A2(n_632),
.B1(n_638),
.B2(n_642),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_825),
.B(n_632),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_692),
.B(n_638),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_723),
.A2(n_642),
.B1(n_660),
.B2(n_573),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_775),
.B(n_568),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_750),
.B(n_295),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_745),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_716),
.A2(n_599),
.B(n_576),
.Y(n_949)
);

AOI21xp33_ASAP7_75t_L g950 ( 
.A1(n_729),
.A2(n_316),
.B(n_318),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_745),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_692),
.B(n_573),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_691),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_692),
.B(n_576),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_819),
.A2(n_525),
.B(n_628),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_751),
.A2(n_303),
.B(n_325),
.C(n_335),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_819),
.A2(n_525),
.B(n_628),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_753),
.B(n_333),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_676),
.A2(n_525),
.B(n_583),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_789),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_730),
.A2(n_791),
.B(n_827),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_791),
.B(n_583),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_789),
.B(n_585),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_816),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_783),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_791),
.A2(n_525),
.B(n_585),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_773),
.B(n_599),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_697),
.A2(n_624),
.B(n_604),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_686),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_692),
.B(n_604),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_805),
.A2(n_645),
.B(n_658),
.C(n_652),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_700),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_698),
.A2(n_624),
.B(n_621),
.Y(n_973)
);

AOI33xp33_ASAP7_75t_L g974 ( 
.A1(n_833),
.A2(n_414),
.A3(n_440),
.B1(n_439),
.B2(n_436),
.B3(n_435),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_683),
.B(n_621),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_698),
.A2(n_637),
.B(n_658),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_728),
.A2(n_629),
.B(n_652),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_765),
.B(n_645),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_822),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_772),
.B(n_324),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_781),
.A2(n_648),
.B1(n_326),
.B2(n_344),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_684),
.B(n_328),
.C(n_331),
.Y(n_982)
);

AND2x6_ASAP7_75t_L g983 ( 
.A(n_807),
.B(n_648),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_686),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_699),
.B(n_660),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_741),
.A2(n_660),
.B(n_503),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_L g987 ( 
.A(n_812),
.B(n_339),
.C(n_338),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_692),
.B(n_485),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_821),
.B(n_349),
.C(n_335),
.Y(n_989)
);

NOR2x2_ASAP7_75t_L g990 ( 
.A(n_731),
.B(n_333),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_771),
.B(n_779),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_816),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_737),
.A2(n_503),
.B(n_497),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_799),
.A2(n_343),
.B(n_336),
.C(n_341),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_SL g995 ( 
.A1(n_708),
.A2(n_342),
.B(n_336),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_699),
.B(n_497),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_739),
.A2(n_497),
.B(n_491),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_699),
.B(n_485),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_777),
.B(n_485),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_689),
.B(n_415),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_701),
.A2(n_491),
.B1(n_487),
.B2(n_440),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_839),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_696),
.B(n_487),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_777),
.B(n_487),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_703),
.B(n_16),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_741),
.A2(n_342),
.B(n_436),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_696),
.B(n_333),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_742),
.A2(n_439),
.B(n_435),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_793),
.A2(n_350),
.B1(n_425),
.B2(n_423),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_717),
.B(n_21),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_736),
.A2(n_430),
.B(n_425),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_749),
.A2(n_430),
.B(n_423),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_736),
.A2(n_422),
.B(n_421),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_757),
.B(n_422),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_743),
.A2(n_421),
.B(n_419),
.C(n_350),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_790),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_726),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_766),
.A2(n_419),
.B(n_139),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_799),
.A2(n_350),
.B(n_24),
.C(n_25),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_790),
.B(n_22),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_790),
.B(n_735),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_769),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_766),
.A2(n_133),
.B(n_174),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_787),
.B(n_350),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_797),
.A2(n_169),
.B(n_163),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_797),
.A2(n_157),
.B(n_156),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_811),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_743),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_823),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_778),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_784),
.A2(n_153),
.B(n_152),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_784),
.A2(n_151),
.B(n_150),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1027),
.B(n_726),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_856),
.A2(n_784),
.B(n_708),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_845),
.B(n_831),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_862),
.B(n_726),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_972),
.A2(n_823),
.B1(n_814),
.B2(n_708),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_961),
.A2(n_749),
.B(n_760),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_943),
.A2(n_726),
.B1(n_761),
.B2(n_784),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_848),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_869),
.B(n_841),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_861),
.A2(n_804),
.B(n_755),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_848),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_893),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_1016),
.B(n_761),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_943),
.A2(n_761),
.B1(n_787),
.B2(n_754),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_849),
.A2(n_804),
.B(n_755),
.Y(n_1047)
);

INVx3_ASAP7_75t_SL g1048 ( 
.A(n_990),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_872),
.A2(n_754),
.B(n_829),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_878),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_845),
.B(n_761),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_920),
.B(n_740),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_969),
.B(n_787),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_842),
.A2(n_740),
.B(n_841),
.C(n_808),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_917),
.A2(n_829),
.B(n_696),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_871),
.A2(n_829),
.B1(n_820),
.B2(n_841),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_SL g1057 ( 
.A(n_937),
.B(n_989),
.C(n_982),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_935),
.A2(n_746),
.B(n_818),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_989),
.B(n_810),
.C(n_802),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_860),
.A2(n_824),
.B(n_696),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1030),
.B(n_840),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_R g1062 ( 
.A(n_895),
.B(n_836),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_991),
.B(n_840),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_958),
.B(n_817),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_979),
.B(n_817),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_879),
.B(n_896),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_871),
.B(n_696),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_873),
.B(n_837),
.Y(n_1068)
);

AO22x1_ASAP7_75t_L g1069 ( 
.A1(n_982),
.A2(n_807),
.B1(n_832),
.B2(n_837),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_895),
.B(n_800),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_882),
.A2(n_696),
.B(n_824),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_868),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1002),
.B(n_834),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_878),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_SL g1075 ( 
.A1(n_894),
.A2(n_807),
.B1(n_832),
.B2(n_837),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_873),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_885),
.A2(n_696),
.B(n_824),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_847),
.A2(n_824),
.B(n_830),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_909),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1000),
.B(n_908),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_947),
.B(n_801),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_SL g1082 ( 
.A(n_956),
.B(n_802),
.C(n_800),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_898),
.A2(n_824),
.B(n_838),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_950),
.A2(n_815),
.B(n_838),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_843),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_928),
.B(n_815),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_978),
.A2(n_913),
.B(n_850),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_965),
.B(n_834),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_883),
.B(n_801),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_843),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_846),
.B(n_837),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_932),
.A2(n_824),
.B(n_832),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_SL g1093 ( 
.A1(n_851),
.A2(n_824),
.B(n_832),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_909),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_967),
.A2(n_807),
.B(n_148),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_910),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1000),
.B(n_32),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_908),
.B(n_851),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_853),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_864),
.A2(n_34),
.B(n_37),
.C(n_38),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_853),
.B(n_145),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_933),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_933),
.B(n_878),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_38),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1022),
.B(n_39),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_880),
.A2(n_117),
.B(n_114),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_878),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_881),
.A2(n_112),
.B(n_109),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_852),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_952),
.A2(n_107),
.B(n_104),
.Y(n_1110)
);

CKINVDCx14_ASAP7_75t_R g1111 ( 
.A(n_918),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1015),
.A2(n_40),
.B(n_42),
.C(n_46),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1021),
.A2(n_951),
.B1(n_867),
.B2(n_858),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_855),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_887),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_901),
.B(n_92),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_980),
.A2(n_47),
.B(n_48),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_974),
.B(n_50),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1024),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_952),
.A2(n_90),
.B(n_86),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1005),
.A2(n_889),
.B(n_1012),
.C(n_1010),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_879),
.B(n_896),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_888),
.A2(n_84),
.B1(n_81),
.B2(n_62),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_901),
.B(n_60),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_901),
.B(n_61),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_954),
.A2(n_72),
.B(n_64),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_857),
.A2(n_63),
.B(n_68),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_901),
.B(n_69),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_987),
.A2(n_71),
.B1(n_1020),
.B2(n_980),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1015),
.A2(n_956),
.B(n_1029),
.C(n_1028),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_964),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_964),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_977),
.A2(n_886),
.B(n_1007),
.Y(n_1133)
);

OR2x6_ASAP7_75t_SL g1134 ( 
.A(n_981),
.B(n_999),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_921),
.B(n_987),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_859),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_927),
.B(n_865),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_984),
.B(n_1010),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_983),
.Y(n_1139)
);

AND2x4_ASAP7_75t_SL g1140 ( 
.A(n_921),
.B(n_892),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_907),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_892),
.B(n_939),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_939),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_948),
.B(n_960),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_953),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_924),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1029),
.A2(n_1028),
.B(n_1019),
.C(n_891),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_854),
.A2(n_874),
.B(n_995),
.C(n_1004),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_975),
.B(n_953),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_954),
.A2(n_970),
.B(n_912),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_983),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_934),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_970),
.A2(n_844),
.B(n_904),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_905),
.A2(n_931),
.B(n_944),
.Y(n_1155)
);

INVx3_ASAP7_75t_SL g1156 ( 
.A(n_1017),
.Y(n_1156)
);

OAI22x1_ASAP7_75t_L g1157 ( 
.A1(n_924),
.A2(n_911),
.B1(n_1007),
.B2(n_1017),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_863),
.A2(n_866),
.B(n_914),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_891),
.A2(n_994),
.B(n_1013),
.C(n_1011),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_985),
.A2(n_926),
.B(n_875),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_983),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1006),
.A2(n_906),
.B(n_876),
.C(n_916),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1014),
.B(n_897),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1026),
.B(n_1025),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_SL g1166 ( 
.A1(n_897),
.A2(n_1003),
.B(n_988),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1009),
.B(n_915),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_983),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_884),
.A2(n_902),
.B(n_922),
.C(n_890),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_996),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_877),
.B(n_945),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_983),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_899),
.B(n_903),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_923),
.A2(n_1008),
.B(n_929),
.C(n_942),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1009),
.B(n_1001),
.C(n_1018),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_870),
.B(n_986),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_998),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_936),
.B(n_963),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_919),
.A2(n_949),
.B(n_925),
.C(n_993),
.Y(n_1179)
);

NOR2x1p5_ASAP7_75t_L g1180 ( 
.A(n_938),
.B(n_946),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_940),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_971),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_962),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_962),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_962),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_931),
.A2(n_944),
.B1(n_900),
.B2(n_988),
.Y(n_1186)
);

CKINVDCx8_ASAP7_75t_R g1187 ( 
.A(n_962),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1003),
.B(n_976),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_966),
.A2(n_930),
.B(n_941),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_962),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1023),
.Y(n_1191)
);

BUFx2_ASAP7_75t_SL g1192 ( 
.A(n_1044),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1109),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1070),
.A2(n_997),
.B(n_968),
.C(n_973),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1121),
.A2(n_959),
.B1(n_955),
.B2(n_957),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1051),
.B(n_1070),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1138),
.A2(n_1035),
.B(n_1062),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1087),
.A2(n_1042),
.B(n_1047),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1100),
.A2(n_1127),
.B(n_1101),
.C(n_1054),
.Y(n_1199)
);

BUFx2_ASAP7_75t_SL g1200 ( 
.A(n_1090),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1114),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1035),
.B(n_1099),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1168),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1051),
.B(n_1061),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1138),
.B(n_1052),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1034),
.A2(n_1039),
.B(n_1154),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1049),
.A2(n_1171),
.B(n_1060),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1153),
.B(n_1181),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1139),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1149),
.A2(n_1089),
.A3(n_1186),
.B(n_1188),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1068),
.B(n_1041),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1098),
.A2(n_1046),
.B1(n_1033),
.B2(n_1080),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_1188),
.A3(n_1113),
.B(n_1151),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1167),
.A2(n_1166),
.B(n_1171),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1058),
.A2(n_1055),
.B(n_1077),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1071),
.A2(n_1152),
.B(n_1139),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1139),
.A2(n_1152),
.B(n_1165),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1129),
.A2(n_1147),
.B(n_1160),
.C(n_1130),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1037),
.B(n_1134),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1086),
.A2(n_1175),
.B(n_1174),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1139),
.A2(n_1152),
.B(n_1170),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1086),
.A2(n_1150),
.B(n_1064),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1115),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1074),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1152),
.A2(n_1170),
.B(n_1092),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1161),
.A2(n_1133),
.B(n_1155),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1163),
.A2(n_1159),
.B(n_1178),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1191),
.A2(n_1157),
.A3(n_1182),
.B(n_1078),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1068),
.B(n_1045),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1048),
.A2(n_1101),
.B1(n_1128),
.B2(n_1125),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1177),
.B(n_1063),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1168),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1146),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1105),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1085),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1082),
.A2(n_1093),
.B(n_1081),
.C(n_1084),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1111),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1159),
.A2(n_1178),
.B(n_1169),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1143),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_SL g1243 ( 
.A1(n_1104),
.A2(n_1118),
.B(n_1126),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1191),
.A2(n_1083),
.A3(n_1150),
.B(n_1095),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1159),
.A2(n_1176),
.B(n_1179),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1176),
.A2(n_1179),
.B(n_1067),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1116),
.A2(n_1135),
.B(n_1124),
.C(n_1128),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1082),
.A2(n_1164),
.B(n_1059),
.C(n_1112),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1056),
.A2(n_1184),
.A3(n_1106),
.B(n_1108),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1036),
.B(n_1088),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1116),
.A2(n_1124),
.B(n_1125),
.C(n_1103),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1048),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1102),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1173),
.A2(n_1144),
.B(n_1137),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1091),
.B(n_1050),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1076),
.B(n_1180),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1065),
.A2(n_1073),
.B(n_1103),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1105),
.A2(n_1062),
.B1(n_1097),
.B2(n_1119),
.Y(n_1258)
);

AO32x2_ASAP7_75t_L g1259 ( 
.A1(n_1075),
.A2(n_1123),
.A3(n_1183),
.B1(n_1050),
.B2(n_1069),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1045),
.A2(n_1187),
.B1(n_1162),
.B2(n_1172),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1145),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1053),
.A2(n_1120),
.B(n_1110),
.C(n_1136),
.Y(n_1262)
);

AOI221xp5_ASAP7_75t_L g1263 ( 
.A1(n_1119),
.A2(n_1148),
.B1(n_1141),
.B2(n_1043),
.C(n_1040),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1168),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1183),
.A2(n_1168),
.B(n_1122),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1094),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_SL g1267 ( 
.A(n_1074),
.B(n_1190),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1045),
.A2(n_1156),
.B1(n_1096),
.B2(n_1131),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1038),
.A2(n_1132),
.B(n_1066),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_SL g1270 ( 
.A1(n_1107),
.A2(n_1185),
.B(n_1142),
.C(n_1156),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1122),
.A2(n_1140),
.B1(n_1107),
.B2(n_1074),
.Y(n_1271)
);

NAND4xp25_ASAP7_75t_L g1272 ( 
.A(n_1142),
.B(n_463),
.C(n_470),
.D(n_449),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1074),
.B(n_1185),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1070),
.A2(n_705),
.B(n_809),
.C(n_704),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1044),
.B(n_733),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1040),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1051),
.B(n_705),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1057),
.A2(n_705),
.B1(n_845),
.B2(n_559),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1035),
.B(n_705),
.Y(n_1284)
);

NAND3x1_ASAP7_75t_L g1285 ( 
.A(n_1129),
.B(n_463),
.C(n_470),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1121),
.A2(n_1100),
.B(n_1127),
.C(n_1101),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1051),
.B(n_705),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1070),
.A2(n_705),
.B(n_809),
.C(n_704),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1035),
.B(n_869),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1044),
.B(n_733),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1117),
.A2(n_705),
.B(n_704),
.Y(n_1295)
);

AOI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1057),
.A2(n_562),
.B1(n_449),
.B2(n_705),
.C(n_809),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1044),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1168),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1035),
.B(n_869),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1057),
.A2(n_705),
.B1(n_845),
.B2(n_559),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1087),
.A2(n_1154),
.B(n_1179),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_1090),
.Y(n_1305)
);

CKINVDCx9p33_ASAP7_75t_R g1306 ( 
.A(n_1085),
.Y(n_1306)
);

OAI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1117),
.A2(n_705),
.B(n_704),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1044),
.B(n_733),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1033),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1044),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1057),
.A2(n_705),
.B(n_704),
.C(n_950),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1121),
.A2(n_705),
.B1(n_943),
.B2(n_871),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1090),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1176),
.A2(n_1133),
.B(n_1069),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1121),
.A2(n_1100),
.B(n_1127),
.C(n_1101),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1109),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1035),
.B(n_705),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1074),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1057),
.A2(n_705),
.B1(n_895),
.B2(n_1129),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1044),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1109),
.Y(n_1324)
);

AO21x1_ASAP7_75t_L g1325 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1130),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1070),
.A2(n_705),
.B(n_809),
.C(n_704),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1121),
.A2(n_705),
.B(n_785),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1121),
.A2(n_705),
.B1(n_943),
.B2(n_871),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1121),
.A2(n_705),
.B(n_785),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1057),
.A2(n_705),
.B1(n_845),
.B2(n_559),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1168),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1109),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1121),
.A2(n_705),
.B(n_785),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1158),
.A2(n_1161),
.B(n_1189),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1121),
.A2(n_705),
.B1(n_943),
.B2(n_871),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1087),
.A2(n_695),
.B(n_856),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1051),
.B(n_705),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1121),
.A2(n_870),
.A3(n_1087),
.B(n_1149),
.Y(n_1341)
);

AO22x2_ASAP7_75t_L g1342 ( 
.A1(n_1057),
.A2(n_1127),
.B1(n_894),
.B2(n_989),
.Y(n_1342)
);

AOI221x1_ASAP7_75t_L g1343 ( 
.A1(n_1127),
.A2(n_1100),
.B1(n_1121),
.B2(n_1117),
.C(n_989),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1044),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1310),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1201),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_1283),
.B2(n_1332),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1193),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1227),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1298),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1280),
.B(n_1287),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1340),
.B(n_1205),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1306),
.Y(n_1353)
);

INVx6_ASAP7_75t_L g1354 ( 
.A(n_1298),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1266),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1226),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1232),
.B(n_1214),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1277),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1296),
.A2(n_1295),
.B1(n_1307),
.B2(n_1327),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1242),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1322),
.A2(n_1285),
.B1(n_1301),
.B2(n_1289),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1196),
.B(n_1204),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1329),
.A2(n_1336),
.B1(n_1325),
.B2(n_1322),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1305),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1318),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1342),
.A2(n_1258),
.B1(n_1197),
.B2(n_1222),
.Y(n_1366)
);

BUFx2_ASAP7_75t_SL g1367 ( 
.A(n_1261),
.Y(n_1367)
);

INVx3_ASAP7_75t_SL g1368 ( 
.A(n_1236),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1342),
.A2(n_1258),
.B1(n_1272),
.B2(n_1223),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1299),
.A2(n_1288),
.B1(n_1275),
.B2(n_1326),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1324),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1313),
.A2(n_1338),
.B1(n_1328),
.B2(n_1237),
.Y(n_1372)
);

CKINVDCx14_ASAP7_75t_R g1373 ( 
.A(n_1240),
.Y(n_1373)
);

OAI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1202),
.A2(n_1309),
.B1(n_1256),
.B2(n_1334),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1333),
.Y(n_1375)
);

BUFx4f_ASAP7_75t_SL g1376 ( 
.A(n_1323),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1314),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1221),
.A2(n_1312),
.B1(n_1208),
.B2(n_1308),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1237),
.A2(n_1233),
.B1(n_1243),
.B2(n_1217),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1209),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1214),
.B(n_1232),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1344),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1333),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1343),
.A2(n_1234),
.B1(n_1250),
.B2(n_1225),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1213),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1253),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1231),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1276),
.A2(n_1290),
.B1(n_1248),
.B2(n_1239),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1252),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1192),
.A2(n_1200),
.B1(n_1238),
.B2(n_1215),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1263),
.A2(n_1254),
.B1(n_1230),
.B2(n_1241),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1297),
.Y(n_1392)
);

BUFx4_ASAP7_75t_R g1393 ( 
.A(n_1267),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1203),
.B(n_1235),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1268),
.A2(n_1260),
.B1(n_1220),
.B2(n_1224),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1245),
.A2(n_1257),
.B1(n_1286),
.B2(n_1317),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1212),
.B(n_1247),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1227),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1320),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1199),
.A2(n_1251),
.B1(n_1255),
.B2(n_1271),
.Y(n_1400)
);

BUFx8_ASAP7_75t_SL g1401 ( 
.A(n_1320),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1320),
.Y(n_1402)
);

INVxp67_ASAP7_75t_SL g1403 ( 
.A(n_1269),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1231),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1211),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1212),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1211),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1246),
.A2(n_1302),
.B1(n_1218),
.B2(n_1195),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1203),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1235),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1270),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1264),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1302),
.A2(n_1207),
.B1(n_1206),
.B2(n_1198),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1265),
.A2(n_1228),
.B1(n_1259),
.B2(n_1316),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1273),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1274),
.A2(n_1339),
.B1(n_1293),
.B2(n_1291),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1273),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1262),
.A2(n_1255),
.B1(n_1315),
.B2(n_1194),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1259),
.A2(n_1294),
.B1(n_1335),
.B2(n_1321),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1216),
.B(n_1294),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1219),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1216),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1282),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1244),
.Y(n_1425)
);

BUFx2_ASAP7_75t_SL g1426 ( 
.A(n_1304),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1244),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1330),
.A2(n_1331),
.B1(n_1229),
.B2(n_1300),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1249),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1281),
.B(n_1292),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1292),
.B(n_1311),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1341),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1292),
.Y(n_1434)
);

OAI21xp33_ASAP7_75t_L g1435 ( 
.A1(n_1210),
.A2(n_1337),
.B(n_1278),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1249),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1249),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1279),
.A2(n_1303),
.B1(n_1294),
.B2(n_1311),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1311),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_SL g1440 ( 
.A(n_1316),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1316),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1321),
.A2(n_1284),
.B1(n_1319),
.B2(n_705),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1321),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1335),
.A2(n_1284),
.B1(n_1319),
.B2(n_1322),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1335),
.Y(n_1445)
);

INVx3_ASAP7_75t_SL g1446 ( 
.A(n_1341),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_449),
.B2(n_825),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1298),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1266),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1296),
.A2(n_1319),
.B1(n_1284),
.B2(n_1307),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1266),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_705),
.B2(n_1296),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1266),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1284),
.B(n_1319),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1242),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_705),
.B2(n_1296),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1201),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1305),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1298),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_449),
.B2(n_825),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1296),
.A2(n_1319),
.B1(n_1284),
.B2(n_1307),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1298),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1193),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1305),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1284),
.B(n_1319),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1323),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1193),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1296),
.A2(n_562),
.B(n_1283),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1296),
.A2(n_1319),
.B1(n_1284),
.B2(n_1307),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1296),
.A2(n_1319),
.B1(n_1284),
.B2(n_1307),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_1322),
.B2(n_1296),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1193),
.Y(n_1472)
);

CKINVDCx16_ASAP7_75t_R g1473 ( 
.A(n_1305),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1193),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1201),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_SL g1476 ( 
.A(n_1201),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1298),
.B(n_1139),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1193),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1201),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1284),
.A2(n_1319),
.B1(n_1322),
.B2(n_1296),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1434),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1420),
.B(n_1432),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1406),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1382),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1439),
.Y(n_1487)
);

AOI222xp33_ASAP7_75t_L g1488 ( 
.A1(n_1468),
.A2(n_1347),
.B1(n_1471),
.B2(n_1480),
.C1(n_1470),
.C2(n_1469),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1431),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1378),
.B(n_1400),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1380),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1393),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1404),
.Y(n_1493)
);

AOI222xp33_ASAP7_75t_L g1494 ( 
.A1(n_1471),
.A2(n_1480),
.B1(n_1470),
.B2(n_1469),
.C1(n_1450),
.C2(n_1461),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1385),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1362),
.B(n_1452),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1429),
.A2(n_1418),
.B(n_1416),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1447),
.A2(n_1460),
.B1(n_1369),
.B2(n_1461),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1443),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1441),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1440),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1429),
.A2(n_1416),
.B(n_1438),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1386),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1440),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1387),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1454),
.B(n_1465),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1447),
.A2(n_1460),
.B1(n_1369),
.B2(n_1450),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1438),
.A2(n_1435),
.B(n_1437),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1425),
.B(n_1397),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1437),
.A2(n_1396),
.B(n_1391),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1391),
.A2(n_1396),
.B(n_1363),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1422),
.B(n_1419),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1456),
.A2(n_1366),
.B1(n_1359),
.B2(n_1444),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1348),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1417),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1443),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1433),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1417),
.Y(n_1518)
);

AO21x1_ASAP7_75t_L g1519 ( 
.A1(n_1442),
.A2(n_1444),
.B(n_1384),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1403),
.Y(n_1520)
);

INVx4_ASAP7_75t_SL g1521 ( 
.A(n_1446),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1421),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1365),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1403),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1371),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1390),
.A2(n_1388),
.B1(n_1422),
.B2(n_1395),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1384),
.A2(n_1370),
.B(n_1361),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1374),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1422),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1475),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1356),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1428),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1426),
.B(n_1436),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1419),
.B(n_1446),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1345),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1366),
.A2(n_1359),
.B1(n_1363),
.B2(n_1372),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1463),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1436),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1430),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1372),
.A2(n_1423),
.B1(n_1445),
.B2(n_1379),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1421),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1467),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1379),
.A2(n_1414),
.B(n_1408),
.C(n_1474),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1421),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1472),
.B(n_1478),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1408),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1414),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1376),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1355),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1477),
.A2(n_1410),
.B(n_1451),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1358),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1417),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1477),
.A2(n_1449),
.B(n_1453),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1413),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_SL g1556 ( 
.A(n_1476),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1383),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1354),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1413),
.A2(n_1392),
.B(n_1412),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1411),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1411),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1411),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1394),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1409),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1398),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1353),
.B(n_1473),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1375),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1354),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1375),
.A2(n_1462),
.B(n_1381),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1376),
.B(n_1466),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1462),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1357),
.B(n_1455),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1393),
.A2(n_1415),
.B(n_1367),
.C(n_1399),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1373),
.A2(n_1349),
.B1(n_1402),
.B2(n_1389),
.C(n_1457),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1466),
.B(n_1360),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1350),
.A2(n_1448),
.B(n_1405),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1360),
.B(n_1399),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1498),
.A2(n_1373),
.B(n_1377),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1520),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1507),
.A2(n_1368),
.B1(n_1479),
.B2(n_1346),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1483),
.B(n_1350),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1491),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1502),
.A2(n_1407),
.B(n_1459),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1368),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

AO21x1_ASAP7_75t_L g1586 ( 
.A1(n_1492),
.A2(n_1459),
.B(n_1464),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1494),
.A2(n_1488),
.B(n_1490),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1540),
.B(n_1464),
.Y(n_1588)
);

AND2x6_ASAP7_75t_L g1589 ( 
.A(n_1516),
.B(n_1407),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1501),
.B(n_1401),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1490),
.A2(n_1407),
.B(n_1364),
.C(n_1458),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1496),
.B(n_1483),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1506),
.B(n_1535),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1531),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1486),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1519),
.A2(n_1497),
.B(n_1502),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1540),
.B(n_1487),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1544),
.A2(n_1513),
.B(n_1536),
.C(n_1526),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1487),
.B(n_1484),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1556),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1546),
.B(n_1483),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1527),
.A2(n_1511),
.B1(n_1541),
.B2(n_1492),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1510),
.A2(n_1547),
.B(n_1548),
.C(n_1559),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1504),
.B(n_1569),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1510),
.A2(n_1547),
.B(n_1548),
.C(n_1555),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1533),
.B(n_1528),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1546),
.B(n_1563),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1573),
.A2(n_1511),
.B(n_1576),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1504),
.B(n_1569),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1570),
.A2(n_1560),
.B1(n_1561),
.B2(n_1562),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1527),
.A2(n_1555),
.B1(n_1524),
.B2(n_1534),
.C(n_1489),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1565),
.B(n_1495),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1550),
.B(n_1552),
.Y(n_1613)
);

AOI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1527),
.A2(n_1511),
.B(n_1522),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1574),
.A2(n_1511),
.B1(n_1561),
.B2(n_1562),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1530),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1550),
.B(n_1552),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1560),
.A2(n_1554),
.B(n_1551),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1503),
.B(n_1514),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1485),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1534),
.A2(n_1489),
.B1(n_1512),
.B2(n_1549),
.C(n_1525),
.Y(n_1621)
);

AO32x1_ASAP7_75t_L g1622 ( 
.A1(n_1493),
.A2(n_1482),
.A3(n_1485),
.B1(n_1481),
.B2(n_1505),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1508),
.A2(n_1538),
.B(n_1493),
.Y(n_1623)
);

AO21x1_ASAP7_75t_L g1624 ( 
.A1(n_1567),
.A2(n_1571),
.B(n_1564),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1572),
.B(n_1509),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1533),
.B(n_1499),
.Y(n_1626)
);

NOR2xp67_ASAP7_75t_L g1627 ( 
.A(n_1515),
.B(n_1553),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1538),
.A2(n_1532),
.B(n_1517),
.Y(n_1628)
);

AO32x2_ASAP7_75t_L g1629 ( 
.A1(n_1558),
.A2(n_1568),
.A3(n_1515),
.B1(n_1518),
.B2(n_1553),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1587),
.A2(n_1512),
.B1(n_1545),
.B2(n_1522),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1592),
.B(n_1566),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1620),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1604),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1579),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1582),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1585),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1623),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1537),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1604),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1623),
.B(n_1529),
.Y(n_1641)
);

INVx5_ASAP7_75t_L g1642 ( 
.A(n_1626),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1604),
.B(n_1521),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1589),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1482),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1624),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1525),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1523),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.B(n_1500),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1592),
.A2(n_1542),
.B1(n_1522),
.B2(n_1545),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1583),
.B(n_1481),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1622),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1629),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1632),
.Y(n_1657)
);

AOI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1639),
.A2(n_1598),
.B1(n_1580),
.B2(n_1578),
.C(n_1603),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

AOI33xp33_ASAP7_75t_L g1661 ( 
.A1(n_1630),
.A2(n_1602),
.A3(n_1621),
.B1(n_1595),
.B2(n_1588),
.B3(n_1597),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1633),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1656),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1641),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1631),
.B(n_1584),
.Y(n_1665)
);

OAI33xp33_ASAP7_75t_L g1666 ( 
.A1(n_1639),
.A2(n_1593),
.A3(n_1617),
.B1(n_1613),
.B2(n_1601),
.B3(n_1600),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1638),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1647),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1656),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1641),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1645),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1644),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1654),
.Y(n_1676)
);

AO21x2_ASAP7_75t_L g1677 ( 
.A1(n_1648),
.A2(n_1614),
.B(n_1618),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1648),
.A2(n_1598),
.B1(n_1603),
.B2(n_1605),
.C(n_1602),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1654),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1634),
.B(n_1629),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1644),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1610),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1652),
.B(n_1605),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1652),
.B(n_1612),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1678),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1684),
.B(n_1657),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1680),
.B(n_1640),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1683),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1680),
.B(n_1640),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1649),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1672),
.B(n_1651),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1660),
.B(n_1649),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1681),
.B(n_1651),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1674),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1655),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1674),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1662),
.B(n_1650),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1662),
.B(n_1637),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1683),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1702),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1679),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1676),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1688),
.B(n_1679),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1705),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1690),
.B(n_1682),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1702),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1708),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1705),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1707),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1702),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1707),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1701),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1701),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1703),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1688),
.B(n_1676),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.B(n_1682),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1694),
.B(n_1661),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1694),
.B(n_1661),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1695),
.Y(n_1730)
);

AO22x1_ASAP7_75t_L g1731 ( 
.A1(n_1690),
.A2(n_1590),
.B1(n_1600),
.B2(n_1581),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1708),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1695),
.B(n_1682),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1698),
.B(n_1685),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1695),
.B(n_1675),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1706),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1686),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1699),
.B(n_1685),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1616),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1706),
.A2(n_1658),
.B1(n_1630),
.B2(n_1683),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1700),
.B(n_1675),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1704),
.B(n_1658),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1700),
.B(n_1675),
.Y(n_1746)
);

AO22x1_ASAP7_75t_L g1747 ( 
.A1(n_1696),
.A2(n_1590),
.B1(n_1668),
.B2(n_1616),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1692),
.B(n_1669),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1686),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1686),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1599),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1735),
.B(n_1700),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1716),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1670),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1710),
.B(n_1696),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1735),
.B(n_1675),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1732),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1745),
.B(n_1697),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1728),
.B(n_1729),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1740),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1734),
.B(n_1697),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1735),
.B(n_1675),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1740),
.Y(n_1763)
);

AOI31xp33_ASAP7_75t_L g1764 ( 
.A1(n_1743),
.A2(n_1591),
.A3(n_1683),
.B(n_1726),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1749),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1721),
.B(n_1697),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_1659),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1749),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1733),
.B(n_1659),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1709),
.Y(n_1771)
);

NAND2x1p5_ASAP7_75t_L g1772 ( 
.A(n_1738),
.B(n_1646),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1736),
.B(n_1692),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1714),
.B(n_1689),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1721),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1750),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1714),
.B(n_1689),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1742),
.B(n_1666),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1750),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1722),
.B(n_1697),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1741),
.B(n_1693),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1725),
.B(n_1689),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1722),
.B(n_1693),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1725),
.B(n_1689),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1723),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1733),
.B(n_1691),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1723),
.B(n_1693),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1747),
.B(n_1691),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1788),
.B(n_1727),
.Y(n_1789)
);

AO221x1_ASAP7_75t_L g1790 ( 
.A1(n_1766),
.A2(n_1727),
.B1(n_1747),
.B2(n_1719),
.C(n_1715),
.Y(n_1790)
);

OAI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1764),
.A2(n_1615),
.B1(n_1608),
.B2(n_1642),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1752),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1759),
.B(n_1594),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1778),
.A2(n_1666),
.B1(n_1731),
.B2(n_1586),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1759),
.B(n_1751),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1758),
.A2(n_1731),
.B1(n_1677),
.B2(n_1659),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1755),
.A2(n_1591),
.B(n_1566),
.C(n_1575),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1764),
.B(n_1594),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1758),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1760),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1755),
.A2(n_1659),
.B1(n_1671),
.B2(n_1744),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1788),
.A2(n_1677),
.B1(n_1659),
.B2(n_1671),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1772),
.A2(n_1671),
.B1(n_1744),
.B2(n_1642),
.Y(n_1803)
);

OAI322xp33_ASAP7_75t_L g1804 ( 
.A1(n_1753),
.A2(n_1709),
.A3(n_1715),
.B1(n_1719),
.B2(n_1711),
.C1(n_1748),
.C2(n_1739),
.Y(n_1804)
);

NAND2x1_ASAP7_75t_L g1805 ( 
.A(n_1770),
.B(n_1744),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1760),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1763),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1752),
.B(n_1737),
.Y(n_1808)
);

OAI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1754),
.A2(n_1717),
.B(n_1713),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1753),
.B(n_1590),
.Y(n_1810)
);

O2A1O1Ixp5_ASAP7_75t_L g1811 ( 
.A1(n_1757),
.A2(n_1713),
.B(n_1717),
.C(n_1718),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1770),
.B(n_1737),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1772),
.A2(n_1720),
.B(n_1718),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1800),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1805),
.Y(n_1816)
);

O2A1O1Ixp33_ASAP7_75t_L g1817 ( 
.A1(n_1798),
.A2(n_1791),
.B(n_1797),
.C(n_1814),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1799),
.B(n_1757),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1792),
.B(n_1761),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1806),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1798),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1807),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1794),
.A2(n_1772),
.B1(n_1770),
.B2(n_1761),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1789),
.Y(n_1824)
);

NAND4xp25_ASAP7_75t_SL g1825 ( 
.A(n_1796),
.B(n_1777),
.C(n_1774),
.D(n_1784),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1813),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1812),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1791),
.A2(n_1775),
.B(n_1785),
.C(n_1766),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1808),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1790),
.B(n_1766),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1810),
.A2(n_1795),
.B1(n_1793),
.B2(n_1802),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1797),
.A2(n_1785),
.B(n_1780),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1803),
.Y(n_1833)
);

NOR3xp33_ASAP7_75t_L g1834 ( 
.A(n_1809),
.B(n_1780),
.C(n_1767),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1824),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1821),
.B(n_1804),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1829),
.B(n_1801),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1830),
.A2(n_1768),
.B1(n_1677),
.B2(n_1767),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1817),
.A2(n_1811),
.B(n_1787),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1824),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1818),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1818),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1816),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1830),
.A2(n_1811),
.B1(n_1769),
.B2(n_1779),
.C(n_1763),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1826),
.B(n_1774),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1828),
.A2(n_1787),
.B(n_1783),
.C(n_1781),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1839),
.A2(n_1823),
.B(n_1825),
.C(n_1831),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1836),
.B(n_1826),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1844),
.A2(n_1832),
.B1(n_1833),
.B2(n_1827),
.C(n_1816),
.Y(n_1849)
);

NAND4xp25_ASAP7_75t_L g1850 ( 
.A(n_1836),
.B(n_1834),
.C(n_1822),
.D(n_1820),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1846),
.A2(n_1815),
.B1(n_1816),
.B2(n_1819),
.C(n_1779),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1835),
.Y(n_1852)
);

OAI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1838),
.A2(n_1783),
.B1(n_1773),
.B2(n_1781),
.C(n_1769),
.Y(n_1853)
);

NAND4xp75_ASAP7_75t_L g1854 ( 
.A(n_1841),
.B(n_1762),
.C(n_1756),
.D(n_1765),
.Y(n_1854)
);

AOI211xp5_ASAP7_75t_L g1855 ( 
.A1(n_1842),
.A2(n_1773),
.B(n_1762),
.C(n_1756),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1848),
.Y(n_1856)
);

NAND4xp75_ASAP7_75t_L g1857 ( 
.A(n_1849),
.B(n_1840),
.C(n_1843),
.D(n_1845),
.Y(n_1857)
);

OAI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1847),
.A2(n_1837),
.B1(n_1765),
.B2(n_1776),
.C(n_1771),
.Y(n_1858)
);

NAND4xp25_ASAP7_75t_L g1859 ( 
.A(n_1850),
.B(n_1837),
.C(n_1776),
.D(n_1771),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1854),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1860),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1858),
.A2(n_1851),
.B(n_1852),
.C(n_1853),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1856),
.B(n_1768),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1859),
.A2(n_1855),
.B1(n_1771),
.B2(n_1768),
.C(n_1782),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1857),
.A2(n_1768),
.B1(n_1784),
.B2(n_1782),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1860),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_SL g1867 ( 
.A(n_1861),
.B(n_1518),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1861),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1863),
.B(n_1777),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1862),
.B(n_1786),
.C(n_1577),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1866),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1869),
.B(n_1865),
.Y(n_1872)
);

NOR3xp33_ASAP7_75t_L g1873 ( 
.A(n_1871),
.B(n_1864),
.C(n_1786),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1868),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1874),
.Y(n_1875)
);

AO22x2_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1872),
.B1(n_1873),
.B2(n_1870),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1876),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1876),
.B(n_1875),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1877),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1878),
.A2(n_1867),
.B(n_1720),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1879),
.A2(n_1711),
.B(n_1724),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1880),
.A2(n_1748),
.B(n_1739),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1881),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1882),
.B(n_1724),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1884),
.Y(n_1885)
);

OAI221xp5_ASAP7_75t_R g1886 ( 
.A1(n_1885),
.A2(n_1744),
.B1(n_1653),
.B2(n_1746),
.C(n_1668),
.Y(n_1886)
);

AOI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_1627),
.B(n_1557),
.C(n_1558),
.Y(n_1887)
);


endmodule