module fake_jpeg_26818_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_16),
.Y(n_54)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_55),
.B1(n_60),
.B2(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_18),
.B1(n_25),
.B2(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_31),
.A2(n_36),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_28),
.B1(n_30),
.B2(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_83),
.B1(n_33),
.B2(n_46),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_40),
.C(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_71),
.B1(n_78),
.B2(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_79),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_77),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_40),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_47),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_51),
.B1(n_56),
.B2(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_26),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_19),
.C(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_27),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_37),
.C(n_17),
.Y(n_81)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_17),
.A3(n_21),
.B1(n_29),
.B2(n_51),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_33),
.B1(n_16),
.B2(n_19),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_59),
.B(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_28),
.B(n_30),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_71),
.B1(n_78),
.B2(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_46),
.B1(n_49),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_78),
.B1(n_68),
.B2(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_102),
.B1(n_105),
.B2(n_83),
.Y(n_114)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_23),
.B(n_24),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_23),
.B(n_24),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_80),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_76),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_69),
.C(n_66),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_17),
.C(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_100),
.B1(n_93),
.B2(n_99),
.Y(n_135)
);

OAI21x1_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_81),
.B(n_75),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_93),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_90),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_127),
.B1(n_103),
.B2(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_67),
.B(n_62),
.C(n_65),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_95),
.B(n_105),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_63),
.B1(n_62),
.B2(n_23),
.Y(n_123)
);

OAI22x1_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_128),
.B1(n_17),
.B2(n_21),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_26),
.B1(n_81),
.B2(n_29),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_101),
.B1(n_86),
.B2(n_89),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_135),
.B1(n_120),
.B2(n_127),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_140),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_141),
.B(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_95),
.B1(n_98),
.B2(n_91),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_104),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_82),
.B(n_21),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_108),
.B1(n_125),
.B2(n_117),
.Y(n_161)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_112),
.B1(n_16),
.B2(n_19),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_106),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_103),
.B(n_21),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_19),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_21),
.B(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_165),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_157),
.A2(n_159),
.B1(n_166),
.B2(n_138),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_133),
.B(n_143),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_139),
.C(n_7),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_147),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_118),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_20),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_20),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_148),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_170),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_135),
.A3(n_136),
.B1(n_150),
.B2(n_146),
.C1(n_141),
.C2(n_145),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_168),
.B(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_150),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.C(n_185),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_151),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_151),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_155),
.B(n_153),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_5),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_152),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_188),
.B(n_192),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_155),
.B(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_197),
.B1(n_5),
.B2(n_13),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_199),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_5),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_192),
.B1(n_194),
.B2(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_182),
.B1(n_176),
.B2(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_183),
.C(n_173),
.Y(n_201)
);

OAI211xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_3),
.B(n_10),
.C(n_14),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_4),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_195),
.C(n_196),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_4),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_210),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_9),
.B(n_13),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_202),
.B(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_200),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_3),
.C(n_10),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_208),
.C(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_215),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_213),
.B(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_0),
.C(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_0),
.Y(n_224)
);


endmodule