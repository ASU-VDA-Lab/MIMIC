module fake_jpeg_5732_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx12_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_4),
.A3(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_14),
.A2(n_18),
.B1(n_15),
.B2(n_24),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_21),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_28),
.B(n_24),
.C(n_25),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_32),
.B2(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_30),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_21),
.A3(n_22),
.B1(n_25),
.B2(n_28),
.C1(n_29),
.C2(n_34),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_22),
.CI(n_35),
.CON(n_37),
.SN(n_37)
);


endmodule