module fake_jpeg_26942_n_43 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_43);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_8),
.B1(n_13),
.B2(n_11),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_0),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_9),
.B1(n_14),
.B2(n_4),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_18),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.C(n_31),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_20),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_1),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_23),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_36),
.C(n_21),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_21),
.C(n_18),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B1(n_27),
.B2(n_2),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_21),
.B(n_2),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_1),
.B(n_4),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_35),
.B(n_6),
.Y(n_43)
);


endmodule