module fake_jpeg_2114_n_328 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_47),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_27),
.B2(n_33),
.Y(n_60)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

OR2x4_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_20),
.Y(n_59)
);

NOR2x1_ASAP7_75t_R g113 ( 
.A(n_59),
.B(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_23),
.B1(n_34),
.B2(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_72),
.B1(n_18),
.B2(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_32),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_15),
.B1(n_28),
.B2(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_15),
.B1(n_28),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_63),
.B1(n_18),
.B2(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_33),
.B1(n_27),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_46),
.B1(n_33),
.B2(n_49),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_16),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_53),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_81),
.B(n_86),
.Y(n_153)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_44),
.B1(n_41),
.B2(n_45),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_104),
.Y(n_132)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_91),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_22),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_46),
.B(n_17),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_20),
.B(n_26),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_95),
.B(n_107),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_106),
.Y(n_152)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_103),
.B1(n_26),
.B2(n_1),
.Y(n_151)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_17),
.B1(n_25),
.B2(n_22),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_112),
.B1(n_118),
.B2(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_117),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_24),
.B1(n_33),
.B2(n_48),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_39),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_24),
.B1(n_33),
.B2(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_51),
.C(n_37),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_20),
.C(n_77),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_57),
.B1(n_31),
.B2(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_76),
.B(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_124),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_29),
.B1(n_28),
.B2(n_18),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_20),
.B1(n_26),
.B2(n_2),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_18),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_20),
.A3(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_128),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_20),
.C(n_77),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_120),
.C(n_129),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_151),
.B1(n_100),
.B2(n_97),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_145),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_125),
.B1(n_127),
.B2(n_126),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_96),
.B1(n_92),
.B2(n_94),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_83),
.B1(n_116),
.B2(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_171),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_178),
.B1(n_184),
.B2(n_190),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_116),
.B1(n_94),
.B2(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_104),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_96),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_82),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_182),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_106),
.B1(n_115),
.B2(n_114),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_146),
.B1(n_156),
.B2(n_142),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_109),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_181),
.Y(n_203)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_111),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_85),
.B1(n_89),
.B2(n_26),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_189),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_149),
.B(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_188),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_0),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_159),
.B1(n_155),
.B2(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_12),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_154),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_134),
.B1(n_131),
.B2(n_148),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_136),
.C(n_137),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_198),
.C(n_204),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_161),
.C(n_152),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_152),
.A3(n_145),
.B1(n_144),
.B2(n_150),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_152),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_178),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_217),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_150),
.C(n_144),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_156),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_190),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_138),
.B1(n_134),
.B2(n_142),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_184),
.B1(n_186),
.B2(n_188),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_154),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_179),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_148),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_168),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_240),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_165),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_239),
.B1(n_241),
.B2(n_207),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_165),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_188),
.B1(n_165),
.B2(n_192),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_131),
.A3(n_140),
.B1(n_180),
.B2(n_133),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_243),
.B(n_206),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_140),
.B(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_195),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_242),
.C(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_213),
.B1(n_196),
.B2(n_197),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_241),
.A2(n_207),
.B1(n_203),
.B2(n_220),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_259),
.B1(n_261),
.B2(n_264),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_194),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_205),
.B1(n_212),
.B2(n_209),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_214),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_205),
.B1(n_201),
.B2(n_133),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_238),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_265),
.B(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_222),
.C(n_223),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_277),
.C(n_269),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_253),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_239),
.B1(n_235),
.B2(n_221),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_281),
.B1(n_254),
.B2(n_261),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_227),
.C(n_237),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_10),
.B1(n_1),
.B2(n_3),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_264),
.B(n_246),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_0),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_247),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_292),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_280),
.C(n_267),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_245),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_297),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_267),
.B(n_270),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_267),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_284),
.C(n_291),
.Y(n_300)
);

OAI321xp33_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_293),
.C(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_309),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_293),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_296),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_283),
.C(n_5),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_4),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_298),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_305),
.B1(n_297),
.B2(n_299),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_317),
.B(n_319),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_307),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_5),
.B(n_7),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_5),
.C(n_8),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_308),
.B1(n_311),
.B2(n_309),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_322),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_316),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_319),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.C(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_314),
.Y(n_328)
);


endmodule