module fake_jpeg_1214_n_56 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_56);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_20),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_15),
.B1(n_13),
.B2(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_23),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_21),
.B(n_22),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_25),
.B(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_24),
.C(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_25),
.B1(n_38),
.B2(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_19),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_16),
.B(n_17),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_42),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_25),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_16),
.C(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_7),
.C(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_4),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_3),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_50),
.B(n_53),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_51),
.B(n_53),
.C(n_6),
.Y(n_56)
);


endmodule