module fake_jpeg_12912_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_3),
.Y(n_7)
);

OR2x2_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_3),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

OR2x2_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_22),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_6),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_13),
.C(n_20),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_39),
.B1(n_32),
.B2(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_17),
.B1(n_19),
.B2(n_35),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_31),
.B(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_31),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_45),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_44),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_48),
.Y(n_52)
);


endmodule