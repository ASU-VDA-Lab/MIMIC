module fake_netlist_6_4253_n_1553 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1553);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1553;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_47),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_43),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_52),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_37),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_0),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g154 ( 
.A(n_44),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_53),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_30),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_40),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_50),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_11),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_50),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_60),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_28),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_36),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_42),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_51),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_44),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_52),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_69),
.Y(n_181)
);

BUFx8_ASAP7_75t_SL g182 ( 
.A(n_141),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_12),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_26),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_23),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_9),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_41),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_57),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_105),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_112),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_41),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_47),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_17),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_18),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_35),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_20),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_27),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_73),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_30),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_3),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_34),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_82),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_20),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_102),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_84),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_14),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_122),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_58),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_18),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_78),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_129),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_71),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_97),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_16),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_111),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_24),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_7),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_74),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_143),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_38),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_64),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_85),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_77),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_49),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_119),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_76),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_118),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_1),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_65),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_80),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_108),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_81),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_35),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_93),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_135),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_107),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_15),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_149),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_250),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_182),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_146),
.B(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_149),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_2),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_149),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_179),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_174),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_181),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_174),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_174),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_193),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_188),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_145),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_192),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_174),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_284),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_199),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_201),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_237),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_202),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_147),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_171),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_203),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_187),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_187),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_218),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_237),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_205),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_226),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_228),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_229),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_232),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_234),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_176),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_151),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_205),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_238),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_242),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_154),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_148),
.B(n_6),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_153),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_158),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_160),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_164),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_248),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_251),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_154),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_189),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_253),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_175),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_148),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_196),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_346),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_196),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_317),
.B(n_169),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_298),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_294),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_292),
.B(n_360),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_297),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_173),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_299),
.B(n_204),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_299),
.B(n_204),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_302),
.B(n_256),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_301),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_306),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_290),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_309),
.B(n_256),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_308),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_309),
.B(n_274),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_310),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_311),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_315),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_330),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_331),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_274),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_336),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_337),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_295),
.B(n_190),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_344),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_322),
.B(n_173),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_355),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_357),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_304),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_328),
.B(n_184),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_329),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_325),
.B(n_144),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_400),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_414),
.A2(n_279),
.B1(n_206),
.B2(n_233),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_423),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_364),
.B(n_356),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_373),
.B(n_166),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_184),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_321),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

NAND2x1p5_ASAP7_75t_L g445 ( 
.A(n_380),
.B(n_152),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_400),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_327),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_183),
.C(n_180),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_373),
.B(n_334),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_386),
.B(n_335),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g452 ( 
.A(n_381),
.B(n_273),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_273),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_207),
.B1(n_266),
.B2(n_258),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_361),
.B(n_353),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_387),
.B(n_338),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_361),
.B(n_353),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_397),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_329),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_390),
.B(n_190),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_400),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_342),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_388),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_178),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_393),
.A2(n_359),
.B1(n_305),
.B2(n_300),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_144),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_375),
.B(n_163),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_361),
.B(n_358),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_414),
.A2(n_190),
.B1(n_198),
.B2(n_209),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_L g479 ( 
.A(n_428),
.B(n_191),
.C(n_185),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_414),
.A2(n_209),
.B1(n_198),
.B2(n_358),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_395),
.B(n_150),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_379),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_414),
.A2(n_366),
.B1(n_363),
.B2(n_381),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_363),
.A2(n_209),
.B1(n_198),
.B2(n_354),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_381),
.B(n_392),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_378),
.Y(n_496)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_396),
.B(n_288),
.C(n_223),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_402),
.B(n_159),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_404),
.A2(n_159),
.B1(n_286),
.B2(n_285),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_366),
.B(n_236),
.C(n_200),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_381),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_381),
.A2(n_209),
.B1(n_198),
.B2(n_354),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_416),
.B(n_333),
.Y(n_506)
);

NOR2x1p5_ASAP7_75t_L g507 ( 
.A(n_405),
.B(n_151),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_388),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_392),
.B(n_186),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_426),
.A2(n_208),
.B1(n_211),
.B2(n_210),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_333),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_408),
.B(n_165),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_364),
.B(n_169),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_423),
.B(n_341),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_409),
.B(n_165),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_415),
.B(n_417),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_384),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_411),
.B(n_348),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_418),
.B(n_216),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_369),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_411),
.B(n_167),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_412),
.A2(n_220),
.B1(n_240),
.B2(n_168),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_412),
.B(n_167),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_376),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_376),
.B(n_169),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_399),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_418),
.B(n_222),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_382),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_413),
.B(n_170),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_403),
.B(n_212),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_380),
.B(n_209),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_368),
.B(n_293),
.Y(n_535)
);

BUFx4f_ASAP7_75t_L g536 ( 
.A(n_406),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_413),
.B(n_421),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_369),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_369),
.B(n_224),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_369),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_383),
.B(n_293),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_401),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_401),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_401),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_425),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_427),
.B(n_348),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_383),
.B(n_170),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_407),
.B(n_222),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_425),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_429),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_435),
.B(n_225),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_435),
.B(n_227),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_230),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_452),
.B(n_231),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_452),
.A2(n_265),
.B1(n_246),
.B2(n_262),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_495),
.B(n_241),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_541),
.A2(n_470),
.B1(n_475),
.B2(n_544),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_495),
.B(n_264),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_495),
.B(n_267),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_259),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_432),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_537),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_544),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_460),
.B(n_260),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_489),
.B(n_550),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_503),
.B(n_281),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_439),
.A2(n_278),
.B1(n_260),
.B2(n_263),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_436),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_517),
.B(n_410),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_434),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_517),
.B(n_410),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_526),
.B(n_419),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_526),
.B(n_419),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_524),
.B(n_341),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_545),
.B(n_419),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_511),
.B(n_343),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_488),
.B(n_263),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_474),
.B(n_486),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_462),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_509),
.A2(n_347),
.B(n_345),
.C(n_343),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_438),
.A2(n_269),
.B1(n_272),
.B2(n_278),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_500),
.B(n_272),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_511),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_440),
.Y(n_599)
);

BUFx8_ASAP7_75t_L g600 ( 
.A(n_447),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_462),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_506),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_514),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_478),
.A2(n_482),
.B1(n_430),
.B2(n_456),
.Y(n_605)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_439),
.A2(n_168),
.B1(n_172),
.B2(n_162),
.C(n_155),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_422),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_471),
.B(n_472),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_213),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_447),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_512),
.B(n_214),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_524),
.B(n_280),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_518),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_472),
.B(n_215),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_515),
.B(n_219),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g617 ( 
.A(n_473),
.B(n_501),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_536),
.B(n_280),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_449),
.B(n_221),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_479),
.B(n_235),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_441),
.A2(n_280),
.B1(n_249),
.B2(n_245),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_549),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_502),
.B(n_243),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_476),
.B(n_254),
.Y(n_624)
);

AND2x6_ASAP7_75t_SL g625 ( 
.A(n_451),
.B(n_287),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_481),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_476),
.B(n_255),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_525),
.B(n_239),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_441),
.A2(n_244),
.B1(n_283),
.B2(n_277),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_480),
.B(n_155),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_480),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_536),
.B(n_156),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_528),
.B(n_156),
.C(n_283),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_444),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_483),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_536),
.B(n_157),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_483),
.B(n_157),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_441),
.A2(n_261),
.B1(n_277),
.B2(n_275),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_507),
.B(n_161),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_485),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_481),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_446),
.B(n_162),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_493),
.B(n_172),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_496),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_441),
.A2(n_275),
.B1(n_271),
.B2(n_287),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_466),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_431),
.B(n_287),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_441),
.A2(n_195),
.B1(n_154),
.B2(n_66),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_457),
.B(n_62),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_432),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_521),
.B(n_195),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_469),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_431),
.B(n_8),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_546),
.B(n_55),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_455),
.A2(n_140),
.B1(n_139),
.B2(n_130),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_455),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_L g659 ( 
.A(n_535),
.B(n_10),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_432),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_445),
.B(n_106),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_522),
.B(n_13),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_443),
.B(n_95),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_458),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_457),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_432),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_523),
.B(n_13),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_531),
.B(n_15),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_520),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_455),
.A2(n_90),
.B1(n_89),
.B2(n_88),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_445),
.B(n_86),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_508),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_522),
.B(n_19),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_459),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_455),
.A2(n_75),
.B1(n_68),
.B2(n_25),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_459),
.B(n_54),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_513),
.B(n_19),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_455),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_477),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_464),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_583),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_610),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_557),
.B(n_467),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_626),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_654),
.Y(n_685)
);

AO22x1_ASAP7_75t_L g686 ( 
.A1(n_662),
.A2(n_497),
.B1(n_510),
.B2(n_455),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_559),
.A2(n_548),
.B(n_547),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_592),
.B(n_437),
.C(n_516),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_569),
.B(n_507),
.Y(n_689)
);

O2A1O1Ixp5_ASAP7_75t_L g690 ( 
.A1(n_667),
.A2(n_551),
.B(n_533),
.C(n_539),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_653),
.A2(n_477),
.B(n_542),
.C(n_540),
.Y(n_691)
);

AO21x1_ASAP7_75t_L g692 ( 
.A1(n_667),
.A2(n_445),
.B(n_477),
.Y(n_692)
);

BUFx4f_ASAP7_75t_L g693 ( 
.A(n_588),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_561),
.A2(n_491),
.B1(n_504),
.B2(n_540),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_561),
.A2(n_543),
.B1(n_542),
.B2(n_538),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_583),
.Y(n_697)
);

BUFx12f_ASAP7_75t_L g698 ( 
.A(n_600),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_565),
.B(n_592),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_598),
.B(n_519),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_578),
.A2(n_494),
.B(n_453),
.Y(n_701)
);

BUFx8_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_570),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_652),
.A2(n_454),
.B(n_453),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_666),
.A2(n_454),
.B(n_453),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_668),
.A2(n_487),
.B(n_530),
.C(n_527),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_653),
.A2(n_461),
.B(n_492),
.C(n_498),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_597),
.B(n_520),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_562),
.B(n_573),
.Y(n_709)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_612),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_611),
.B(n_492),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_608),
.B(n_484),
.Y(n_712)
);

BUFx8_ASAP7_75t_SL g713 ( 
.A(n_664),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_554),
.B(n_498),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_611),
.B(n_29),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_616),
.A2(n_463),
.B1(n_534),
.B2(n_468),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_651),
.B(n_499),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_553),
.B(n_505),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_642),
.B(n_505),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_616),
.B(n_568),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_600),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_568),
.B(n_29),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_648),
.B(n_490),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_668),
.A2(n_464),
.B(n_463),
.C(n_534),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_582),
.A2(n_463),
.B(n_534),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_584),
.A2(n_463),
.B(n_534),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_586),
.A2(n_463),
.B(n_534),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_619),
.A2(n_463),
.B(n_534),
.C(n_33),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_567),
.A2(n_463),
.B(n_534),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_587),
.A2(n_31),
.B(n_32),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_606),
.B(n_32),
.C(n_33),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_589),
.A2(n_38),
.B(n_45),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_643),
.B(n_45),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_636),
.B(n_641),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_605),
.A2(n_46),
.B1(n_48),
.B2(n_679),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_583),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_660),
.A2(n_46),
.B(n_48),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_643),
.B(n_613),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_660),
.A2(n_555),
.B(n_556),
.Y(n_740)
);

O2A1O1Ixp5_ASAP7_75t_L g741 ( 
.A1(n_618),
.A2(n_579),
.B(n_563),
.C(n_566),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_672),
.B(n_576),
.Y(n_742)
);

O2A1O1Ixp5_ASAP7_75t_L g743 ( 
.A1(n_618),
.A2(n_579),
.B(n_563),
.C(n_566),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_644),
.B(n_646),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_576),
.B(n_591),
.C(n_677),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_614),
.B(n_622),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_651),
.A2(n_679),
.B1(n_617),
.B2(n_665),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_649),
.Y(n_748)
);

NAND2x1_ASAP7_75t_L g749 ( 
.A(n_660),
.B(n_680),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_628),
.B(n_593),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_601),
.B(n_602),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_591),
.B(n_677),
.C(n_619),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_656),
.A2(n_661),
.B(n_671),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_552),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_603),
.B(n_604),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_588),
.B(n_629),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_607),
.B(n_680),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_560),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_590),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_574),
.B(n_585),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_590),
.B(n_629),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_564),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_674),
.B(n_575),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_661),
.A2(n_671),
.B(n_663),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_631),
.B(n_638),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_673),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_659),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_645),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_609),
.B(n_627),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_615),
.B(n_624),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_650),
.B(n_657),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_599),
.B(n_635),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_676),
.B(n_647),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_623),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_620),
.A2(n_623),
.B(n_637),
.C(n_633),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_633),
.A2(n_637),
.B(n_595),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_658),
.A2(n_580),
.B1(n_621),
.B2(n_639),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_670),
.A2(n_675),
.B(n_596),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_630),
.B(n_678),
.Y(n_780)
);

NAND2x1_ASAP7_75t_L g781 ( 
.A(n_634),
.B(n_640),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_625),
.A2(n_571),
.B(n_495),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_577),
.A2(n_559),
.B(n_558),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_571),
.A2(n_495),
.B(n_669),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_571),
.A2(n_495),
.B(n_669),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_577),
.A2(n_559),
.B(n_558),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_577),
.B(n_529),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_653),
.A2(n_577),
.B(n_667),
.C(n_668),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_571),
.A2(n_495),
.B(n_669),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_592),
.B(n_529),
.Y(n_790)
);

AO21x1_ASAP7_75t_L g791 ( 
.A1(n_667),
.A2(n_668),
.B(n_577),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_565),
.B(n_592),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_653),
.A2(n_577),
.B(n_667),
.C(n_668),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_592),
.B(n_450),
.C(n_557),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_667),
.A2(n_668),
.B(n_577),
.C(n_618),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_592),
.B(n_450),
.C(n_557),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_577),
.A2(n_561),
.B1(n_592),
.B2(n_558),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_667),
.A2(n_668),
.B(n_565),
.C(n_577),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_653),
.A2(n_577),
.B(n_667),
.C(n_668),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_557),
.B(n_594),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_557),
.B(n_594),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_577),
.B(n_529),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_577),
.B(n_529),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_577),
.B(n_529),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_577),
.A2(n_592),
.B1(n_565),
.B2(n_611),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_583),
.Y(n_806)
);

OAI321xp33_ASAP7_75t_L g807 ( 
.A1(n_667),
.A2(n_668),
.A3(n_606),
.B1(n_677),
.B2(n_653),
.C(n_658),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_557),
.B(n_594),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_610),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_583),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_610),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_685),
.Y(n_812)
);

AOI21xp33_ASAP7_75t_L g813 ( 
.A1(n_721),
.A2(n_775),
.B(n_752),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_807),
.A2(n_715),
.B(n_805),
.C(n_723),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_783),
.A2(n_786),
.B(n_753),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_790),
.B(n_766),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_810),
.B(n_681),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_788),
.A2(n_799),
.B(n_793),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_694),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_776),
.B(n_798),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_797),
.A2(n_745),
.B(n_787),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_802),
.B(n_803),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_740),
.A2(n_764),
.B(n_708),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_804),
.B(n_770),
.Y(n_824)
);

AOI21x1_ASAP7_75t_SL g825 ( 
.A1(n_774),
.A2(n_780),
.B(n_771),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_800),
.B(n_683),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_718),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_784),
.A2(n_789),
.B(n_785),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_SL g829 ( 
.A(n_794),
.B(n_796),
.C(n_792),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_767),
.B(n_742),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_769),
.B(n_684),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_718),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_809),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_681),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_682),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_741),
.A2(n_743),
.B(n_774),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_699),
.B(n_688),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_691),
.A2(n_777),
.B(n_707),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_687),
.A2(n_711),
.B(n_712),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_718),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_739),
.B(n_801),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_808),
.B(n_761),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_749),
.A2(n_719),
.B(n_712),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_701),
.A2(n_705),
.B(n_704),
.Y(n_844)
);

BUFx4_ASAP7_75t_SL g845 ( 
.A(n_722),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_779),
.A2(n_778),
.B(n_756),
.C(n_734),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_690),
.A2(n_725),
.B(n_696),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_747),
.A2(n_780),
.B1(n_744),
.B2(n_735),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_735),
.B(n_744),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_698),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_763),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_757),
.A2(n_706),
.B(n_726),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_730),
.A2(n_695),
.B(n_727),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_728),
.A2(n_716),
.B(n_763),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_703),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_811),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_746),
.A2(n_709),
.B1(n_750),
.B2(n_751),
.Y(n_857)
);

AO21x1_ASAP7_75t_L g858 ( 
.A1(n_736),
.A2(n_731),
.B(n_733),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_746),
.B(n_709),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_717),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_750),
.B(n_751),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_759),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_732),
.A2(n_755),
.B(n_729),
.C(n_693),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_748),
.B(n_710),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_755),
.B(n_718),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_759),
.B(n_754),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_759),
.B(n_754),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_754),
.A2(n_693),
.B1(n_760),
.B2(n_806),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_692),
.A2(n_700),
.B(n_773),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_737),
.Y(n_870)
);

OA22x2_ASAP7_75t_L g871 ( 
.A1(n_689),
.A2(n_781),
.B1(n_724),
.B2(n_714),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_765),
.Y(n_872)
);

AOI221xp5_ASAP7_75t_SL g873 ( 
.A1(n_782),
.A2(n_738),
.B1(n_720),
.B2(n_758),
.C(n_762),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_686),
.B(n_791),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_681),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_737),
.A2(n_689),
.B(n_772),
.C(n_806),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_772),
.B(n_697),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_772),
.A2(n_697),
.B(n_806),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_697),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_772),
.A2(n_689),
.B(n_702),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_772),
.B(n_702),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_768),
.A2(n_786),
.B(n_783),
.Y(n_882)
);

BUFx2_ASAP7_75t_SL g883 ( 
.A(n_713),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_768),
.B(n_721),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_721),
.B(n_790),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_775),
.B(n_770),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_783),
.A2(n_786),
.B(n_753),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_790),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_783),
.A2(n_786),
.B(n_753),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_721),
.B(n_790),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_800),
.B(n_683),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_721),
.B(n_790),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_694),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_775),
.B(n_721),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_721),
.B(n_790),
.Y(n_895)
);

AND2x6_ASAP7_75t_L g896 ( 
.A(n_775),
.B(n_770),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_783),
.A2(n_786),
.B(n_753),
.Y(n_897)
);

OAI22x1_ASAP7_75t_L g898 ( 
.A1(n_721),
.A2(n_522),
.B1(n_673),
.B2(n_662),
.Y(n_898)
);

AOI21x1_ASAP7_75t_SL g899 ( 
.A1(n_775),
.A2(n_774),
.B(n_780),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_788),
.A2(n_799),
.B(n_793),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_694),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_681),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_783),
.A2(n_786),
.B(n_753),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_721),
.B(n_790),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_759),
.B(n_754),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_759),
.B(n_754),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_718),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_721),
.B(n_790),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_721),
.B(n_790),
.Y(n_909)
);

AND3x2_ASAP7_75t_L g910 ( 
.A(n_721),
.B(n_612),
.C(n_715),
.Y(n_910)
);

O2A1O1Ixp5_ASAP7_75t_L g911 ( 
.A1(n_788),
.A2(n_793),
.B(n_799),
.C(n_721),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_721),
.B(n_790),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_721),
.B(n_790),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_788),
.A2(n_799),
.B(n_793),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_721),
.B(n_790),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_800),
.B(n_683),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_759),
.B(n_754),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_759),
.B(n_754),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_810),
.B(n_681),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_713),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_775),
.B(n_721),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_810),
.B(n_681),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_721),
.B(n_790),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_835),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_881),
.B(n_876),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_812),
.Y(n_926)
);

OA22x2_ASAP7_75t_L g927 ( 
.A1(n_910),
.A2(n_898),
.B1(n_841),
.B2(n_842),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_827),
.B(n_832),
.Y(n_928)
);

CKINVDCx6p67_ASAP7_75t_R g929 ( 
.A(n_850),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_885),
.B(n_888),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_883),
.Y(n_931)
);

OR2x6_ASAP7_75t_SL g932 ( 
.A(n_884),
.B(n_868),
.Y(n_932)
);

INVx8_ASAP7_75t_L g933 ( 
.A(n_875),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_890),
.B(n_892),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_826),
.B(n_891),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_845),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_835),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_870),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_916),
.B(n_830),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_815),
.A2(n_889),
.B(n_887),
.Y(n_940)
);

CKINVDCx6p67_ASAP7_75t_R g941 ( 
.A(n_920),
.Y(n_941)
);

INVx3_ASAP7_75t_SL g942 ( 
.A(n_864),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_814),
.A2(n_911),
.B(n_900),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_895),
.B(n_904),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_860),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_862),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_881),
.B(n_877),
.Y(n_947)
);

AOI21xp33_ASAP7_75t_L g948 ( 
.A1(n_814),
.A2(n_914),
.B(n_818),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_816),
.B(n_894),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_908),
.B(n_909),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_870),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_866),
.B(n_867),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_829),
.A2(n_813),
.B1(n_837),
.B2(n_894),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_833),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_855),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_912),
.B(n_913),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_897),
.A2(n_903),
.B(n_828),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_827),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_897),
.A2(n_903),
.B(n_828),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_856),
.Y(n_960)
);

OR2x2_ASAP7_75t_SL g961 ( 
.A(n_829),
.B(n_915),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_833),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_856),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_866),
.B(n_867),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_876),
.B(n_905),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_831),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_921),
.B(n_923),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_921),
.B(n_911),
.C(n_846),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_882),
.A2(n_824),
.B(n_821),
.C(n_820),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_905),
.B(n_906),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_863),
.A2(n_848),
.B(n_857),
.C(n_861),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_910),
.A2(n_886),
.B1(n_896),
.B2(n_858),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_859),
.B(n_849),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_862),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_906),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_863),
.A2(n_882),
.B(n_822),
.C(n_874),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_917),
.B(n_918),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_851),
.A2(n_827),
.B1(n_840),
.B2(n_907),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_917),
.B(n_918),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_879),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_839),
.A2(n_823),
.B(n_838),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_845),
.Y(n_982)
);

INVx3_ASAP7_75t_SL g983 ( 
.A(n_871),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_832),
.B(n_840),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_875),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_872),
.B(n_893),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_875),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_875),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_865),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_819),
.B(n_901),
.Y(n_990)
);

CKINVDCx8_ASAP7_75t_R g991 ( 
.A(n_886),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_886),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_834),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_886),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_880),
.B(n_834),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_832),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_836),
.A2(n_853),
.B(n_847),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_902),
.B(n_840),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_902),
.B(n_840),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_817),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_853),
.A2(n_852),
.B(n_854),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_832),
.B(n_907),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_873),
.B(n_896),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_896),
.B(n_869),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_896),
.B(n_878),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_907),
.B(n_919),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_922),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_907),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_843),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_825),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_825),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_899),
.B(n_844),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_814),
.A2(n_721),
.B1(n_888),
.B2(n_885),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_814),
.A2(n_911),
.B(n_900),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_812),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_860),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_885),
.B(n_888),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_881),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_815),
.A2(n_889),
.B(n_887),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_826),
.B(n_891),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_885),
.B(n_888),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_835),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_885),
.B(n_888),
.Y(n_1024)
);

BUFx10_ASAP7_75t_L g1025 ( 
.A(n_881),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_829),
.A2(n_721),
.B1(n_775),
.B2(n_664),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_812),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_849),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_875),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_835),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_860),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_860),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_866),
.B(n_867),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_826),
.B(n_891),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_881),
.B(n_876),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_875),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_829),
.B(n_388),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_830),
.B(n_721),
.Y(n_1038)
);

INVx8_ASAP7_75t_L g1039 ( 
.A(n_875),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_870),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_815),
.A2(n_889),
.B(n_887),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_870),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_814),
.A2(n_721),
.B1(n_888),
.B2(n_885),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_888),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_925),
.B(n_1035),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1028),
.B(n_969),
.Y(n_1046)
);

INVx4_ASAP7_75t_SL g1047 ( 
.A(n_992),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_965),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_965),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_936),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_927),
.A2(n_948),
.B1(n_1026),
.B2(n_1043),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_996),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_965),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_925),
.B(n_1035),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_927),
.A2(n_948),
.B1(n_1043),
.B2(n_1014),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_SL g1056 ( 
.A(n_929),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_1019),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_950),
.A2(n_961),
.B1(n_1018),
.B2(n_934),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_963),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_926),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_924),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_967),
.B(n_949),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_945),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1014),
.A2(n_1037),
.B1(n_953),
.B2(n_968),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_925),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_973),
.B(n_947),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_930),
.B(n_934),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1017),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_933),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1031),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1032),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_1002),
.Y(n_1072)
);

CKINVDCx11_ASAP7_75t_R g1073 ( 
.A(n_941),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_930),
.B(n_944),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1016),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_933),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_943),
.A2(n_1015),
.B1(n_1038),
.B2(n_983),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_944),
.B(n_956),
.Y(n_1078)
);

BUFx2_ASAP7_75t_R g1079 ( 
.A(n_982),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1035),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1023),
.Y(n_1081)
);

OAI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_956),
.A2(n_1044),
.B1(n_1024),
.B2(n_1018),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_931),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_971),
.A2(n_976),
.B(n_1001),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1022),
.B(n_1024),
.Y(n_1085)
);

INVxp33_ASAP7_75t_L g1086 ( 
.A(n_935),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_990),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_937),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_942),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1022),
.B(n_1044),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_SL g1091 ( 
.A1(n_943),
.A2(n_1015),
.B1(n_989),
.B2(n_966),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_1003),
.B(n_958),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_997),
.B(n_1001),
.Y(n_1094)
);

OAI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_932),
.A2(n_937),
.B1(n_960),
.B2(n_991),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1011),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_995),
.B(n_952),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1021),
.A2(n_1034),
.B1(n_939),
.B2(n_1012),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_986),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_933),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_960),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1027),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_954),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_962),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_979),
.B(n_1030),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1004),
.Y(n_1107)
);

AO21x2_ASAP7_75t_L g1108 ( 
.A1(n_957),
.A2(n_959),
.B(n_981),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_995),
.B(n_977),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_972),
.A2(n_1004),
.B1(n_994),
.B2(n_1025),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1039),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1019),
.A2(n_1025),
.B1(n_974),
.B2(n_946),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_975),
.B(n_1033),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1005),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_985),
.Y(n_1115)
);

BUFx4f_ASAP7_75t_SL g1116 ( 
.A(n_1000),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_975),
.B(n_964),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_952),
.B(n_977),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_940),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_L g1120 ( 
.A1(n_940),
.A2(n_1020),
.B(n_1041),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_980),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_987),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1009),
.B(n_1007),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1039),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1029),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_964),
.B(n_1033),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1029),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_928),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_978),
.A2(n_970),
.B1(n_951),
.B2(n_938),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1013),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_987),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1039),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_1013),
.A2(n_984),
.B(n_999),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_998),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_951),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_998),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1036),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_999),
.A2(n_1036),
.B(n_1040),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1006),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_993),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1042),
.B(n_1006),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1006),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_988),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1010),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_925),
.B(n_1035),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_963),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_950),
.B(n_885),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_950),
.B(n_885),
.Y(n_1149)
);

INVx8_ASAP7_75t_L g1150 ( 
.A(n_933),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_967),
.B(n_949),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1062),
.B(n_1151),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1045),
.B(n_1146),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1082),
.B(n_1067),
.Y(n_1154)
);

AO21x1_ASAP7_75t_SL g1155 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_1084),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1086),
.B(n_1148),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1062),
.B(n_1151),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1045),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1088),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1081),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1145),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1107),
.B(n_1114),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1120),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1045),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1114),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1107),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1073),
.Y(n_1167)
);

INVxp33_ASAP7_75t_SL g1168 ( 
.A(n_1073),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1146),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1067),
.B(n_1074),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1146),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1119),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1081),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1074),
.B(n_1078),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1149),
.B(n_1058),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1051),
.A2(n_1046),
.B(n_1077),
.Y(n_1176)
);

CKINVDCx9p33_ASAP7_75t_R g1177 ( 
.A(n_1106),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1049),
.B2(n_1065),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1094),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1131),
.A2(n_1134),
.B(n_1094),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1078),
.B(n_1085),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1054),
.B(n_1065),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1131),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1046),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1090),
.B(n_1093),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1108),
.A2(n_1099),
.B(n_1096),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1108),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1093),
.B(n_1071),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1096),
.A2(n_1099),
.B(n_1139),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1054),
.B(n_1080),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1063),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1054),
.B(n_1080),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1054),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1068),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1049),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1091),
.B(n_1066),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1053),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1095),
.B(n_1102),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1047),
.B(n_1072),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1102),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1092),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1059),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1110),
.A2(n_1066),
.B(n_1136),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1124),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1124),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1136),
.A2(n_1135),
.B(n_1137),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1087),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1104),
.B(n_1147),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1147),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1180),
.B(n_1052),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1179),
.B(n_1097),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1195),
.B(n_1047),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1172),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1155),
.A2(n_1098),
.B1(n_1097),
.B2(n_1109),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1180),
.B(n_1109),
.Y(n_1219)
);

OAI33xp33_ASAP7_75t_L g1220 ( 
.A1(n_1210),
.A2(n_1121),
.A3(n_1100),
.B1(n_1105),
.B2(n_1122),
.B3(n_1141),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1188),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1154),
.B(n_1143),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1160),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1173),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1165),
.B(n_1113),
.Y(n_1225)
);

OR2x2_ASAP7_75t_SL g1226 ( 
.A(n_1206),
.B(n_1057),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1155),
.A2(n_1109),
.B1(n_1089),
.B2(n_1117),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1180),
.B(n_1143),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1180),
.B(n_1142),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1162),
.B(n_1142),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1162),
.B(n_1072),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1165),
.B(n_1144),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1175),
.A2(n_1089),
.B1(n_1118),
.B2(n_1112),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_1137),
.B(n_1135),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1166),
.B(n_1144),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1203),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1188),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1207),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1207),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1154),
.B(n_1140),
.Y(n_1240)
);

INVxp67_ASAP7_75t_L g1241 ( 
.A(n_1159),
.Y(n_1241)
);

BUFx2_ASAP7_75t_SL g1242 ( 
.A(n_1203),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1186),
.B(n_1126),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1186),
.B(n_1128),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1161),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1176),
.A2(n_1118),
.B1(n_1127),
.B2(n_1075),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1186),
.B(n_1198),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1186),
.B(n_1138),
.Y(n_1248)
);

NOR2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1195),
.B(n_1129),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1163),
.A2(n_1111),
.B(n_1101),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1187),
.B(n_1115),
.Y(n_1251)
);

INVx4_ASAP7_75t_SL g1252 ( 
.A(n_1202),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1209),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1191),
.A2(n_1111),
.B(n_1101),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1245),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1219),
.B(n_1187),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1226),
.B(n_1189),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1219),
.B(n_1183),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_SL g1259 ( 
.A(n_1249),
.B(n_1201),
.Y(n_1259)
);

OAI221xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1233),
.A2(n_1201),
.B1(n_1199),
.B2(n_1205),
.C(n_1156),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1233),
.A2(n_1199),
.B1(n_1184),
.B2(n_1170),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1227),
.A2(n_1178),
.B1(n_1203),
.B2(n_1183),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1246),
.A2(n_1170),
.B1(n_1181),
.B2(n_1184),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1241),
.B(n_1223),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1214),
.A2(n_1192),
.B1(n_1194),
.B2(n_1183),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1229),
.B(n_1183),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1241),
.B(n_1182),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1229),
.B(n_1183),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1229),
.B(n_1192),
.Y(n_1269)
);

OAI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1218),
.A2(n_1234),
.B1(n_1240),
.B2(n_1222),
.C(n_1211),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1234),
.B(n_1208),
.C(n_1204),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1214),
.A2(n_1240),
.B1(n_1222),
.B2(n_1211),
.C(n_1247),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1251),
.B(n_1192),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1224),
.B(n_1208),
.C(n_1204),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1251),
.B(n_1192),
.Y(n_1275)
);

NAND4xp25_ASAP7_75t_L g1276 ( 
.A(n_1214),
.B(n_1210),
.C(n_1168),
.D(n_1185),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1251),
.B(n_1194),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1230),
.B(n_1174),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1230),
.B(n_1174),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1228),
.B(n_1194),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1243),
.B(n_1185),
.C(n_1200),
.Y(n_1282)
);

AND2x2_ASAP7_75t_SL g1283 ( 
.A(n_1226),
.B(n_1194),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1225),
.B(n_1190),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1242),
.A2(n_1167),
.B1(n_1083),
.B2(n_1177),
.Y(n_1285)
);

OAI221xp5_ASAP7_75t_L g1286 ( 
.A1(n_1243),
.A2(n_1171),
.B1(n_1158),
.B2(n_1169),
.C(n_1164),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1225),
.B(n_1190),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1228),
.B(n_1198),
.Y(n_1288)
);

NAND2x1_ASAP7_75t_L g1289 ( 
.A(n_1250),
.B(n_1153),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1215),
.B(n_1231),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1215),
.B(n_1152),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1244),
.B(n_1200),
.C(n_1196),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1215),
.B(n_1152),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1228),
.B(n_1157),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1216),
.B(n_1153),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1231),
.B(n_1157),
.Y(n_1296)
);

OAI221xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1247),
.A2(n_1164),
.B1(n_1158),
.B2(n_1169),
.C(n_1171),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1231),
.B(n_1158),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1232),
.B(n_1164),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1244),
.B(n_1206),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1235),
.B(n_1171),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1244),
.A2(n_1193),
.B(n_1197),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1300),
.B(n_1248),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1257),
.B(n_1248),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1255),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1255),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1257),
.B(n_1248),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1300),
.B(n_1250),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1289),
.B(n_1250),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1294),
.B(n_1250),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1288),
.Y(n_1311)
);

AND2x2_ASAP7_75t_SL g1312 ( 
.A(n_1283),
.B(n_1153),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1283),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1294),
.B(n_1250),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1288),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1256),
.B(n_1213),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1256),
.B(n_1213),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1283),
.B(n_1213),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1280),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1264),
.B(n_1238),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1284),
.B(n_1238),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1280),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1258),
.B(n_1252),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1269),
.B(n_1213),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1302),
.B(n_1292),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1289),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1287),
.B(n_1239),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1266),
.B(n_1253),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1266),
.B(n_1221),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1268),
.B(n_1221),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1282),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1302),
.B(n_1217),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1299),
.B(n_1239),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1258),
.B(n_1252),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1273),
.B(n_1237),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1292),
.Y(n_1336)
);

BUFx2_ASAP7_75t_SL g1337 ( 
.A(n_1295),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1281),
.B(n_1217),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1273),
.B(n_1252),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1309),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1305),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1331),
.B(n_1278),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1305),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1340),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1325),
.A2(n_1260),
.B(n_1261),
.Y(n_1346)
);

NOR2x1_ASAP7_75t_R g1347 ( 
.A(n_1337),
.B(n_1050),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1313),
.B(n_1275),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1313),
.B(n_1275),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1306),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1309),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1306),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1323),
.B(n_1252),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1326),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1309),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1311),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1311),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1304),
.B(n_1290),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1304),
.B(n_1267),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1325),
.A2(n_1276),
.B1(n_1261),
.B2(n_1270),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1331),
.B(n_1340),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1312),
.B(n_1279),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1337),
.B(n_1316),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1316),
.B(n_1296),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1315),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1323),
.B(n_1334),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1320),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1336),
.B(n_1291),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_R g1371 ( 
.A(n_1339),
.B(n_1050),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1307),
.B(n_1301),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1307),
.B(n_1293),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1336),
.B(n_1272),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1316),
.B(n_1298),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1315),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1317),
.B(n_1339),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1317),
.B(n_1265),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1354),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1342),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1346),
.B(n_1338),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1342),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1354),
.B(n_1323),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1347),
.B(n_1285),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1346),
.B(n_1338),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1344),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1362),
.A2(n_1363),
.B(n_1347),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1344),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1374),
.A2(n_1259),
.B(n_1345),
.C(n_1276),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1350),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1350),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1368),
.B(n_1334),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1370),
.B(n_1320),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1352),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1370),
.B(n_1321),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1353),
.B(n_1339),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1374),
.A2(n_1285),
.B1(n_1297),
.B2(n_1271),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1353),
.B(n_1339),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1352),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1343),
.B(n_1335),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1371),
.B(n_1079),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1354),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1357),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1354),
.B(n_1334),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1363),
.B(n_1334),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1357),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1368),
.B(n_1318),
.Y(n_1408)
);

NAND2x1_ASAP7_75t_L g1409 ( 
.A(n_1368),
.B(n_1318),
.Y(n_1409)
);

AOI21xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1345),
.A2(n_1262),
.B(n_1318),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1361),
.B(n_1324),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1358),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1358),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1367),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1367),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1343),
.B(n_1335),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1378),
.A2(n_1263),
.B1(n_1220),
.B2(n_1271),
.Y(n_1417)
);

OAI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1369),
.A2(n_1332),
.B(n_1286),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1364),
.B(n_1328),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1360),
.B(n_1321),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1381),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1382),
.B(n_1364),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1381),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1404),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1383),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1394),
.B(n_1360),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1384),
.B(n_1377),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1384),
.B(n_1377),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1387),
.Y(n_1431)
);

AOI222xp33_ASAP7_75t_L g1432 ( 
.A1(n_1386),
.A2(n_1263),
.B1(n_1371),
.B2(n_1332),
.C1(n_1378),
.C2(n_1365),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1385),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1389),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1409),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1379),
.B(n_1365),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1417),
.B(n_1366),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1396),
.B(n_1373),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1388),
.B(n_1361),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1242),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1421),
.B(n_1373),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1420),
.B(n_1359),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1379),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1391),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1405),
.B(n_1348),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1379),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1392),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1395),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1393),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1407),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1393),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1393),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1412),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1418),
.B(n_1366),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1380),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1390),
.A2(n_1274),
.B(n_1236),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1410),
.B(n_1348),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1433),
.B(n_1398),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1440),
.A2(n_1439),
.B1(n_1456),
.B2(n_1457),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1439),
.A2(n_1406),
.B1(n_1403),
.B2(n_1380),
.C(n_1415),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1432),
.B(n_1402),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_SL g1462 ( 
.A(n_1437),
.B(n_1406),
.C(n_1419),
.Y(n_1462)
);

AOI31xp33_ASAP7_75t_L g1463 ( 
.A1(n_1457),
.A2(n_1403),
.A3(n_1405),
.B(n_1408),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1424),
.B(n_1408),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1454),
.B(n_1411),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1422),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_SL g1469 ( 
.A(n_1423),
.B(n_1083),
.C(n_1401),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1425),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1440),
.A2(n_1452),
.B1(n_1446),
.B2(n_1451),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1431),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1435),
.A2(n_1408),
.B(n_1351),
.C(n_1308),
.Y(n_1474)
);

AOI21xp33_ASAP7_75t_L g1475 ( 
.A1(n_1440),
.A2(n_1400),
.B(n_1413),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1440),
.A2(n_1359),
.B1(n_1351),
.B2(n_1372),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1446),
.A2(n_1414),
.B(n_1400),
.Y(n_1477)
);

AOI31xp33_ASAP7_75t_L g1478 ( 
.A1(n_1451),
.A2(n_1056),
.A3(n_1220),
.B(n_1349),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1428),
.B(n_1372),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1441),
.B(n_1333),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1349),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1436),
.A2(n_1351),
.B1(n_1249),
.B2(n_1216),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1464),
.B(n_1424),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1445),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1467),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1458),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1465),
.B(n_1429),
.Y(n_1487)
);

NOR3xp33_ASAP7_75t_L g1488 ( 
.A(n_1461),
.B(n_1455),
.C(n_1435),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1468),
.B(n_1443),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1472),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1460),
.B(n_1471),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1473),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1471),
.B(n_1429),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1470),
.B(n_1430),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1479),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1459),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1480),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1481),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1477),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1463),
.Y(n_1501)
);

AOI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1469),
.A2(n_1450),
.B1(n_1434),
.B2(n_1447),
.C1(n_1453),
.C2(n_1444),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1491),
.A2(n_1469),
.B1(n_1436),
.B2(n_1443),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1500),
.A2(n_1478),
.B(n_1475),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1488),
.B(n_1474),
.C(n_1482),
.Y(n_1505)
);

AOI21xp33_ASAP7_75t_L g1506 ( 
.A1(n_1501),
.A2(n_1455),
.B(n_1476),
.Y(n_1506)
);

AOI322xp5_ASAP7_75t_L g1507 ( 
.A1(n_1497),
.A2(n_1436),
.A3(n_1430),
.B1(n_1435),
.B2(n_1443),
.C1(n_1448),
.C2(n_1351),
.Y(n_1507)
);

AOI211xp5_ASAP7_75t_L g1508 ( 
.A1(n_1488),
.A2(n_1442),
.B(n_1341),
.C(n_1356),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1486),
.B(n_1502),
.C(n_1489),
.Y(n_1509)
);

NOR3xp33_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1485),
.C(n_1494),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1483),
.Y(n_1511)
);

AOI31xp33_ASAP7_75t_L g1512 ( 
.A1(n_1484),
.A2(n_1116),
.A3(n_1309),
.B(n_1355),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1496),
.Y(n_1513)
);

XNOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1509),
.B(n_1499),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1510),
.B(n_1493),
.C(n_1498),
.Y(n_1516)
);

NOR3x1_ASAP7_75t_L g1517 ( 
.A(n_1504),
.B(n_1495),
.C(n_1492),
.Y(n_1517)
);

NOR3xp33_ASAP7_75t_L g1518 ( 
.A(n_1506),
.B(n_1490),
.C(n_1487),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_L g1519 ( 
.A(n_1513),
.B(n_1060),
.Y(n_1519)
);

NOR4xp25_ASAP7_75t_L g1520 ( 
.A(n_1505),
.B(n_1341),
.C(n_1356),
.D(n_1355),
.Y(n_1520)
);

NOR2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1507),
.B(n_1060),
.Y(n_1521)
);

OAI322xp33_ASAP7_75t_L g1522 ( 
.A1(n_1503),
.A2(n_1341),
.A3(n_1356),
.B1(n_1355),
.B2(n_1376),
.C1(n_1326),
.C2(n_1327),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1520),
.A2(n_1508),
.B1(n_1512),
.B2(n_1376),
.C(n_1326),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1516),
.B(n_1075),
.Y(n_1524)
);

NOR2x1p5_ASAP7_75t_SL g1525 ( 
.A(n_1514),
.B(n_1327),
.Y(n_1525)
);

OAI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1518),
.A2(n_1103),
.B1(n_1236),
.B2(n_1212),
.C(n_1333),
.Y(n_1526)
);

NAND4xp75_ASAP7_75t_L g1527 ( 
.A(n_1517),
.B(n_1076),
.C(n_1308),
.D(n_1317),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1524),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1525),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1527),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1526),
.A2(n_1521),
.B1(n_1515),
.B2(n_1519),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1523),
.B(n_1375),
.Y(n_1532)
);

NOR2x2_ASAP7_75t_L g1533 ( 
.A(n_1527),
.B(n_1522),
.Y(n_1533)
);

OAI211xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1531),
.A2(n_1103),
.B(n_1319),
.C(n_1322),
.Y(n_1534)
);

NOR3xp33_ASAP7_75t_L g1535 ( 
.A(n_1529),
.B(n_1069),
.C(n_1076),
.Y(n_1535)
);

NAND4xp75_ASAP7_75t_L g1536 ( 
.A(n_1528),
.B(n_1308),
.C(n_1314),
.D(n_1310),
.Y(n_1536)
);

NAND3x1_ASAP7_75t_SL g1537 ( 
.A(n_1533),
.B(n_1123),
.C(n_1310),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1532),
.B(n_1319),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1538),
.Y(n_1539)
);

NAND4xp25_ASAP7_75t_SL g1540 ( 
.A(n_1535),
.B(n_1530),
.C(n_1274),
.D(n_1310),
.Y(n_1540)
);

XNOR2xp5_ASAP7_75t_L g1541 ( 
.A(n_1537),
.B(n_1125),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1539),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1542),
.Y(n_1543)
);

AOI221x1_ASAP7_75t_L g1544 ( 
.A1(n_1543),
.A2(n_1534),
.B1(n_1541),
.B2(n_1540),
.C(n_1536),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1543),
.A2(n_1375),
.B(n_1069),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1544),
.A2(n_1254),
.B(n_1314),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1545),
.B(n_1322),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1546),
.A2(n_1123),
.B1(n_1057),
.B2(n_1303),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1547),
.A2(n_1069),
.B(n_1125),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1549),
.A2(n_1548),
.B(n_1150),
.Y(n_1550)
);

AOI322xp5_ASAP7_75t_L g1551 ( 
.A1(n_1550),
.A2(n_1314),
.A3(n_1303),
.B1(n_1324),
.B2(n_1328),
.C1(n_1329),
.C2(n_1330),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1551),
.A2(n_1057),
.B1(n_1133),
.B2(n_1132),
.C(n_1212),
.Y(n_1552)
);

AOI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1552),
.A2(n_1133),
.B(n_1212),
.C(n_1236),
.Y(n_1553)
);


endmodule