module real_jpeg_11949_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_275, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_275;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_244;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_2),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_35),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_3),
.A2(n_35),
.B1(n_146),
.B2(n_158),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_7),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_41),
.B1(n_44),
.B2(n_150),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_7),
.A2(n_98),
.B1(n_99),
.B2(n_150),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_9),
.A2(n_43),
.B1(n_98),
.B2(n_99),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_9),
.A2(n_43),
.B1(n_146),
.B2(n_158),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_27),
.C(n_46),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_28),
.B1(n_41),
.B2(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_10),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_10),
.B(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_28),
.B1(n_98),
.B2(n_99),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_55),
.B(n_99),
.C(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_28),
.B1(n_146),
.B2(n_158),
.Y(n_163)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_254),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_235),
.B(n_253),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_214),
.B(n_234),
.Y(n_14)
);

AOI321xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_174),
.A3(n_207),
.B1(n_212),
.B2(n_213),
.C(n_275),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_137),
.B(n_173),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_114),
.B(n_136),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_91),
.B(n_113),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_69),
.B(n_90),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_36),
.B1(n_37),
.B2(n_59),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_23),
.B(n_87),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_33),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_109)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_27),
.B(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_28),
.A2(n_44),
.B(n_56),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_28),
.B(n_99),
.C(n_127),
.Y(n_145)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_30),
.A2(n_87),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_32),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_80),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_33),
.A2(n_149),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_39),
.B(n_66),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_39),
.A2(n_171),
.B(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_40),
.B(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_45),
.B(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_45),
.Y(n_172)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_57),
.C(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_53),
.B(n_104),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_53),
.A2(n_101),
.B(n_104),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_53),
.A2(n_167),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_54),
.B(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_56),
.B1(n_98),
.B2(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_68),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_83),
.B(n_89),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_77),
.B(n_82),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_81),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_93),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_105),
.C(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_99),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_100),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_102),
.B(n_131),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_102),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_106),
.A2(n_172),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_106),
.B(n_118),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_108),
.A2(n_109),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_108),
.A2(n_109),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_109),
.B(n_231),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_109),
.A2(n_242),
.B(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_135),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_135),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_122),
.B1(n_123),
.B2(n_134),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.C(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_142),
.C(n_152),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.CI(n_129),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_126),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_126),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_128),
.B1(n_146),
.B2(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_130),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_130),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_139),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_152),
.B2(n_153),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_148),
.B2(n_151),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_166),
.C(n_169),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_161),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_160),
.A2(n_163),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_179),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_169),
.A2(n_170),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_201),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_201),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_186),
.C(n_197),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_184),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_178),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_194),
.C(n_195),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_206),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_203),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_211),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_216),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_233),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_229),
.B2(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_230),
.C(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_222),
.C(n_227),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.C(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B(n_252),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_252),
.A2(n_261),
.B1(n_262),
.B2(n_272),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_273),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);


endmodule