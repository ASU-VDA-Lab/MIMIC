module fake_jpeg_32046_n_360 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_14),
.B(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_49),
.B(n_82),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_26),
.A2(n_16),
.B1(n_35),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_56),
.A2(n_40),
.B1(n_15),
.B2(n_7),
.Y(n_143)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_59),
.B(n_60),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_8),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_64),
.B(n_66),
.Y(n_113)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_67),
.B(n_73),
.Y(n_128)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_10),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_26),
.B(n_0),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_10),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_12),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_90),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_29),
.B(n_0),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_92),
.Y(n_149)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_21),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_94),
.Y(n_150)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_33),
.B1(n_44),
.B2(n_35),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_13),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_47),
.B(n_43),
.C(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_104),
.B(n_65),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_117),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_43),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_35),
.B1(n_33),
.B2(n_44),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_137),
.B1(n_84),
.B2(n_95),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_44),
.B1(n_30),
.B2(n_42),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_138),
.B1(n_83),
.B2(n_94),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_50),
.Y(n_127)
);

OR2x4_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_24),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_72),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_140),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_24),
.B1(n_37),
.B2(n_23),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_76),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_51),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_32),
.B1(n_40),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_143),
.B1(n_74),
.B2(n_63),
.Y(n_160)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_111),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_153),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_59),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_48),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_175),
.B1(n_102),
.B2(n_101),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_164),
.A2(n_174),
.B1(n_186),
.B2(n_109),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_167),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_48),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_105),
.B(n_3),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_52),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_53),
.B1(n_98),
.B2(n_52),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_145),
.A3(n_121),
.B1(n_125),
.B2(n_99),
.Y(n_209)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_98),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_3),
.B1(n_5),
.B2(n_136),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_100),
.A2(n_3),
.B1(n_5),
.B2(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_177),
.A2(n_131),
.B1(n_100),
.B2(n_102),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_150),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_133),
.B1(n_124),
.B2(n_145),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_107),
.B(n_106),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_144),
.B(n_108),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_104),
.B(n_137),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_124),
.B(n_103),
.C(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_175),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_203),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_144),
.B1(n_108),
.B2(n_145),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_142),
.B1(n_130),
.B2(n_146),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_147),
.B1(n_146),
.B2(n_109),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_184),
.B(n_166),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_112),
.A3(n_123),
.B1(n_121),
.B2(n_114),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_165),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_216),
.B1(n_171),
.B2(n_161),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_153),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_218),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_153),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_223),
.B1(n_203),
.B2(n_176),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_159),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_157),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_167),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_169),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_173),
.C(n_154),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_206),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_154),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_236),
.B(n_189),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_238),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_211),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_216),
.B1(n_202),
.B2(n_206),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_245),
.B1(n_254),
.B2(n_255),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_246),
.C(n_207),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_197),
.B1(n_209),
.B2(n_213),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_213),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_221),
.B(n_233),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_251),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_205),
.B1(n_201),
.B2(n_164),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_234),
.A2(n_205),
.B1(n_208),
.B2(n_171),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_217),
.B1(n_211),
.B2(n_207),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_236),
.B(n_220),
.C(n_228),
.D(n_230),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_263),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_223),
.B1(n_226),
.B2(n_232),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_267),
.B1(n_271),
.B2(n_260),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_229),
.B(n_237),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_241),
.B(n_251),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_229),
.B1(n_231),
.B2(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.C(n_258),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_178),
.C(n_172),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_277),
.A2(n_245),
.B1(n_240),
.B2(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_284),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_275),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_244),
.C(n_246),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_282),
.C(n_286),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_257),
.B(n_252),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_289),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_247),
.B1(n_249),
.B2(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_267),
.B1(n_262),
.B2(n_272),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_252),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_242),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_241),
.B1(n_196),
.B2(n_238),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_266),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_204),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_302),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_297),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_263),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_295),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_309),
.B1(n_279),
.B2(n_280),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_294),
.C(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_238),
.C(n_204),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_280),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_312),
.B(n_316),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_320),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_293),
.B1(n_291),
.B2(n_288),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_293),
.B1(n_285),
.B2(n_261),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_300),
.A3(n_304),
.B1(n_303),
.B2(n_287),
.C1(n_295),
.C2(n_270),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_298),
.B(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_325),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_296),
.C(n_306),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_287),
.B(n_268),
.C(n_273),
.D(n_191),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_328),
.B(n_329),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_278),
.B(n_224),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_310),
.C(n_320),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_337),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_315),
.C(n_321),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_335),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_322),
.C(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_314),
.C(n_199),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_191),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_339),
.B(n_198),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_199),
.C(n_158),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_162),
.B(n_198),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_336),
.A2(n_328),
.B(n_171),
.C(n_214),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_342),
.A2(n_112),
.B1(n_151),
.B2(n_156),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_344),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_338),
.A2(n_168),
.B(n_186),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_345),
.A2(n_99),
.B(n_125),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_347),
.A2(n_183),
.B1(n_179),
.B2(n_152),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_341),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_349),
.B(n_352),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_350),
.A2(n_342),
.B(n_156),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_352),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_353),
.A2(n_349),
.B(n_351),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_357),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_354),
.C(n_148),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_181),
.B(n_329),
.Y(n_360)
);


endmodule