module real_jpeg_31272_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_17),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_1),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_63),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

INVx3_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_3),
.A2(n_57),
.B1(n_70),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_3),
.A2(n_70),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_3),
.B(n_112),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_3),
.B(n_100),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_3),
.B(n_390),
.C(n_393),
.Y(n_389)
);

NAND2xp67_ASAP7_75t_L g405 ( 
.A(n_3),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_3),
.B(n_27),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_6),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_6),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_105),
.B1(n_149),
.B2(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_7),
.A2(n_105),
.B1(n_231),
.B2(n_235),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_9),
.Y(n_303)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

OAI211xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_207),
.B(n_446),
.C(n_448),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_18),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_15),
.B(n_447),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_16),
.B(n_18),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_206),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_186),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_20),
.B(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_145),
.C(n_158),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_22),
.A2(n_145),
.B1(n_146),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_22),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_109),
.B2(n_144),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_67),
.B2(n_68),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_26),
.B(n_191),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_43),
.B(n_61),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_43),
.B1(n_61),
.B2(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_27),
.B(n_148),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_27),
.A2(n_148),
.B(n_162),
.Y(n_244)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_29),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_29)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_30),
.Y(n_236)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_32),
.Y(n_182)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_32),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_32),
.Y(n_234)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_36),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_38),
.Y(n_184)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_L g162 ( 
.A(n_44),
.B(n_163),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_45),
.A2(n_164),
.B(n_221),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B1(n_54),
.B2(n_57),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_53),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_53),
.Y(n_350)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_60),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_63),
.A2(n_178),
.B(n_183),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_68),
.B(n_185),
.C(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_81),
.B1(n_100),
.B2(n_101),
.Y(n_68)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_69),
.A2(n_81),
.B(n_82),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_76),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_74),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_75),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_76),
.Y(n_365)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_92),
.B1(n_95),
.B2(n_99),
.Y(n_91)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

NOR2x1p5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_85),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_85),
.Y(n_359)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

NOR2x1p5_ASAP7_75t_L g247 ( 
.A(n_110),
.B(n_248),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g272 ( 
.A1(n_110),
.A2(n_245),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_110),
.B(n_220),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

AO22x2_ASAP7_75t_L g216 ( 
.A1(n_111),
.A2(n_157),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_111),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_123),
.B(n_136),
.Y(n_111)
);

OAI22x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_115),
.Y(n_292)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2x1_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_134),
.Y(n_299)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_140),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_159),
.B1(n_168),
.B2(n_185),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_189),
.B1(n_190),
.B2(n_203),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_145),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_156),
.B(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_157),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_157),
.B(n_218),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_157),
.B(n_220),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_158),
.B(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2x1_ASAP7_75t_SL g271 ( 
.A(n_160),
.B(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_168),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

NAND2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OR2x6_ASAP7_75t_L g285 ( 
.A(n_170),
.B(n_252),
.Y(n_285)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_175),
.Y(n_406)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_185),
.B(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_201),
.B2(n_202),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_197),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_207),
.B(n_449),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_436),
.B(n_443),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_423),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_336),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_310),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_275),
.Y(n_211)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_212),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_264),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_213),
.B(n_264),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_242),
.C(n_246),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_240),
.B2(n_241),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_216),
.B(n_250),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_216),
.A2(n_240),
.B1(n_283),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_219),
.A2(n_247),
.B(n_261),
.Y(n_270)
);

NAND2x1p5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_251),
.Y(n_250)
);

XOR2x2_ASAP7_75t_SL g281 ( 
.A(n_220),
.B(n_222),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_220),
.A2(n_251),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_220),
.Y(n_316)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_220),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_220),
.A2(n_284),
.B1(n_285),
.B2(n_316),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_220),
.A2(n_316),
.B1(n_384),
.B2(n_385),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_230),
.B1(n_237),
.B2(n_239),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_230),
.B1(n_252),
.B2(n_257),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_249),
.B(n_261),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_263),
.B(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AND3x1_ASAP7_75t_L g319 ( 
.A(n_263),
.B(n_320),
.C(n_321),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_266),
.B(n_271),
.C(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_267),
.B(n_284),
.C(n_334),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_267),
.A2(n_340),
.B(n_342),
.C(n_366),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_267),
.B(n_374),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_270),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_275),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_276),
.B(n_278),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_282),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_281),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_287),
.Y(n_331)
);

NAND2x1p5_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_343),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_284),
.A2(n_285),
.B1(n_334),
.B2(n_335),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_284),
.B(n_371),
.C(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_284),
.B(n_413),
.Y(n_412)
);

CKINVDCx11_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_285),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_285),
.B(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_285),
.B(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_295),
.B(n_300),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx4f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_304),
.B(n_309),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_324),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_311),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_322),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_312),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_318),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_318),
.B1(n_319),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_325),
.B(n_328),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.C(n_332),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_329),
.B(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_342),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_331),
.B(n_333),
.Y(n_421)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI21x1_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_418),
.B(n_422),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_376),
.B(n_417),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_367),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_339),
.B(n_367),
.Y(n_417)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_370),
.C(n_372),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_347),
.B(n_355),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_360),
.B(n_364),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_372),
.B1(n_373),
.B2(n_375),
.Y(n_367)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI21x1_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_381),
.B(n_416),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_401),
.B(n_414),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_397),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_412),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_410),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_420),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_427),
.B(n_433),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_441),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);


endmodule