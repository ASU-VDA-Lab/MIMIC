module fake_jpeg_21984_n_160 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_1),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_32),
.B(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_16),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_39),
.B(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_18),
.B1(n_16),
.B2(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_41),
.B1(n_27),
.B2(n_29),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_44),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_18),
.B1(n_14),
.B2(n_24),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_49),
.B1(n_58),
.B2(n_31),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_53),
.Y(n_66)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_30),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_41),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_25),
.B(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_59),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_44),
.B1(n_43),
.B2(n_26),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_69),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_33),
.B1(n_28),
.B2(n_34),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_75),
.B1(n_58),
.B2(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_30),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_30),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_76),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_44),
.C(n_43),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_56),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_49),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_83),
.B(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_60),
.B1(n_56),
.B2(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_52),
.B(n_55),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_71),
.B(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_48),
.B1(n_45),
.B2(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_95),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_51),
.B(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_45),
.B1(n_26),
.B2(n_24),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_49),
.B1(n_22),
.B2(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_83),
.B(n_72),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_106),
.B(n_87),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_96),
.C(n_66),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_108),
.C(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_67),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_69),
.C(n_70),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_94),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_123),
.C(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_119),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_107),
.A3(n_110),
.B1(n_12),
.B2(n_17),
.C(n_23),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_120),
.Y(n_129)
);

AO221x1_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_74),
.B1(n_78),
.B2(n_90),
.C(n_57),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_121),
.B(n_110),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_81),
.B1(n_88),
.B2(n_91),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_97),
.B(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_97),
.B1(n_65),
.B2(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_65),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_97),
.C(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_103),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_128),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_132),
.C(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_116),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_108),
.C(n_104),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_134),
.B(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_119),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_137),
.B(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_141),
.C(n_114),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_119),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_142),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_122),
.C(n_125),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_145),
.B(n_146),
.Y(n_153)
);

OAI31xp33_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_122),
.A3(n_119),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_92),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_149),
.A3(n_49),
.B1(n_15),
.B2(n_19),
.C1(n_17),
.C2(n_23),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_115),
.B(n_120),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_19),
.A3(n_12),
.B1(n_15),
.B2(n_22),
.C1(n_6),
.C2(n_7),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_6),
.A3(n_10),
.B1(n_9),
.B2(n_4),
.C1(n_11),
.C2(n_7),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_6),
.A3(n_10),
.B1(n_9),
.B2(n_4),
.C1(n_11),
.C2(n_7),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_10),
.C(n_2),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_157),
.B(n_1),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_158)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_159),
.B1(n_3),
.B2(n_77),
.C(n_142),
.Y(n_160)
);


endmodule