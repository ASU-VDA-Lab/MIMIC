module fake_jpeg_8327_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_24),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_31),
.B1(n_20),
.B2(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_48),
.B1(n_24),
.B2(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_26),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_20),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_57),
.C(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_20),
.B1(n_31),
.B2(n_18),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_39),
.B1(n_22),
.B2(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_54),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_61),
.Y(n_109)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_34),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_85),
.B(n_38),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_77),
.B1(n_78),
.B2(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_17),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_40),
.B1(n_22),
.B2(n_25),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_43),
.B1(n_34),
.B2(n_38),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_40),
.B1(n_25),
.B2(n_39),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_32),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_45),
.B(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_27),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_116),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_27),
.B1(n_16),
.B2(n_28),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_54),
.B1(n_59),
.B2(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_103),
.B1(n_70),
.B2(n_61),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_29),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_115),
.B1(n_102),
.B2(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_53),
.B1(n_29),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_27),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_120),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_121),
.B1(n_126),
.B2(n_128),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_82),
.B1(n_69),
.B2(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_111),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_127),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_85),
.B1(n_73),
.B2(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_87),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_85),
.B1(n_88),
.B2(n_68),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_130),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_60),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_64),
.B1(n_21),
.B2(n_30),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_19),
.B(n_17),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_163)
);

AO21x2_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_62),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_64),
.B1(n_21),
.B2(n_32),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_107),
.B(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_11),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_28),
.B(n_17),
.C(n_83),
.D(n_80),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_112),
.B1(n_106),
.B2(n_28),
.C(n_17),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_158),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_100),
.B(n_93),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_150),
.B(n_153),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_175),
.B(n_126),
.C(n_118),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_93),
.B(n_116),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_162),
.C(n_165),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_16),
.B(n_19),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_104),
.B1(n_98),
.B2(n_92),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_171),
.B1(n_139),
.B2(n_120),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_19),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_123),
.C(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_67),
.C(n_98),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_172),
.C(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_169),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_98),
.B1(n_16),
.B2(n_19),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_19),
.C(n_1),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_19),
.B(n_1),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_0),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_198),
.B1(n_199),
.B2(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_193),
.B1(n_197),
.B2(n_187),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_192),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_172),
.B(n_160),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_143),
.C(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_165),
.C(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_152),
.A2(n_126),
.B1(n_117),
.B2(n_145),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_126),
.B1(n_133),
.B2(n_137),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_207),
.C(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_166),
.B1(n_175),
.B2(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_150),
.B1(n_146),
.B2(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_180),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_156),
.B(n_173),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_209),
.B(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_162),
.C(n_158),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_146),
.B1(n_160),
.B2(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_177),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_137),
.C(n_1),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_0),
.C(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_191),
.C(n_188),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_9),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_177),
.B(n_180),
.C(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_227),
.B1(n_230),
.B2(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_228),
.C(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_183),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_194),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_186),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_209),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_221),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_202),
.B1(n_217),
.B2(n_205),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_241),
.B1(n_243),
.B2(n_194),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_223),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_201),
.B1(n_206),
.B2(n_211),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_214),
.B1(n_194),
.B2(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_238),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_223),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_255),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_234),
.CI(n_232),
.CON(n_251),
.SN(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_254),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_236),
.B(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_8),
.C(n_13),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_243),
.B(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_12),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_8),
.B(n_13),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_11),
.B(n_15),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_270),
.B1(n_259),
.B2(n_266),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_269),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_258),
.B(n_257),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_251),
.A3(n_10),
.B1(n_5),
.B2(n_7),
.C1(n_12),
.C2(n_13),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_275),
.A3(n_5),
.B1(n_10),
.B2(n_12),
.C1(n_15),
.C2(n_3),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_251),
.A3(n_256),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_4),
.B(n_274),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_4),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_4),
.Y(n_281)
);


endmodule