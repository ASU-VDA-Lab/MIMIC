module fake_aes_9073_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx3_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_1), .B(n_2), .Y(n_4) );
O2A1O1Ixp33_ASAP7_75t_SL g5 ( .A1(n_4), .A2(n_3), .B(n_1), .C(n_0), .Y(n_5) );
OAI22xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B1(n_2), .B2(n_4), .Y(n_6) );
INVxp67_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx4_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_11), .Y(n_12) );
endmodule