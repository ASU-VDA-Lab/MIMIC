module fake_netlist_5_661_n_1003 (n_137, n_294, n_82, n_194, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_286, n_122, n_282, n_10, n_24, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_9, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1003);

input n_137;
input n_294;
input n_82;
input n_194;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_9;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1003;

wire n_924;
wire n_676;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_525;
wire n_397;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_823;
wire n_983;
wire n_725;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_526;
wire n_915;
wire n_719;
wire n_443;
wire n_372;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_498;
wire n_516;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_812;
wire n_842;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_883;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_519;
wire n_406;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_918;
wire n_942;
wire n_381;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_428;
wire n_379;
wire n_833;
wire n_514;
wire n_457;
wire n_570;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_839;
wire n_901;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_369;
wire n_675;
wire n_888;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_517;
wire n_342;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_388;
wire n_761;
wire n_903;
wire n_740;
wire n_329;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_907;
wire n_722;
wire n_458;
wire n_770;
wire n_844;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_585;
wire n_349;
wire n_616;
wire n_953;
wire n_601;
wire n_917;
wire n_966;
wire n_987;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_868;
wire n_803;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_533;
wire n_950;
wire n_747;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_39),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_292),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_301),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_305),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_79),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_138),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_295),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_16),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_240),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_107),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_86),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_156),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_126),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_153),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_239),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_261),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_8),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_34),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_139),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_217),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_277),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_182),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_185),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_142),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_161),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_66),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_242),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_28),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_150),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_237),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_293),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_153),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_13),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_231),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_83),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_243),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_244),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_144),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_249),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_129),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_256),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_145),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_230),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_41),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_53),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_228),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_213),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_120),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_139),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_297),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_45),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_104),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_290),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_51),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_219),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_14),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_38),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_48),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_127),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_302),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_59),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_275),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_57),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_235),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_128),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_304),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_257),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_236),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_49),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_160),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_168),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_285),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_303),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_162),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_300),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_43),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_177),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_124),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_103),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_312),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_131),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_227),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_233),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_116),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_74),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_269),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_110),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_215),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_263),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_82),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_280),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_322),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_317),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_318),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_376),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_316),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_422),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_319),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_424),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_324),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_323),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_326),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_336),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_328),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_332),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_330),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_337),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_338),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_397),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_340),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_341),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_321),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_366),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_339),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_327),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_363),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_327),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_387),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_343),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_346),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_411),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_349),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_352),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_468),
.A2(n_380),
.B1(n_379),
.B2(n_364),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_431),
.B(n_396),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_453),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_432),
.B(n_347),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_448),
.B(n_367),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_437),
.B(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_460),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_439),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_437),
.A2(n_342),
.B1(n_353),
.B2(n_345),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_461),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_450),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_462),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_451),
.B(n_425),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_446),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_442),
.A2(n_384),
.B(n_357),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_386),
.B(n_354),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_423),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_465),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_467),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_474),
.B(n_392),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_327),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_426),
.B(n_378),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_475),
.B(n_408),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_471),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_476),
.B(n_410),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_473),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_478),
.A2(n_356),
.B1(n_359),
.B2(n_355),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_413),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_403),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_481),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_482),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_483),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_477),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_487),
.B(n_455),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_539),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_486),
.A2(n_469),
.B1(n_479),
.B2(n_457),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_527),
.B(n_485),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_497),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_535),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_507),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_512),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_514),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_535),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

CKINVDCx8_ASAP7_75t_R g555 ( 
.A(n_513),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_529),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_537),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_499),
.B(n_447),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_536),
.Y(n_560)
);

BUFx6f_ASAP7_75t_SL g561 ( 
.A(n_505),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_538),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_494),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_459),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_488),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_489),
.A2(n_374),
.B1(n_382),
.B2(n_372),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_503),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_491),
.B(n_358),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_447),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_500),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_490),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_525),
.B(n_463),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_498),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_501),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_530),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_533),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_525),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_593),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_575),
.B(n_519),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_559),
.B(n_516),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_L g597 ( 
.A(n_542),
.B(n_528),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_562),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_562),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_524),
.C(n_532),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_526),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_510),
.C(n_504),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_570),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_582),
.B(n_526),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_534),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_534),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_571),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_522),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_573),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_463),
.C(n_385),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_578),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_553),
.B(n_417),
.Y(n_614)
);

OAI21xp33_ASAP7_75t_L g615 ( 
.A1(n_566),
.A2(n_395),
.B(n_383),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_574),
.B(n_362),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_540),
.B(n_371),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_567),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_543),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_546),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_547),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_549),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_415),
.C(n_409),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_550),
.B(n_373),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_561),
.A2(n_377),
.B1(n_381),
.B2(n_375),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_388),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_552),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_554),
.B(n_394),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_556),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_563),
.B(n_398),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_557),
.Y(n_633)
);

INVx8_ASAP7_75t_L g634 ( 
.A(n_561),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_563),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_563),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_558),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_583),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_418),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_577),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_583),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_572),
.B(n_399),
.Y(n_642)
);

NOR3xp33_ASAP7_75t_L g643 ( 
.A(n_544),
.B(n_421),
.C(n_419),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_584),
.B(n_400),
.Y(n_646)
);

BUFx8_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_548),
.B(n_402),
.Y(n_648)
);

BUFx2_ASAP7_75t_SL g649 ( 
.A(n_555),
.Y(n_649)
);

NAND2x1_ASAP7_75t_L g650 ( 
.A(n_585),
.B(n_403),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_548),
.B(n_404),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_565),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_560),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_649),
.B(n_589),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_L g655 ( 
.A1(n_596),
.A2(n_615),
.B1(n_612),
.B2(n_602),
.C(n_605),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_609),
.Y(n_656)
);

AO22x2_ASAP7_75t_L g657 ( 
.A1(n_603),
.A2(n_601),
.B1(n_594),
.B2(n_625),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_595),
.A2(n_580),
.B1(n_585),
.B2(n_579),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_623),
.B(n_568),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_599),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_621),
.B(n_568),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_606),
.A2(n_579),
.B1(n_590),
.B2(n_591),
.C(n_589),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_600),
.B(n_589),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_616),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_600),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_629),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_634),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_643),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_610),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_613),
.Y(n_673)
);

NAND2x1p5_ASAP7_75t_L g674 ( 
.A(n_641),
.B(n_591),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_641),
.B(n_159),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_607),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_620),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_406),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_631),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_647),
.Y(n_681)
);

OAI221xp5_ASAP7_75t_L g682 ( 
.A1(n_622),
.A2(n_624),
.B1(n_637),
.B2(n_633),
.C(n_617),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

NAND2x1p5_ASAP7_75t_L g684 ( 
.A(n_635),
.B(n_163),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_616),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_636),
.Y(n_686)
);

BUFx8_ASAP7_75t_L g687 ( 
.A(n_635),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_634),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_652),
.A2(n_11),
.B1(n_18),
.B2(n_5),
.Y(n_690)
);

AO22x2_ASAP7_75t_L g691 ( 
.A1(n_640),
.A2(n_12),
.B1(n_19),
.B2(n_6),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_597),
.A2(n_165),
.B1(n_166),
.B2(n_164),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_645),
.A2(n_653),
.B1(n_650),
.B2(n_611),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_636),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_638),
.B(n_6),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_638),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_627),
.B(n_7),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_644),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_683),
.A2(n_626),
.B1(n_630),
.B2(n_628),
.Y(n_700)
);

CKINVDCx8_ASAP7_75t_R g701 ( 
.A(n_654),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_664),
.A2(n_651),
.B(n_648),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_682),
.A2(n_632),
.B(n_614),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_646),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_659),
.B(n_7),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_655),
.A2(n_169),
.B(n_167),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_661),
.B(n_8),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_687),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_663),
.A2(n_171),
.B(n_170),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_679),
.A2(n_173),
.B(n_172),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_658),
.A2(n_175),
.B(n_174),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_666),
.B(n_10),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_670),
.B(n_13),
.Y(n_713)
);

BUFx8_ASAP7_75t_L g714 ( 
.A(n_665),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_698),
.B(n_14),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_667),
.B(n_176),
.Y(n_716)
);

AOI21x1_ASAP7_75t_L g717 ( 
.A1(n_693),
.A2(n_179),
.B(n_178),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_657),
.A2(n_680),
.B1(n_668),
.B2(n_678),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_667),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_669),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_15),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_672),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_674),
.A2(n_181),
.B(n_180),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_673),
.B(n_17),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_675),
.B(n_183),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_695),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_657),
.B(n_17),
.Y(n_727)
);

CKINVDCx10_ASAP7_75t_R g728 ( 
.A(n_689),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_699),
.B(n_184),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_688),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_694),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_660),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_686),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_697),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_696),
.B(n_22),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_662),
.A2(n_187),
.B(n_186),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_681),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_676),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_L g739 ( 
.A1(n_671),
.A2(n_25),
.B(n_26),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_692),
.A2(n_189),
.B(n_188),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_677),
.B(n_27),
.C(n_28),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_691),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_728),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_740),
.A2(n_690),
.B(n_31),
.C(n_29),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_718),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_715),
.B(n_30),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_704),
.B(n_700),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_732),
.B(n_190),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_722),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_727),
.B(n_32),
.Y(n_751)
);

CKINVDCx16_ASAP7_75t_R g752 ( 
.A(n_708),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_719),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_743),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_733),
.B(n_191),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_734),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_712),
.B(n_33),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_721),
.B(n_739),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_713),
.B(n_35),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_719),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_720),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_705),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_707),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_724),
.B(n_737),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_735),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_711),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_741),
.B(n_703),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_741),
.B(n_192),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_716),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_701),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_714),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_738),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_730),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_725),
.B(n_193),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_40),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_706),
.B(n_40),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_710),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_723),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_731),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_702),
.B(n_41),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_736),
.B(n_42),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_709),
.B(n_43),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_726),
.B(n_44),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

OR2x2_ASAP7_75t_SL g787 ( 
.A(n_752),
.B(n_44),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_786),
.B(n_194),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_762),
.B(n_46),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_748),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_764),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_744),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_770),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_758),
.B(n_47),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_770),
.Y(n_795)
);

NOR2x1_ASAP7_75t_SL g796 ( 
.A(n_767),
.B(n_769),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_754),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_780),
.A2(n_315),
.B(n_314),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_776),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_751),
.B(n_50),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_778),
.A2(n_196),
.B(n_195),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_763),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_761),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_760),
.B(n_197),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_782),
.A2(n_313),
.B(n_311),
.Y(n_805)
);

BUFx2_ASAP7_75t_R g806 ( 
.A(n_771),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_779),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_807)
);

AOI221x1_ASAP7_75t_L g808 ( 
.A1(n_777),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.C(n_57),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_765),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_757),
.B(n_58),
.Y(n_810)
);

AOI221xp5_ASAP7_75t_L g811 ( 
.A1(n_775),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.C(n_63),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_756),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_768),
.B(n_198),
.Y(n_813)
);

O2A1O1Ixp5_ASAP7_75t_SL g814 ( 
.A1(n_772),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_759),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_785),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_755),
.B(n_199),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_784),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_747),
.B(n_67),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_773),
.B(n_781),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_749),
.B(n_200),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_774),
.A2(n_783),
.B(n_746),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_786),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_767),
.A2(n_202),
.B(n_201),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_750),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_753),
.Y(n_826)
);

NOR2x1_ASAP7_75t_L g827 ( 
.A(n_748),
.B(n_203),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_750),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_745),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.C(n_71),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_770),
.B(n_204),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_770),
.B(n_205),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_SL g832 ( 
.A1(n_766),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_770),
.B(n_206),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_750),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_744),
.Y(n_835)
);

NOR2x2_ASAP7_75t_L g836 ( 
.A(n_831),
.B(n_72),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_794),
.B(n_207),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_791),
.B(n_73),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_796),
.A2(n_209),
.B(n_208),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_822),
.A2(n_211),
.B(n_210),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_826),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_829),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_820),
.B(n_212),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_816),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_78),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_818),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_802),
.B(n_80),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_809),
.B(n_214),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_835),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_SL g850 ( 
.A(n_806),
.B(n_81),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_827),
.B(n_216),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_797),
.Y(n_852)
);

OA21x2_ASAP7_75t_L g853 ( 
.A1(n_808),
.A2(n_84),
.B(n_85),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_832),
.A2(n_87),
.B(n_88),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_819),
.B(n_218),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_825),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_828),
.Y(n_857)
);

OA22x2_ASAP7_75t_L g858 ( 
.A1(n_807),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_834),
.B(n_90),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_812),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_800),
.B(n_220),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_795),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_793),
.B(n_221),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_789),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_813),
.B(n_222),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_805),
.A2(n_91),
.B(n_92),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_810),
.B(n_223),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_792),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_811),
.B(n_790),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_799),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_801),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_817),
.B(n_92),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_787),
.B(n_93),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_821),
.B(n_94),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_830),
.B(n_833),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_798),
.A2(n_225),
.B(n_224),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_795),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_804),
.B(n_788),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_814),
.B(n_95),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_824),
.A2(n_96),
.B(n_97),
.Y(n_880)
);

OA22x2_ASAP7_75t_L g881 ( 
.A1(n_823),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_803),
.B(n_226),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_858),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_883)
);

AOI211xp5_ASAP7_75t_L g884 ( 
.A1(n_842),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_868),
.Y(n_885)
);

INVx4_ASAP7_75t_SL g886 ( 
.A(n_882),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_853),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_853),
.A2(n_865),
.B1(n_881),
.B2(n_854),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_873),
.A2(n_850),
.B1(n_864),
.B2(n_874),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_840),
.A2(n_108),
.B1(n_105),
.B2(n_106),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_846),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_860),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_856),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_867),
.A2(n_851),
.B1(n_843),
.B2(n_837),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_843),
.A2(n_112),
.B1(n_109),
.B2(n_111),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_866),
.A2(n_880),
.B1(n_879),
.B2(n_878),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_841),
.B(n_111),
.Y(n_897)
);

BUFx4f_ASAP7_75t_SL g898 ( 
.A(n_877),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_870),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_855),
.B(n_113),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_875),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_861),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_871),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_849),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_872),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_845),
.A2(n_847),
.B1(n_838),
.B2(n_859),
.Y(n_906)
);

BUFx4f_ASAP7_75t_SL g907 ( 
.A(n_863),
.Y(n_907)
);

BUFx4f_ASAP7_75t_SL g908 ( 
.A(n_863),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_836),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_848),
.B(n_121),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_839),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_876),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_862),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_857),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_852),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_844),
.B(n_130),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_869),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_852),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_869),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_891),
.B(n_140),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_909),
.B(n_141),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_899),
.Y(n_923)
);

BUFx4f_ASAP7_75t_SL g924 ( 
.A(n_885),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_915),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_903),
.B(n_143),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_901),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_917),
.B(n_146),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_884),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_892),
.B(n_914),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_919),
.B(n_149),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_898),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_911),
.B(n_229),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_900),
.Y(n_934)
);

BUFx12f_ASAP7_75t_L g935 ( 
.A(n_904),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_910),
.A2(n_151),
.B(n_152),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_906),
.B(n_151),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_893),
.B(n_154),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_886),
.B(n_155),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_913),
.B(n_157),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_923),
.B(n_916),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_897),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_925),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_930),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_934),
.B(n_889),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_928),
.B(n_931),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_929),
.A2(n_888),
.B1(n_887),
.B2(n_883),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_926),
.B(n_894),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_935),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_932),
.B(n_896),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_921),
.B(n_905),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_936),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_938),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_937),
.B(n_912),
.C(n_890),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_939),
.B(n_895),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_940),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_933),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_922),
.B(n_902),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_949),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_924),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_952),
.B(n_907),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_908),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_943),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_944),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_941),
.B(n_920),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_946),
.B(n_918),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_942),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_967),
.B(n_945),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_953),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_962),
.B(n_956),
.Y(n_970)
);

AND2x4_ASAP7_75t_SL g971 ( 
.A(n_961),
.B(n_948),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_951),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_960),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_959),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_965),
.B(n_955),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_973),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_975),
.Y(n_978)
);

AOI31xp33_ASAP7_75t_L g979 ( 
.A1(n_974),
.A2(n_954),
.A3(n_947),
.B(n_958),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_976),
.B(n_966),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_979),
.A2(n_971),
.B(n_972),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_978),
.B(n_971),
.Y(n_982)
);

AND3x1_ASAP7_75t_L g983 ( 
.A(n_982),
.B(n_980),
.C(n_977),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_981),
.B(n_969),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_984),
.B(n_970),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_985),
.B(n_983),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_986),
.B(n_968),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_987),
.B(n_238),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_988),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_989),
.B(n_245),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_990),
.B(n_248),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_991),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_992),
.Y(n_993)
);

AOI322xp5_ASAP7_75t_L g994 ( 
.A1(n_993),
.A2(n_250),
.A3(n_251),
.B1(n_252),
.B2(n_253),
.C1(n_254),
.C2(n_255),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_994),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_L g996 ( 
.A(n_995),
.B(n_258),
.C(n_259),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_996),
.A2(n_260),
.B1(n_262),
.B2(n_264),
.Y(n_997)
);

OAI322xp33_ASAP7_75t_L g998 ( 
.A1(n_997),
.A2(n_265),
.A3(n_266),
.B1(n_267),
.B2(n_270),
.C1(n_271),
.C2(n_272),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_998),
.B(n_273),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_999),
.B(n_274),
.Y(n_1000)
);

AOI22x1_ASAP7_75t_L g1001 ( 
.A1(n_1000),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_1001),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.C(n_284),
.Y(n_1002)
);

AOI211xp5_ASAP7_75t_L g1003 ( 
.A1(n_1002),
.A2(n_286),
.B(n_287),
.C(n_288),
.Y(n_1003)
);


endmodule