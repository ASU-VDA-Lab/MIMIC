module fake_jpeg_25562_n_41 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_4),
.B(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_11),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_6),
.B1(n_16),
.B2(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_30),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_30),
.C(n_17),
.Y(n_36)
);

XOR2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.C(n_33),
.Y(n_38)
);

OAI21x1_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_34),
.B(n_14),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_20),
.A3(n_19),
.B1(n_15),
.B2(n_28),
.C(n_29),
.Y(n_41)
);


endmodule