module real_aes_319_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g507 ( .A(n_0), .B(n_199), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_1), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g133 ( .A(n_2), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_3), .B(n_510), .Y(n_529) );
NAND2xp33_ASAP7_75t_SL g500 ( .A(n_4), .B(n_154), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_5), .B(n_167), .Y(n_190) );
INVx1_ASAP7_75t_L g492 ( .A(n_6), .Y(n_492) );
INVx1_ASAP7_75t_L g224 ( .A(n_7), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g815 ( .A(n_8), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_9), .Y(n_241) );
AND2x2_ASAP7_75t_L g527 ( .A(n_10), .B(n_123), .Y(n_527) );
INVx2_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_12), .Y(n_478) );
INVx1_ASAP7_75t_L g200 ( .A(n_13), .Y(n_200) );
AOI221x1_ASAP7_75t_L g495 ( .A1(n_14), .A2(n_156), .B1(n_496), .B2(n_498), .C(n_499), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_15), .B(n_510), .Y(n_563) );
INVx1_ASAP7_75t_L g481 ( .A(n_16), .Y(n_481) );
NOR2xp33_ASAP7_75t_SL g812 ( .A(n_16), .B(n_482), .Y(n_812) );
INVx1_ASAP7_75t_L g197 ( .A(n_17), .Y(n_197) );
INVx1_ASAP7_75t_SL g145 ( .A(n_18), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_19), .B(n_148), .Y(n_170) );
AOI33xp33_ASAP7_75t_L g215 ( .A1(n_20), .A2(n_50), .A3(n_130), .B1(n_141), .B2(n_216), .B3(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_21), .A2(n_498), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_22), .B(n_199), .Y(n_532) );
AOI221xp5_ASAP7_75t_SL g572 ( .A1(n_23), .A2(n_41), .B1(n_498), .B2(n_510), .C(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g234 ( .A(n_24), .Y(n_234) );
OR2x2_ASAP7_75t_L g125 ( .A(n_25), .B(n_90), .Y(n_125) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_25), .A2(n_90), .B(n_124), .Y(n_158) );
INVxp67_ASAP7_75t_L g494 ( .A(n_26), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_27), .B(n_202), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_28), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g521 ( .A(n_29), .B(n_122), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_30), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_31), .B(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_32), .A2(n_103), .B1(n_809), .B2(n_816), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_33), .A2(n_498), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_34), .B(n_202), .Y(n_574) );
AND2x2_ASAP7_75t_L g135 ( .A(n_35), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g140 ( .A(n_35), .Y(n_140) );
AND2x2_ASAP7_75t_L g154 ( .A(n_35), .B(n_133), .Y(n_154) );
OR2x6_ASAP7_75t_L g479 ( .A(n_36), .B(n_480), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_36), .B(n_478), .C(n_814), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_37), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_38), .B(n_128), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_39), .A2(n_157), .B1(n_163), .B2(n_167), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_40), .B(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_42), .A2(n_82), .B1(n_138), .B2(n_498), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_43), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_44), .B(n_199), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_45), .B(n_174), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_46), .B(n_148), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_47), .Y(n_166) );
AND2x2_ASAP7_75t_L g511 ( .A(n_48), .B(n_122), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_49), .B(n_122), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_51), .B(n_148), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_52), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_52), .A2(n_62), .B1(n_413), .B2(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g131 ( .A(n_53), .Y(n_131) );
INVx1_ASAP7_75t_L g150 ( .A(n_53), .Y(n_150) );
AND2x2_ASAP7_75t_L g266 ( .A(n_54), .B(n_122), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g222 ( .A1(n_55), .A2(n_75), .B1(n_128), .B2(n_138), .C(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_56), .B(n_128), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_57), .B(n_510), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_58), .B(n_157), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g179 ( .A1(n_59), .A2(n_138), .B(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g548 ( .A(n_60), .B(n_122), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_61), .B(n_202), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_62), .Y(n_804) );
INVx1_ASAP7_75t_L g193 ( .A(n_63), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_64), .B(n_199), .Y(n_546) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_65), .B(n_123), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_66), .A2(n_498), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g264 ( .A(n_67), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_68), .B(n_202), .Y(n_533) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_69), .B(n_174), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_70), .A2(n_101), .B1(n_777), .B2(n_778), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_70), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_71), .A2(n_138), .B(n_263), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_72), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_72), .Y(n_802) );
INVx1_ASAP7_75t_L g136 ( .A(n_73), .Y(n_136) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_74), .B(n_128), .Y(n_218) );
AND2x2_ASAP7_75t_L g155 ( .A(n_76), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g194 ( .A(n_77), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_78), .A2(n_138), .B(n_144), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_79), .A2(n_138), .B(n_169), .C(n_173), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_80), .A2(n_85), .B1(n_128), .B2(n_510), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_81), .B(n_510), .Y(n_547) );
INVx1_ASAP7_75t_L g482 ( .A(n_83), .Y(n_482) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_84), .B(n_156), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_86), .A2(n_138), .B1(n_213), .B2(n_214), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_87), .B(n_199), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_88), .B(n_199), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_89), .A2(n_498), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g181 ( .A(n_91), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_92), .B(n_202), .Y(n_545) );
AND2x2_ASAP7_75t_L g219 ( .A(n_93), .B(n_156), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_94), .A2(n_232), .B(n_233), .C(n_235), .Y(n_231) );
INVxp67_ASAP7_75t_L g497 ( .A(n_95), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_96), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_97), .B(n_202), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_98), .A2(n_498), .B(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_SL g106 ( .A(n_99), .Y(n_106) );
BUFx2_ASAP7_75t_L g789 ( .A(n_99), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_100), .B(n_148), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_101), .Y(n_778) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B(n_786), .Y(n_103) );
CKINVDCx11_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx8_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_783), .Y(n_107) );
AOI21xp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_775), .B(n_779), .Y(n_108) );
OAI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_476), .B1(n_483), .B2(n_771), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_111), .A2(n_476), .B1(n_484), .B2(n_785), .Y(n_784) );
AND3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_470), .C(n_473), .Y(n_111) );
NAND5xp2_ASAP7_75t_L g112 ( .A(n_113), .B(n_370), .C(n_400), .D(n_414), .E(n_440), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_114), .A2(n_413), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g798 ( .A(n_114), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_319), .Y(n_114) );
NOR3xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_267), .C(n_301), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_184), .B(n_206), .C(n_245), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_159), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_119), .B(n_257), .Y(n_322) );
AND2x2_ASAP7_75t_L g409 ( .A(n_119), .B(n_187), .Y(n_409) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g205 ( .A(n_120), .B(n_176), .Y(n_205) );
INVx1_ASAP7_75t_L g247 ( .A(n_120), .Y(n_247) );
INVx2_ASAP7_75t_L g252 ( .A(n_120), .Y(n_252) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_120), .Y(n_280) );
INVx1_ASAP7_75t_L g294 ( .A(n_120), .Y(n_294) );
AND2x2_ASAP7_75t_L g298 ( .A(n_120), .B(n_189), .Y(n_298) );
AND2x2_ASAP7_75t_L g379 ( .A(n_120), .B(n_188), .Y(n_379) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_126), .B(n_155), .Y(n_120) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_121), .A2(n_515), .B(n_521), .Y(n_514) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_121), .A2(n_542), .B(n_548), .Y(n_541) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_121), .A2(n_515), .B(n_521), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_122), .A2(n_572), .B(n_576), .Y(n_571) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x4_ASAP7_75t_L g167 ( .A(n_124), .B(n_125), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_137), .Y(n_126) );
INVx1_ASAP7_75t_L g244 ( .A(n_128), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_128), .A2(n_138), .B1(n_491), .B2(n_493), .Y(n_490) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_134), .Y(n_128) );
INVx1_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
OR2x6_ASAP7_75t_L g146 ( .A(n_130), .B(n_142), .Y(n_146) );
INVxp33_ASAP7_75t_L g216 ( .A(n_130), .Y(n_216) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g143 ( .A(n_131), .B(n_133), .Y(n_143) );
AND2x4_ASAP7_75t_L g202 ( .A(n_131), .B(n_151), .Y(n_202) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g498 ( .A(n_135), .B(n_143), .Y(n_498) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
AND2x6_ASAP7_75t_L g199 ( .A(n_136), .B(n_149), .Y(n_199) );
INVxp67_ASAP7_75t_L g242 ( .A(n_138), .Y(n_242) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NOR2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx1_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_146), .B(n_147), .C(n_153), .Y(n_144) );
INVx2_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_153), .B(n_181), .C(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_146), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_146), .A2(n_153), .B(n_224), .C(n_225), .Y(n_223) );
INVxp67_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_146), .A2(n_153), .B(n_264), .C(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
AND2x4_ASAP7_75t_L g510 ( .A(n_148), .B(n_154), .Y(n_510) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_153), .A2(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_153), .B(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_153), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_153), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_153), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_153), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_153), .A2(n_566), .B(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_153), .A2(n_574), .B(n_575), .Y(n_573) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_154), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_156), .A2(n_231), .B1(n_236), .B2(n_237), .Y(n_230) );
INVx3_ASAP7_75t_L g237 ( .A(n_156), .Y(n_237) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_157), .B(n_240), .Y(n_239) );
AOI21x1_ASAP7_75t_L g503 ( .A1(n_157), .A2(n_504), .B(n_511), .Y(n_503) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
AND2x4_ASAP7_75t_SL g159 ( .A(n_160), .B(n_175), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
AND2x2_ASAP7_75t_L g248 ( .A(n_161), .B(n_189), .Y(n_248) );
AND2x2_ASAP7_75t_L g269 ( .A(n_161), .B(n_176), .Y(n_269) );
INVx1_ASAP7_75t_L g292 ( .A(n_161), .Y(n_292) );
AND2x4_ASAP7_75t_L g359 ( .A(n_161), .B(n_188), .Y(n_359) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_168), .Y(n_161) );
NOR3xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .C(n_166), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_167), .A2(n_179), .B(n_183), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_167), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_167), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_167), .B(n_497), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g499 ( .A(n_167), .B(n_195), .C(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_167), .A2(n_529), .B(n_530), .Y(n_528) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_211), .B(n_219), .Y(n_210) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_173), .A2(n_211), .B(n_219), .Y(n_274) );
AOI21x1_ASAP7_75t_L g536 ( .A1(n_173), .A2(n_537), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_174), .A2(n_222), .B(n_226), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_174), .A2(n_563), .B(n_564), .Y(n_562) );
AND2x4_ASAP7_75t_L g375 ( .A(n_175), .B(n_292), .Y(n_375) );
OR2x2_ASAP7_75t_L g416 ( .A(n_175), .B(n_417), .Y(n_416) );
NOR2xp67_ASAP7_75t_SL g435 ( .A(n_175), .B(n_308), .Y(n_435) );
NOR2x1_ASAP7_75t_L g453 ( .A(n_175), .B(n_367), .Y(n_453) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2x1_ASAP7_75t_SL g253 ( .A(n_176), .B(n_189), .Y(n_253) );
AND2x4_ASAP7_75t_L g291 ( .A(n_176), .B(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_176), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_176), .B(n_251), .Y(n_329) );
INVx2_ASAP7_75t_L g343 ( .A(n_176), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_176), .B(n_295), .Y(n_365) );
AND2x2_ASAP7_75t_L g457 ( .A(n_176), .B(n_315), .Y(n_457) );
OR2x6_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2x1_ASAP7_75t_L g185 ( .A(n_186), .B(n_205), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_187), .B(n_294), .Y(n_308) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_187), .B(n_297), .Y(n_317) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_204), .Y(n_187) );
INVx1_ASAP7_75t_L g295 ( .A(n_188), .Y(n_295) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g315 ( .A(n_189), .Y(n_315) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_196), .B(n_203), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_195), .B(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B1(n_200), .B2(n_201), .Y(n_196) );
INVxp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVxp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g348 ( .A(n_204), .Y(n_348) );
INVx2_ASAP7_75t_SL g393 ( .A(n_205), .Y(n_393) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_227), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_208), .B(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g339 ( .A(n_208), .Y(n_339) );
AND2x2_ASAP7_75t_L g463 ( .A(n_208), .B(n_288), .Y(n_463) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AND2x4_ASAP7_75t_L g276 ( .A(n_209), .B(n_258), .Y(n_276) );
INVx1_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
AND2x2_ASAP7_75t_L g318 ( .A(n_209), .B(n_273), .Y(n_318) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_210), .B(n_221), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_210), .B(n_259), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_212), .B(n_218), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g256 ( .A(n_221), .Y(n_256) );
AND2x4_ASAP7_75t_L g324 ( .A(n_221), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g336 ( .A(n_221), .Y(n_336) );
INVx1_ASAP7_75t_L g378 ( .A(n_221), .Y(n_378) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_221), .Y(n_390) );
AND2x2_ASAP7_75t_L g406 ( .A(n_221), .B(n_229), .Y(n_406) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g353 ( .A(n_228), .B(n_311), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_228), .Y(n_355) );
AND2x2_ASAP7_75t_L g376 ( .A(n_228), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g255 ( .A(n_229), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g283 ( .A(n_229), .Y(n_283) );
INVx2_ASAP7_75t_L g289 ( .A(n_229), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_229), .B(n_259), .Y(n_304) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_238), .Y(n_229) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_237), .A2(n_260), .B(n_266), .Y(n_259) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_237), .A2(n_260), .B(n_266), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_242), .B1(n_243), .B2(n_244), .Y(n_238) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B(n_254), .Y(n_245) );
INVx1_ASAP7_75t_L g385 ( .A(n_246), .Y(n_385) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g305 ( .A(n_248), .Y(n_305) );
AND2x2_ASAP7_75t_L g361 ( .A(n_248), .B(n_297), .Y(n_361) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g275 ( .A(n_250), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_250), .B(n_291), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_250), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_250), .B(n_375), .Y(n_382) );
AND2x2_ASAP7_75t_L g456 ( .A(n_250), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_251), .Y(n_444) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_252), .Y(n_364) );
AND2x2_ASAP7_75t_L g277 ( .A(n_253), .B(n_278), .Y(n_277) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_253), .A2(n_466), .B(n_468), .Y(n_465) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx3_ASAP7_75t_L g351 ( .A(n_255), .Y(n_351) );
NAND2x1_ASAP7_75t_SL g395 ( .A(n_255), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_255), .B(n_276), .Y(n_398) );
AND2x2_ASAP7_75t_L g310 ( .A(n_257), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g447 ( .A(n_257), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g458 ( .A(n_257), .B(n_406), .Y(n_458) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_258), .B(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g389 ( .A(n_259), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OAI21xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_281), .B(n_284), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B1(n_276), .B2(n_277), .Y(n_268) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_269), .Y(n_326) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
AND2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g405 ( .A(n_271), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_271), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_271), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g288 ( .A(n_273), .B(n_289), .Y(n_288) );
NOR2xp67_ASAP7_75t_L g369 ( .A(n_273), .B(n_289), .Y(n_369) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_273), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
AND2x2_ASAP7_75t_L g333 ( .A(n_274), .B(n_289), .Y(n_333) );
INVx1_ASAP7_75t_L g396 ( .A(n_274), .Y(n_396) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_279), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g426 ( .A(n_282), .B(n_311), .Y(n_426) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g300 ( .A(n_283), .Y(n_300) );
AND2x2_ASAP7_75t_L g323 ( .A(n_283), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g411 ( .A(n_283), .B(n_318), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .B1(n_296), .B2(n_299), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g419 ( .A(n_286), .B(n_420), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g449 ( .A(n_289), .B(n_336), .Y(n_449) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g316 ( .A(n_291), .Y(n_316) );
OAI21xp33_ASAP7_75t_SL g462 ( .A1(n_291), .A2(n_463), .B(n_464), .Y(n_462) );
AND2x4_ASAP7_75t_SL g293 ( .A(n_294), .B(n_295), .Y(n_293) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_294), .Y(n_452) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_SL g394 ( .A1(n_297), .A2(n_395), .B(n_397), .C(n_399), .Y(n_394) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_298), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g399 ( .A(n_298), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_298), .B(n_375), .Y(n_439) );
INVx1_ASAP7_75t_SL g306 ( .A(n_299), .Y(n_306) );
AND2x2_ASAP7_75t_L g387 ( .A(n_300), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g432 ( .A(n_300), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_306), .B2(n_307), .C(n_309), .Y(n_301) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_302), .Y(n_421) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g469 ( .A(n_304), .B(n_312), .Y(n_469) );
OR2x2_ASAP7_75t_L g328 ( .A(n_305), .B(n_329), .Y(n_328) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_305), .B(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_305), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g467 ( .A(n_305), .B(n_364), .Y(n_467) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI32xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .A3(n_316), .B1(n_317), .B2(n_318), .Y(n_309) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_313), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g425 ( .A(n_314), .Y(n_425) );
OAI22xp33_ASAP7_75t_SL g407 ( .A1(n_316), .A2(n_408), .B1(n_410), .B2(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g438 ( .A(n_317), .Y(n_438) );
AOI211x1_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_326), .B(n_327), .C(n_344), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_321), .B(n_406), .Y(n_412) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g368 ( .A(n_324), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g434 ( .A(n_324), .Y(n_434) );
OAI222xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_331), .B2(n_337), .C1(n_338), .C2(n_340), .Y(n_327) );
INVxp67_ASAP7_75t_L g424 ( .A(n_328), .Y(n_424) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_332), .B(n_417), .Y(n_464) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g380 ( .A(n_333), .B(n_377), .Y(n_380) );
INVx3_ASAP7_75t_L g420 ( .A(n_335), .Y(n_420) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g358 ( .A(n_343), .B(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B1(n_352), .B2(n_357), .C(n_360), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_346), .A2(n_403), .B(n_405), .Y(n_402) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g356 ( .A(n_350), .Y(n_356) );
OR2x2_ASAP7_75t_L g460 ( .A(n_351), .B(n_396), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_354), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_357), .A2(n_386), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_358), .A2(n_430), .B(n_437), .Y(n_436) );
INVx4_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
OAI31xp33_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .A3(n_366), .B(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g392 ( .A(n_367), .Y(n_392) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_383), .Y(n_370) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_371), .B(n_383), .C(n_402), .D(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_381), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_379), .B2(n_380), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g443 ( .A(n_375), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_376), .B(n_396), .Y(n_404) );
INVx1_ASAP7_75t_SL g417 ( .A(n_379), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_394), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_388), .B2(n_391), .Y(n_384) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_393), .A2(n_456), .B1(n_458), .B2(n_459), .Y(n_455) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_407), .C(n_413), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g472 ( .A(n_407), .Y(n_472) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g473 ( .A1(n_413), .A2(n_474), .B(n_475), .Y(n_473) );
INVxp33_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
AND2x2_ASAP7_75t_L g797 ( .A(n_414), .B(n_440), .Y(n_797) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_415), .B(n_422), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_419), .B2(n_421), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_419), .A2(n_442), .B(n_445), .Y(n_441) );
INVx2_ASAP7_75t_L g429 ( .A(n_420), .Y(n_429) );
NAND3xp33_ASAP7_75t_SL g422 ( .A(n_423), .B(n_427), .C(n_436), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_433), .B2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVxp33_ASAP7_75t_SL g475 ( .A(n_440), .Y(n_475) );
NOR3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_454), .C(n_461), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g799 ( .A(n_471), .Y(n_799) );
CKINVDCx11_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OR2x6_ASAP7_75t_SL g773 ( .A(n_478), .B(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g782 ( .A(n_478), .B(n_479), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_478), .B(n_774), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_479), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_648), .Y(n_484) );
NOR4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_591), .C(n_630), .D(n_637), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_512), .B1(n_549), .B2(n_558), .C(n_577), .Y(n_486) );
OR2x2_ASAP7_75t_L g721 ( .A(n_487), .B(n_583), .Y(n_721) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g636 ( .A(n_488), .B(n_561), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_488), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_SL g701 ( .A(n_488), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_501), .Y(n_488) );
AND2x4_ASAP7_75t_SL g560 ( .A(n_489), .B(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g582 ( .A(n_489), .Y(n_582) );
AND2x2_ASAP7_75t_L g617 ( .A(n_489), .B(n_590), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_489), .B(n_502), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_489), .B(n_584), .Y(n_669) );
OR2x2_ASAP7_75t_L g747 ( .A(n_489), .B(n_561), .Y(n_747) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_502), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g595 ( .A(n_502), .Y(n_595) );
OR2x2_ASAP7_75t_L g600 ( .A(n_502), .B(n_584), .Y(n_600) );
AND2x2_ASAP7_75t_L g613 ( .A(n_502), .B(n_571), .Y(n_613) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_502), .Y(n_616) );
INVx1_ASAP7_75t_L g628 ( .A(n_502), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_502), .B(n_582), .Y(n_693) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_513), .B(n_522), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g557 ( .A(n_514), .B(n_541), .Y(n_557) );
AND2x4_ASAP7_75t_L g587 ( .A(n_514), .B(n_526), .Y(n_587) );
INVx2_ASAP7_75t_L g621 ( .A(n_514), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_514), .B(n_541), .Y(n_679) );
AND2x2_ASAP7_75t_L g726 ( .A(n_514), .B(n_555), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g714 ( .A1(n_522), .A2(n_586), .B1(n_629), .B2(n_689), .C1(n_715), .C2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .Y(n_523) );
AND2x2_ASAP7_75t_L g633 ( .A(n_524), .B(n_553), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_524), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g762 ( .A(n_524), .B(n_602), .Y(n_762) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_525), .A2(n_593), .B(n_597), .Y(n_592) );
AND2x2_ASAP7_75t_L g673 ( .A(n_525), .B(n_556), .Y(n_673) );
OR2x2_ASAP7_75t_L g698 ( .A(n_525), .B(n_557), .Y(n_698) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx5_ASAP7_75t_L g552 ( .A(n_526), .Y(n_552) );
AND2x2_ASAP7_75t_L g639 ( .A(n_526), .B(n_621), .Y(n_639) );
AND2x2_ASAP7_75t_L g665 ( .A(n_526), .B(n_541), .Y(n_665) );
OR2x2_ASAP7_75t_L g668 ( .A(n_526), .B(n_555), .Y(n_668) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_526), .Y(n_686) );
AND2x4_ASAP7_75t_SL g743 ( .A(n_526), .B(n_620), .Y(n_743) );
OR2x2_ASAP7_75t_L g752 ( .A(n_526), .B(n_579), .Y(n_752) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g585 ( .A(n_534), .Y(n_585) );
AOI221xp5_ASAP7_75t_SL g703 ( .A1(n_534), .A2(n_587), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_703) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_541), .Y(n_534) );
OR2x2_ASAP7_75t_L g642 ( .A(n_535), .B(n_612), .Y(n_642) );
OR2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g678 ( .A(n_535), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g684 ( .A(n_535), .B(n_603), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_535), .B(n_667), .Y(n_696) );
INVx2_ASAP7_75t_L g709 ( .A(n_535), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_535), .B(n_587), .Y(n_730) );
AND2x2_ASAP7_75t_L g734 ( .A(n_535), .B(n_556), .Y(n_734) );
AND2x2_ASAP7_75t_L g742 ( .A(n_535), .B(n_743), .Y(n_742) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g555 ( .A(n_536), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_541), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g586 ( .A(n_541), .B(n_555), .Y(n_586) );
INVx2_ASAP7_75t_L g603 ( .A(n_541), .Y(n_603) );
AND2x4_ASAP7_75t_L g620 ( .A(n_541), .B(n_621), .Y(n_620) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_541), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g732 ( .A(n_551), .B(n_554), .Y(n_732) );
AND2x4_ASAP7_75t_L g578 ( .A(n_552), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g619 ( .A(n_552), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_586), .Y(n_646) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g750 ( .A(n_554), .B(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g602 ( .A(n_555), .B(n_603), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_556), .A2(n_623), .B(n_629), .Y(n_622) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_569), .Y(n_559) );
INVx1_ASAP7_75t_SL g676 ( .A(n_560), .Y(n_676) );
AND2x2_ASAP7_75t_L g706 ( .A(n_560), .B(n_616), .Y(n_706) );
AND2x4_ASAP7_75t_L g717 ( .A(n_560), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g583 ( .A(n_561), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g590 ( .A(n_561), .Y(n_590) );
AND2x4_ASAP7_75t_L g596 ( .A(n_561), .B(n_582), .Y(n_596) );
INVx2_ASAP7_75t_L g607 ( .A(n_561), .Y(n_607) );
INVx1_ASAP7_75t_L g656 ( .A(n_561), .Y(n_656) );
OR2x2_ASAP7_75t_L g677 ( .A(n_561), .B(n_661), .Y(n_677) );
OR2x2_ASAP7_75t_L g691 ( .A(n_561), .B(n_571), .Y(n_691) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_561), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_561), .B(n_613), .Y(n_763) );
OR2x6_ASAP7_75t_L g561 ( .A(n_562), .B(n_568), .Y(n_561) );
INVx1_ASAP7_75t_L g608 ( .A(n_569), .Y(n_608) );
AND2x2_ASAP7_75t_L g741 ( .A(n_569), .B(n_607), .Y(n_741) );
AND2x2_ASAP7_75t_L g766 ( .A(n_569), .B(n_596), .Y(n_766) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g584 ( .A(n_571), .Y(n_584) );
BUFx3_ASAP7_75t_L g626 ( .A(n_571), .Y(n_626) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_571), .Y(n_653) );
INVx1_ASAP7_75t_L g662 ( .A(n_571), .Y(n_662) );
AOI33xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .A3(n_585), .B1(n_586), .B2(n_587), .B3(n_588), .Y(n_577) );
AOI21x1_ASAP7_75t_SL g680 ( .A1(n_578), .A2(n_602), .B(n_664), .Y(n_680) );
INVx2_ASAP7_75t_L g710 ( .A(n_578), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_578), .B(n_709), .Y(n_716) );
AND2x2_ASAP7_75t_L g664 ( .A(n_579), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g627 ( .A(n_582), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g728 ( .A(n_583), .Y(n_728) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_584), .Y(n_718) );
OAI32xp33_ASAP7_75t_L g767 ( .A1(n_585), .A2(n_587), .A3(n_763), .B1(n_768), .B2(n_770), .Y(n_767) );
AND2x2_ASAP7_75t_L g685 ( .A(n_586), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g675 ( .A(n_587), .Y(n_675) );
AND2x2_ASAP7_75t_L g740 ( .A(n_587), .B(n_684), .Y(n_740) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_601), .B1(n_604), .B2(n_618), .C(n_622), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_595), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_596), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_596), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_596), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g645 ( .A(n_600), .Y(n_645) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .C(n_614), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_606), .A2(n_668), .B1(n_708), .B2(n_711), .Y(n_707) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g611 ( .A(n_607), .Y(n_611) );
NOR2x1p5_ASAP7_75t_L g625 ( .A(n_607), .B(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_607), .Y(n_647) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_610), .A2(n_652), .A3(n_675), .B1(n_676), .B2(n_677), .C1(n_678), .C2(n_680), .Y(n_674) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_612), .A2(n_631), .B(n_632), .C(n_634), .Y(n_630) );
OR2x2_ASAP7_75t_L g722 ( .A(n_612), .B(n_676), .Y(n_722) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g629 ( .A(n_613), .B(n_617), .Y(n_629) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g635 ( .A(n_619), .B(n_636), .Y(n_635) );
INVx3_ASAP7_75t_SL g667 ( .A(n_620), .Y(n_667) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_624), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_SL g671 ( .A(n_627), .Y(n_671) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_628), .Y(n_713) );
OR2x6_ASAP7_75t_SL g768 ( .A(n_631), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g758 ( .A1(n_636), .A2(n_759), .B(n_760), .C(n_767), .Y(n_758) );
O2A1O1Ixp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_643), .C(n_647), .Y(n_637) );
OAI211xp5_ASAP7_75t_SL g649 ( .A1(n_638), .A2(n_650), .B(n_657), .C(n_681), .Y(n_649) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_694), .C(n_738), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_653), .Y(n_745) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g700 ( .A(n_656), .Y(n_700) );
NOR3xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_670), .C(n_674), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_663), .B1(n_666), .B2(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g702 ( .A(n_662), .Y(n_702) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_662), .Y(n_769) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_SL g755 ( .A(n_668), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OR2x2_ASAP7_75t_L g705 ( .A(n_671), .B(n_691), .Y(n_705) );
OR2x2_ASAP7_75t_L g756 ( .A(n_671), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g754 ( .A(n_679), .Y(n_754) );
OR2x2_ASAP7_75t_L g770 ( .A(n_679), .B(n_709), .Y(n_770) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B(n_687), .Y(n_681) );
OAI31xp33_ASAP7_75t_L g695 ( .A1(n_682), .A2(n_696), .A3(n_697), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g727 ( .A(n_692), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND4xp25_ASAP7_75t_SL g694 ( .A(n_695), .B(n_703), .C(n_714), .D(n_719), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_702), .Y(n_737) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B1(n_727), .B2(n_729), .C(n_731), .Y(n_719) );
NAND2xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g764 ( .A(n_723), .Y(n_764) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g759 ( .A(n_733), .Y(n_759) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_739), .B(n_758), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_742), .B2(n_744), .C(n_748), .Y(n_739) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_753), .B(n_756), .Y(n_748) );
INVxp33_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_772), .Y(n_785) );
CKINVDCx11_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_776), .B(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_790), .B(n_806), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_795), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g808 ( .A(n_794), .Y(n_808) );
XNOR2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
NAND3x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .C(n_799), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g805 ( .A(n_803), .Y(n_805) );
INVx1_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_SL g817 ( .A(n_810), .Y(n_817) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_SL g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
endmodule