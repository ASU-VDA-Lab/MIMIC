module fake_jpeg_14138_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_27),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_65),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_6),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_5),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_36),
.CON(n_74),
.SN(n_74)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_74),
.A2(n_84),
.B(n_1),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_37),
.B1(n_32),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_83),
.B1(n_90),
.B2(n_114),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_79),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_26),
.B1(n_16),
.B2(n_23),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_31),
.CON(n_84),
.SN(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_86),
.B1(n_105),
.B2(n_107),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_31),
.B1(n_24),
.B2(n_38),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_21),
.B1(n_35),
.B2(n_49),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_18),
.C(n_22),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_41),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_28),
.B1(n_39),
.B2(n_22),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_42),
.A2(n_21),
.B1(n_35),
.B2(n_2),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_49),
.B(n_35),
.C(n_4),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_21),
.B1(n_9),
.B2(n_12),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_43),
.B(n_8),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_8),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_3),
.B(n_4),
.C(n_35),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_132),
.Y(n_163)
);

BUFx2_ASAP7_75t_SL g119 ( 
.A(n_104),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_86),
.B1(n_116),
.B2(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_133),
.B(n_134),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_0),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_142),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_11),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_76),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_80),
.B1(n_95),
.B2(n_84),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_9),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_156),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_47),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_125),
.C(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_155),
.Y(n_186)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_55),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_170),
.B1(n_125),
.B2(n_120),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_74),
.B1(n_89),
.B2(n_107),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_85),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_179),
.C(n_182),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_175),
.B1(n_181),
.B2(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_89),
.B1(n_72),
.B2(n_99),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_100),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_55),
.B1(n_59),
.B2(n_99),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_72),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_71),
.B(n_59),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_184),
.B(n_191),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_138),
.B(n_137),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_122),
.B(n_147),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_145),
.C(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_163),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_139),
.B(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_151),
.A2(n_155),
.B1(n_126),
.B2(n_121),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_195),
.B1(n_164),
.B2(n_185),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_161),
.B(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_141),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_200),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_207),
.C(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_208),
.B1(n_165),
.B2(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_158),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_150),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_135),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_170),
.A2(n_128),
.B1(n_157),
.B2(n_184),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_213),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_171),
.A3(n_191),
.B1(n_188),
.B2(n_172),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_173),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_220),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_183),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_187),
.C(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_214),
.C(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_164),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_229),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_208),
.B1(n_210),
.B2(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_165),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_256),
.C(n_216),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_238),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_197),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_204),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_213),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_230),
.B(n_233),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_214),
.A2(n_206),
.B1(n_205),
.B2(n_221),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_215),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_238),
.B1(n_235),
.B2(n_240),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_259),
.C(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_218),
.B(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_270),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_251),
.A3(n_239),
.B1(n_253),
.B2(n_236),
.C1(n_255),
.C2(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_263),
.B(n_269),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_273),
.B1(n_244),
.B2(n_272),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_254),
.C(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_277),
.C(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_246),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_242),
.B(n_234),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_274),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_237),
.B(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_242),
.C(n_247),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_283),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_249),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_244),
.B1(n_272),
.B2(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_283),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_266),
.C(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

AOI221xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_268),
.B1(n_264),
.B2(n_260),
.C(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_292),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_271),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_273),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_265),
.B1(n_274),
.B2(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_302),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_289),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_279),
.B(n_280),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_305),
.B(n_298),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_286),
.B1(n_299),
.B2(n_303),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_313),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_296),
.C(n_305),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_316),
.Y(n_323)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_294),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_294),
.C(n_302),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_321),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_312),
.B(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_315),
.C(n_307),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_327),
.B(n_319),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_310),
.Y(n_327)
);

OAI211xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_323),
.B(n_320),
.C(n_318),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_325),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_331),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_324),
.Y(n_336)
);


endmodule