module fake_jpeg_10775_n_584 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_584);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_64),
.Y(n_134)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_68),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_9),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_72),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_80),
.B(n_83),
.Y(n_143)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_18),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_86),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_89),
.Y(n_175)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_105),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_17),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_16),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_112),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_28),
.B(n_13),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_31),
.B(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_117),
.Y(n_176)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_11),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_124),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_26),
.B(n_0),
.CON(n_121),
.SN(n_121)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_54),
.Y(n_146)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_32),
.B(n_10),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_131),
.B(n_132),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_135),
.B(n_164),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_151),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_146),
.B(n_22),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_69),
.B(n_44),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_157),
.B(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_55),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_174),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_74),
.B(n_55),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_68),
.B(n_57),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_106),
.B(n_51),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_178),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_65),
.A2(n_56),
.B1(n_57),
.B2(n_53),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_196),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

BUFx16f_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_96),
.B(n_20),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_190),
.B(n_193),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_20),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_108),
.A2(n_53),
.B1(n_57),
.B2(n_42),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_197),
.A2(n_202),
.B1(n_193),
.B2(n_127),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_86),
.B(n_20),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_200),
.B(n_210),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_100),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_201),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_90),
.B(n_42),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_54),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_113),
.B(n_10),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_22),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_42),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_212),
.B(n_250),
.Y(n_287)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_214),
.Y(n_309)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_215),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_134),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_218),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_67),
.B1(n_75),
.B2(n_73),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_217),
.A2(n_277),
.B1(n_196),
.B2(n_200),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_134),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_220),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_138),
.Y(n_222)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_223),
.A2(n_201),
.B(n_204),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_138),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_224),
.B(n_242),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_146),
.A2(n_125),
.B1(n_42),
.B2(n_7),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_227),
.A2(n_269),
.B1(n_188),
.B2(n_208),
.Y(n_308)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_229),
.A2(n_227),
.B1(n_239),
.B2(n_269),
.Y(n_323)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_141),
.B(n_5),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_234),
.B(n_236),
.Y(n_300)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_141),
.B(n_5),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_237),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_6),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_205),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_240),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_152),
.Y(n_241)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_182),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_8),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_137),
.Y(n_247)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_173),
.B(n_8),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_178),
.B(n_176),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_254),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_190),
.Y(n_254)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_155),
.Y(n_258)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_130),
.Y(n_259)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_173),
.B(n_143),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_261),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_143),
.B(n_189),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_266),
.Y(n_334)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_271),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_195),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_267),
.B(n_270),
.Y(n_335)
);

CKINVDCx12_ASAP7_75t_R g268 ( 
.A(n_195),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_268),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_203),
.A2(n_158),
.B1(n_175),
.B2(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_176),
.B(n_172),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_275),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_210),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_274),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_199),
.B(n_206),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_167),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_280),
.A2(n_281),
.B1(n_162),
.B2(n_150),
.Y(n_315)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_198),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_204),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_298),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_290),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_223),
.A2(n_192),
.B(n_180),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_294),
.A2(n_299),
.B(n_251),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_217),
.A2(n_158),
.B1(n_133),
.B2(n_148),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_297),
.A2(n_256),
.B1(n_258),
.B2(n_283),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_163),
.B(n_147),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_229),
.A2(n_136),
.B1(n_154),
.B2(n_128),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_302),
.A2(n_321),
.B1(n_323),
.B2(n_294),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_128),
.B1(n_133),
.B2(n_148),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_305),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_159),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_322),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_232),
.A2(n_150),
.B1(n_181),
.B2(n_156),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_319),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g321 ( 
.A1(n_240),
.A2(n_181),
.B1(n_156),
.B2(n_162),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_212),
.B(n_221),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_225),
.B(n_246),
.CI(n_253),
.CON(n_325),
.SN(n_325)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_325),
.B(n_271),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_212),
.B(n_231),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_230),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_253),
.B(n_235),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_283),
.C(n_222),
.Y(n_343)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_340),
.A2(n_296),
.B1(n_320),
.B2(n_327),
.Y(n_385)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_337),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_331),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_370),
.Y(n_386)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_226),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_346),
.B(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_271),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_352),
.B(n_366),
.Y(n_399)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_354),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_213),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_367),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_360),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_321),
.B1(n_337),
.B2(n_297),
.Y(n_401)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_285),
.B(n_259),
.Y(n_360)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_376),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_245),
.Y(n_370)
);

OAI32xp33_ASAP7_75t_L g371 ( 
.A1(n_316),
.A2(n_215),
.A3(n_265),
.B1(n_255),
.B2(n_237),
.Y(n_371)
);

AOI32xp33_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_290),
.A3(n_308),
.B1(n_323),
.B2(n_286),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_255),
.B(n_233),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_372),
.A2(n_373),
.B(n_299),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_322),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_287),
.C(n_336),
.Y(n_400)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_378),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_287),
.B(n_280),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_324),
.B(n_247),
.Y(n_377)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_326),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_300),
.B(n_334),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_332),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_385),
.A2(n_345),
.B1(n_339),
.B2(n_348),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_365),
.A2(n_380),
.B1(n_358),
.B2(n_351),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_413),
.B1(n_376),
.B2(n_372),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_310),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_363),
.A2(n_357),
.B1(n_380),
.B2(n_365),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_398),
.A2(n_410),
.B(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_350),
.C(n_286),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_401),
.A2(n_402),
.B1(n_375),
.B2(n_361),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_358),
.B1(n_349),
.B2(n_323),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_411),
.B1(n_289),
.B2(n_367),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_343),
.B(n_377),
.Y(n_423)
);

AO22x1_ASAP7_75t_SL g408 ( 
.A1(n_363),
.A2(n_323),
.B1(n_301),
.B2(n_327),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_409),
.Y(n_420)
);

OA22x2_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_295),
.B1(n_328),
.B2(n_303),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_349),
.A2(n_324),
.B1(n_312),
.B2(n_317),
.Y(n_411)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

OAI22x1_ASAP7_75t_SL g413 ( 
.A1(n_371),
.A2(n_312),
.B1(n_317),
.B2(n_332),
.Y(n_413)
);

OA22x2_ASAP7_75t_L g415 ( 
.A1(n_344),
.A2(n_303),
.B1(n_318),
.B2(n_310),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_416),
.A2(n_417),
.B1(n_431),
.B2(n_435),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_387),
.A2(n_369),
.B1(n_359),
.B2(n_362),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_391),
.B(n_356),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_418),
.B(n_426),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_374),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_425),
.C(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_423),
.A2(n_427),
.B(n_395),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_360),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_355),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_428),
.B(n_430),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_386),
.B(n_341),
.Y(n_429)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_335),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_293),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_434),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_412),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_364),
.B1(n_353),
.B2(n_347),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_436),
.A2(n_437),
.B1(n_446),
.B2(n_405),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_396),
.B(n_379),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_445),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_425),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_368),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_307),
.C(n_318),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_439),
.C(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_398),
.A2(n_338),
.B1(n_314),
.B2(n_307),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_438),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_448),
.B(n_450),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_429),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_445),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_451),
.B(n_434),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_416),
.A2(n_401),
.B1(n_408),
.B2(n_406),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_455),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_424),
.A2(n_404),
.B(n_395),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_454),
.A2(n_475),
.B(n_390),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_396),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_461),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_457),
.A2(n_420),
.B1(n_422),
.B2(n_432),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_473),
.C(n_474),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_410),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_471),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_469),
.Y(n_480)
);

INVx3_ASAP7_75t_SL g470 ( 
.A(n_431),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_409),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_408),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_409),
.C(n_414),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_392),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_424),
.A2(n_409),
.B(n_390),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_420),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_476),
.B(n_494),
.Y(n_507)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_479),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_421),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_484),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_460),
.B(n_418),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_486),
.B(n_492),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_487),
.A2(n_453),
.B1(n_472),
.B2(n_471),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_447),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_490),
.Y(n_512)
);

AO22x1_ASAP7_75t_L g490 ( 
.A1(n_475),
.A2(n_427),
.B1(n_443),
.B2(n_441),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_452),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_493),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_414),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_456),
.B(n_444),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_495),
.A2(n_469),
.B1(n_454),
.B2(n_449),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_496),
.B(n_499),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_447),
.B(n_461),
.C(n_455),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_465),
.C(n_449),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_466),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_382),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_501),
.A2(n_503),
.B1(n_490),
.B2(n_484),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_470),
.B1(n_474),
.B2(n_457),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_504),
.A2(n_495),
.B(n_480),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_506),
.B(n_490),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g508 ( 
.A(n_476),
.B(n_463),
.CI(n_415),
.CON(n_508),
.SN(n_508)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_510),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_392),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_494),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_388),
.C(n_382),
.Y(n_510)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_516),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_485),
.B(n_388),
.C(n_381),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_520),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_381),
.C(n_415),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_527),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_488),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_523),
.B(n_526),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_515),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_524),
.A2(n_503),
.B1(n_501),
.B2(n_511),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_518),
.B(n_489),
.Y(n_528)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_528),
.Y(n_542)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_517),
.Y(n_530)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_530),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_481),
.C(n_497),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_533),
.C(n_520),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_502),
.B(n_483),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_507),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_497),
.C(n_491),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_513),
.B(n_478),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_SL g537 ( 
.A(n_534),
.B(n_535),
.Y(n_537)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_514),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_536),
.A2(n_500),
.B1(n_479),
.B2(n_507),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_544),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_539),
.A2(n_541),
.B1(n_543),
.B2(n_532),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_524),
.A2(n_505),
.B1(n_504),
.B2(n_508),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_521),
.A2(n_508),
.B1(n_493),
.B2(n_512),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_509),
.C(n_512),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_546),
.A2(n_525),
.B1(n_531),
.B2(n_529),
.Y(n_552)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_547),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_415),
.C(n_342),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_278),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_522),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_551),
.B(n_553),
.Y(n_562)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_552),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_536),
.C(n_527),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_542),
.A2(n_545),
.B(n_549),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_554),
.A2(n_550),
.B(n_552),
.Y(n_566)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_556),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_546),
.A2(n_532),
.B1(n_314),
.B2(n_257),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_559),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_539),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_560),
.Y(n_568)
);

AOI31xp67_ASAP7_75t_L g563 ( 
.A1(n_557),
.A2(n_537),
.A3(n_541),
.B(n_543),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_354),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_558),
.B(n_544),
.C(n_545),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_565),
.B(n_309),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_566),
.A2(n_547),
.B(n_556),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_562),
.B(n_553),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_569),
.B(n_571),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_570),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_572),
.B(n_573),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_561),
.A2(n_262),
.B1(n_309),
.B2(n_313),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_313),
.C(n_244),
.Y(n_574)
);

AOI21xp33_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_569),
.B(n_568),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_579),
.C(n_575),
.Y(n_580)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_576),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_580),
.A2(n_564),
.B(n_574),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_568),
.B(n_244),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_582),
.B(n_219),
.Y(n_583)
);

AO21x1_ASAP7_75t_L g584 ( 
.A1(n_583),
.A2(n_244),
.B(n_214),
.Y(n_584)
);


endmodule