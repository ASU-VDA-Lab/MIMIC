module fake_netlist_6_1981_n_1070 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_265, n_113, n_39, n_63, n_223, n_270, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1070);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_270;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1070;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_842;
wire n_758;
wire n_611;
wire n_943;
wire n_491;
wire n_843;
wire n_656;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_683;
wire n_811;
wire n_620;
wire n_420;
wire n_878;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_1051;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_474;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_861;
wire n_296;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_672;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_663;
wire n_508;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_10),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_109),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_151),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_215),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_138),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_15),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_156),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_50),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_163),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_46),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_54),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_167),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_65),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_80),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_187),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_145),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_68),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_241),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_195),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_129),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_108),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_98),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_113),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_85),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_192),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_74),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_174),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_176),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_32),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_159),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_168),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_88),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_17),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_124),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_69),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_76),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_153),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_100),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_131),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_170),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_92),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_99),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_169),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_111),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_53),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_49),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_48),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_114),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_173),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_51),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_66),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_207),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_144),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_247),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_72),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_101),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_107),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_193),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_60),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_89),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_161),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_225),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_83),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_197),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_55),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_130),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_235),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_93),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_203),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_148),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_75),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_3),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_141),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_196),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_271),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_265),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_110),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_86),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_94),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_258),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_106),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_7),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_96),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_42),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_27),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_256),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_172),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_4),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_270),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_262),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_127),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_221),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_45),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_233),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_204),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_249),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_189),
.Y(n_392)
);

CKINVDCx6p67_ASAP7_75t_R g393 ( 
.A(n_142),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_37),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_132),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_191),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_213),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_97),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_181),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_44),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_91),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_123),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_120),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_16),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_134),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_95),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_186),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_149),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_232),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_135),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_112),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_18),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_269),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_246),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_56),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_244),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_245),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_121),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_229),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_105),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_23),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_28),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_87),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_2),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_171),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_12),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_71),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_119),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_63),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_243),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_10),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_208),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_90),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_29),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_11),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_137),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_140),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_226),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_240),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_214),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_17),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_212),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_254),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_118),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_188),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_58),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_27),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_185),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_103),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_9),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_282),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_272),
.Y(n_454)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_320),
.B(n_0),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_272),
.Y(n_457)
);

BUFx8_ASAP7_75t_SL g458 ( 
.A(n_291),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_320),
.B(n_385),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_272),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_411),
.B(n_0),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_273),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_295),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_273),
.B(n_1),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_1),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_272),
.B(n_40),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_2),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_294),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_294),
.B(n_3),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_315),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

BUFx8_ASAP7_75t_SL g475 ( 
.A(n_291),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_390),
.B(n_5),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_335),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_335),
.B(n_6),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_334),
.B(n_6),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_343),
.B(n_7),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_354),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_354),
.B(n_367),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

BUFx8_ASAP7_75t_SL g487 ( 
.A(n_422),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_442),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_425),
.B(n_296),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_349),
.B(n_8),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_296),
.B(n_8),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_425),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_448),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_274),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_280),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_284),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_311),
.B(n_344),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_311),
.B(n_43),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_380),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_11),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_405),
.B(n_12),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_344),
.B(n_13),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_352),
.Y(n_504)
);

INVx6_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_275),
.Y(n_506)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_352),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_430),
.B(n_14),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_310),
.B(n_14),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_15),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_287),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_421),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_290),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_276),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_298),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_439),
.B(n_16),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_314),
.B(n_18),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_304),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_305),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_306),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_308),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_313),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_321),
.B(n_19),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_325),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_332),
.B(n_19),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_277),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_278),
.Y(n_533)
);

BUFx12f_ASAP7_75t_L g534 ( 
.A(n_279),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_361),
.B(n_20),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_281),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_362),
.B(n_20),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_364),
.B(n_21),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_365),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_366),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_368),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_382),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_388),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_326),
.B(n_21),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_398),
.B(n_400),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_283),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_285),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_286),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_415),
.B(n_22),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_461),
.A2(n_408),
.B1(n_437),
.B2(n_396),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_464),
.A2(n_416),
.B1(n_419),
.B2(n_417),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_459),
.B(n_414),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_464),
.A2(n_423),
.B1(n_428),
.B2(n_420),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_505),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_456),
.B(n_408),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_469),
.A2(n_479),
.B1(n_465),
.B2(n_467),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_470),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_477),
.A2(n_438),
.B1(n_437),
.B2(n_330),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_469),
.A2(n_434),
.B1(n_440),
.B2(n_433),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_452),
.A2(n_438),
.B1(n_331),
.B2(n_355),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_R g566 ( 
.A1(n_541),
.A2(n_481),
.B1(n_514),
.B2(n_494),
.Y(n_566)
);

AO22x1_ASAP7_75t_SL g567 ( 
.A1(n_512),
.A2(n_449),
.B1(n_450),
.B2(n_447),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_519),
.A2(n_455),
.B1(n_490),
.B2(n_480),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_502),
.A2(n_545),
.B1(n_501),
.B2(n_482),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_455),
.A2(n_503),
.B1(n_509),
.B2(n_491),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

NAND3x1_ASAP7_75t_L g573 ( 
.A(n_511),
.B(n_22),
.C(n_23),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_505),
.A2(n_289),
.B1(n_292),
.B2(n_288),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_500),
.B(n_303),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_R g577 ( 
.A1(n_458),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_518),
.A2(n_372),
.B1(n_446),
.B2(n_359),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_538),
.A2(n_549),
.B1(n_535),
.B2(n_531),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_552),
.A2(n_297),
.B1(n_299),
.B2(n_293),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_546),
.A2(n_445),
.B1(n_444),
.B2(n_443),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_492),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_507),
.A2(n_353),
.B1(n_431),
.B2(n_426),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_506),
.B(n_300),
.Y(n_584)
);

INVx6_ASAP7_75t_L g585 ( 
.A(n_521),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_479),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_516),
.A2(n_496),
.B1(n_550),
.B2(n_534),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_512),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_549),
.A2(n_441),
.B1(n_418),
.B2(n_413),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_527),
.A2(n_410),
.B1(n_407),
.B2(n_406),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_492),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_527),
.A2(n_347),
.B1(n_401),
.B2(n_399),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_486),
.B(n_301),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_538),
.A2(n_402),
.B1(n_397),
.B2(n_395),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_462),
.A2(n_392),
.B1(n_391),
.B2(n_389),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_497),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_468),
.A2(n_387),
.B1(n_386),
.B2(n_384),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_471),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_302),
.Y(n_601)
);

INVx8_ASAP7_75t_L g602 ( 
.A(n_532),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_537),
.A2(n_539),
.B1(n_506),
.B2(n_485),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_485),
.B(n_307),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_521),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_486),
.B(n_309),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_453),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_540),
.Y(n_608)
);

OA22x2_ASAP7_75t_L g609 ( 
.A1(n_463),
.A2(n_381),
.B1(n_379),
.B2(n_378),
.Y(n_609)
);

AO22x2_ASAP7_75t_L g610 ( 
.A1(n_537),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_539),
.A2(n_339),
.B1(n_375),
.B2(n_374),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_489),
.B(n_312),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_493),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_489),
.A2(n_376),
.B1(n_373),
.B2(n_371),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_543),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_R g616 ( 
.A1(n_475),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_498),
.A2(n_370),
.B1(n_369),
.B2(n_363),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_495),
.A2(n_360),
.B1(n_358),
.B2(n_357),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_498),
.A2(n_333),
.B1(n_351),
.B2(n_350),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_495),
.B(n_316),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_495),
.B(n_317),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_472),
.A2(n_356),
.B1(n_348),
.B2(n_346),
.Y(n_622)
);

OA22x2_ASAP7_75t_L g623 ( 
.A1(n_476),
.A2(n_488),
.B1(n_483),
.B2(n_551),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_486),
.B(n_345),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_544),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_513),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_521),
.B(n_523),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_515),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_466),
.A2(n_342),
.B1(n_341),
.B2(n_340),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_466),
.A2(n_327),
.B1(n_337),
.B2(n_336),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_626),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_596),
.B(n_532),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_628),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_607),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_601),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_561),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_553),
.B(n_587),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_579),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_562),
.Y(n_641)
);

INVxp33_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_600),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_604),
.B(n_523),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_582),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_591),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_620),
.B(n_523),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_559),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_613),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_574),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_631),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_597),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_583),
.B(n_532),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_608),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_571),
.B(n_533),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_615),
.Y(n_660)
);

OR2x2_ASAP7_75t_SL g661 ( 
.A(n_566),
.B(n_487),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_625),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_621),
.B(n_528),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_563),
.B(n_466),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_560),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_560),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_622),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_603),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_554),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_609),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_557),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_557),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_564),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_564),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_569),
.B(n_499),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_573),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_558),
.B(n_528),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_629),
.B(n_520),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

XOR2x2_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_33),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_606),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_624),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_627),
.A2(n_522),
.B(n_457),
.Y(n_685)
);

XOR2xp5_ASAP7_75t_L g686 ( 
.A(n_565),
.B(n_318),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_605),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_584),
.B(n_528),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_585),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_588),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_619),
.B(n_529),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_585),
.B(n_529),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_588),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_586),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_610),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_590),
.B(n_529),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_592),
.B(n_533),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_630),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_581),
.B(n_533),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_SL g702 ( 
.A(n_578),
.B(n_319),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_602),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_576),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_595),
.B(n_599),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_611),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_614),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_594),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_580),
.A2(n_457),
.B(n_454),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_576),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_589),
.B(n_536),
.Y(n_711)
);

INVxp33_ASAP7_75t_L g712 ( 
.A(n_617),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_602),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_575),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_642),
.B(n_524),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_636),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_642),
.B(n_524),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_654),
.B(n_670),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_636),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_666),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_666),
.B(n_525),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_669),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_680),
.B(n_536),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_632),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_665),
.B(n_47),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_682),
.B(n_536),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_651),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_678),
.Y(n_730)
);

AND2x6_ASAP7_75t_SL g731 ( 
.A(n_705),
.B(n_577),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_651),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_672),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_707),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_683),
.B(n_525),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_643),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_676),
.B(n_649),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_676),
.B(n_454),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_659),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_640),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_663),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_637),
.B(n_525),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_653),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_708),
.B(n_618),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_700),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_688),
.B(n_547),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_658),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_644),
.B(n_547),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_669),
.B(n_34),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_660),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_673),
.B(n_526),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_673),
.B(n_526),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_679),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_679),
.B(n_526),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_690),
.B(n_693),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_662),
.Y(n_758)
);

AND2x2_ASAP7_75t_SL g759 ( 
.A(n_664),
.B(n_616),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_705),
.B(n_547),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_635),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_706),
.B(n_548),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_684),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_638),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_633),
.B(n_548),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_641),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_703),
.B(n_548),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_677),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_633),
.B(n_530),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_701),
.B(n_322),
.Y(n_770)
);

AND2x2_ASAP7_75t_SL g771 ( 
.A(n_650),
.B(n_530),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_645),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_671),
.B(n_530),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_646),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_647),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_685),
.Y(n_776)
);

OR2x2_ASAP7_75t_SL g777 ( 
.A(n_694),
.B(n_542),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_648),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_711),
.B(n_542),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_652),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_699),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_702),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_674),
.B(n_542),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_708),
.A2(n_338),
.B(n_324),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_675),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_695),
.B(n_696),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_697),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_698),
.B(n_504),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_699),
.B(n_52),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_712),
.A2(n_691),
.B(n_709),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_755),
.B(n_689),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_721),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_768),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_721),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_721),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_721),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_738),
.B(n_677),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_687),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_721),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_740),
.B(n_714),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_719),
.B(n_656),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_755),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_715),
.B(n_667),
.Y(n_803)
);

AND2x6_ASAP7_75t_L g804 ( 
.A(n_726),
.B(n_703),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_789),
.B(n_710),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_719),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_725),
.B(n_713),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_768),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_732),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_740),
.B(n_717),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_732),
.Y(n_811)
);

BUFx12f_ASAP7_75t_L g812 ( 
.A(n_731),
.Y(n_812)
);

INVx6_ASAP7_75t_L g813 ( 
.A(n_781),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_716),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_743),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_725),
.B(n_713),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_759),
.B(n_681),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_740),
.B(n_714),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_787),
.B(n_686),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_755),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_789),
.B(n_692),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_737),
.B(n_640),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_755),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_755),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_763),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_737),
.B(n_704),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_718),
.B(n_667),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_782),
.B(n_661),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_757),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_789),
.B(n_681),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_726),
.B(n_454),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_744),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_740),
.B(n_702),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_723),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_744),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_759),
.B(n_639),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_740),
.B(n_323),
.Y(n_837)
);

AO21x2_ASAP7_75t_L g838 ( 
.A1(n_760),
.A2(n_329),
.B(n_328),
.Y(n_838)
);

CKINVDCx8_ASAP7_75t_R g839 ( 
.A(n_726),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_742),
.B(n_704),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_802),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_809),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_808),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_803),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_820),
.B(n_778),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_827),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_820),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_806),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_811),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_829),
.Y(n_850)
);

INVx3_ASAP7_75t_SL g851 ( 
.A(n_822),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_824),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_795),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_820),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_800),
.A2(n_746),
.B1(n_734),
.B2(n_747),
.Y(n_855)
);

BUFx2_ASAP7_75t_SL g856 ( 
.A(n_823),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_797),
.B(n_735),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_802),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_823),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_826),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_832),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_826),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_797),
.B(n_735),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_829),
.B(n_753),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_792),
.Y(n_865)
);

BUFx2_ASAP7_75t_SL g866 ( 
.A(n_823),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_834),
.Y(n_867)
);

BUFx12f_ASAP7_75t_L g868 ( 
.A(n_812),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_824),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_793),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_825),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_840),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_800),
.B(n_720),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_870),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_844),
.A2(n_817),
.B1(n_819),
.B2(n_836),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_844),
.A2(n_784),
.B1(n_790),
.B2(n_818),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_854),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_849),
.Y(n_878)
);

OAI22xp33_ASAP7_75t_L g879 ( 
.A1(n_855),
.A2(n_830),
.B1(n_818),
.B2(n_839),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_842),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_857),
.B(n_863),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_846),
.A2(n_830),
.B1(n_822),
.B2(n_828),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_855),
.B(n_815),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_846),
.A2(n_814),
.B1(n_801),
.B2(n_733),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_871),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

INVx11_ASAP7_75t_L g887 ( 
.A(n_872),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_873),
.A2(n_830),
.B1(n_771),
.B2(n_801),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_864),
.A2(n_781),
.B1(n_798),
.B2(n_833),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_851),
.Y(n_890)
);

INVx6_ASAP7_75t_L g891 ( 
.A(n_854),
.Y(n_891)
);

CKINVDCx6p67_ASAP7_75t_R g892 ( 
.A(n_851),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_843),
.Y(n_893)
);

BUFx12f_ASAP7_75t_L g894 ( 
.A(n_860),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_867),
.A2(n_833),
.B1(n_810),
.B2(n_814),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_851),
.A2(n_756),
.B1(n_804),
.B2(n_770),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_850),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_848),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_872),
.A2(n_741),
.B1(n_840),
.B2(n_816),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_875),
.A2(n_848),
.B1(n_777),
.B2(n_850),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_878),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_881),
.B(n_743),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_894),
.A2(n_741),
.B1(n_862),
.B2(n_860),
.Y(n_903)
);

OAI222xp33_ASAP7_75t_L g904 ( 
.A1(n_879),
.A2(n_810),
.B1(n_779),
.B2(n_739),
.C1(n_770),
.C2(n_867),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_879),
.A2(n_862),
.B1(n_807),
.B2(n_816),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_888),
.A2(n_756),
.B1(n_744),
.B2(n_838),
.Y(n_906)
);

OAI222xp33_ASAP7_75t_L g907 ( 
.A1(n_882),
.A2(n_739),
.B1(n_805),
.B2(n_837),
.C1(n_751),
.C2(n_849),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_876),
.A2(n_744),
.B1(n_838),
.B2(n_804),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_899),
.A2(n_807),
.B1(n_742),
.B2(n_730),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_897),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_893),
.B(n_773),
.Y(n_911)
);

CKINVDCx8_ASAP7_75t_R g912 ( 
.A(n_886),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_884),
.A2(n_742),
.B1(n_821),
.B2(n_805),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_883),
.B(n_753),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_897),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_889),
.A2(n_831),
.B1(n_852),
.B2(n_869),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_880),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_896),
.A2(n_804),
.B1(n_749),
.B2(n_758),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_895),
.A2(n_804),
.B1(n_749),
.B2(n_758),
.Y(n_919)
);

INVx5_ASAP7_75t_L g920 ( 
.A(n_877),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_885),
.A2(n_837),
.B1(n_727),
.B2(n_736),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_893),
.A2(n_852),
.B1(n_805),
.B2(n_813),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_890),
.A2(n_866),
.B1(n_856),
.B2(n_813),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_SL g924 ( 
.A1(n_874),
.A2(n_762),
.B(n_752),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_874),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_877),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_892),
.A2(n_736),
.B1(n_780),
.B2(n_778),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_898),
.A2(n_778),
.B1(n_766),
.B2(n_775),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_898),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_877),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_902),
.A2(n_772),
.B1(n_761),
.B2(n_764),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_914),
.A2(n_900),
.B1(n_921),
.B2(n_911),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_925),
.B(n_865),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_924),
.B(n_865),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_910),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_906),
.A2(n_772),
.B1(n_764),
.B2(n_761),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_926),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_905),
.A2(n_821),
.B1(n_767),
.B2(n_728),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_909),
.A2(n_887),
.B1(n_821),
.B2(n_751),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_913),
.A2(n_724),
.B1(n_750),
.B2(n_748),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_903),
.A2(n_774),
.B1(n_745),
.B2(n_832),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_916),
.A2(n_774),
.B1(n_745),
.B2(n_835),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_908),
.A2(n_745),
.B1(n_835),
.B2(n_729),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_918),
.A2(n_927),
.B1(n_928),
.B2(n_923),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_922),
.B(n_765),
.C(n_769),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_917),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_919),
.A2(n_783),
.B1(n_861),
.B2(n_868),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_915),
.B(n_853),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_901),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_929),
.A2(n_722),
.B1(n_754),
.B2(n_785),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_929),
.A2(n_722),
.B1(n_785),
.B2(n_794),
.Y(n_951)
);

OA21x2_ASAP7_75t_L g952 ( 
.A1(n_904),
.A2(n_907),
.B(n_799),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_930),
.A2(n_861),
.B1(n_791),
.B2(n_796),
.Y(n_953)
);

AOI222xp33_ASAP7_75t_L g954 ( 
.A1(n_929),
.A2(n_757),
.B1(n_786),
.B2(n_788),
.C1(n_723),
.C2(n_504),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_912),
.B(n_891),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_920),
.A2(n_841),
.B1(n_858),
.B2(n_866),
.Y(n_956)
);

AOI222xp33_ASAP7_75t_L g957 ( 
.A1(n_920),
.A2(n_786),
.B1(n_788),
.B2(n_508),
.C1(n_510),
.C2(n_38),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_911),
.B(n_841),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_925),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_902),
.B(n_858),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_905),
.A2(n_845),
.B1(n_858),
.B2(n_856),
.Y(n_961)
);

NAND4xp25_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_932),
.C(n_954),
.D(n_934),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_932),
.A2(n_510),
.B1(n_508),
.B2(n_37),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_939),
.A2(n_510),
.B1(n_508),
.B2(n_859),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_59),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_946),
.B(n_62),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_SL g967 ( 
.A1(n_938),
.A2(n_859),
.B(n_854),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_935),
.B(n_64),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_937),
.B(n_67),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_949),
.B(n_73),
.Y(n_970)
);

OAI22xp33_ASAP7_75t_L g971 ( 
.A1(n_952),
.A2(n_859),
.B1(n_854),
.B2(n_847),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_958),
.B(n_78),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_960),
.B(n_79),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_961),
.B(n_81),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_955),
.B(n_82),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_933),
.B(n_948),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_940),
.B(n_84),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_941),
.A2(n_859),
.B1(n_854),
.B2(n_776),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_931),
.B(n_102),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_950),
.B(n_859),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_931),
.B(n_952),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_952),
.B(n_104),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_944),
.B(n_947),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_956),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_953),
.B(n_942),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_L g986 ( 
.A(n_962),
.B(n_945),
.C(n_936),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_943),
.Y(n_987)
);

NAND4xp75_ASAP7_75t_L g988 ( 
.A(n_977),
.B(n_115),
.C(n_116),
.D(n_117),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_951),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_951),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_950),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_969),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_975),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_971),
.B(n_457),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_972),
.B(n_122),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_L g996 ( 
.A(n_963),
.B(n_776),
.C(n_474),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_973),
.B(n_125),
.C(n_126),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_963),
.B(n_974),
.Y(n_998)
);

AO21x2_ASAP7_75t_L g999 ( 
.A1(n_971),
.A2(n_128),
.B(n_133),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_974),
.B(n_776),
.C(n_474),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_965),
.B(n_136),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_983),
.A2(n_776),
.B1(n_474),
.B2(n_473),
.Y(n_1002)
);

OA211x2_ASAP7_75t_L g1003 ( 
.A1(n_964),
.A2(n_139),
.B(n_143),
.C(n_146),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_967),
.B(n_776),
.C(n_473),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_989),
.B(n_970),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_998),
.B(n_993),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_986),
.B(n_964),
.C(n_980),
.Y(n_1007)
);

NAND4xp75_ASAP7_75t_L g1008 ( 
.A(n_998),
.B(n_968),
.C(n_966),
.D(n_985),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_992),
.B(n_978),
.Y(n_1009)
);

XNOR2xp5_ASAP7_75t_L g1010 ( 
.A(n_991),
.B(n_979),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_999),
.Y(n_1011)
);

NAND4xp75_ASAP7_75t_SL g1012 ( 
.A(n_990),
.B(n_147),
.C(n_150),
.D(n_152),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_999),
.Y(n_1013)
);

NAND4xp75_ASAP7_75t_SL g1014 ( 
.A(n_990),
.B(n_157),
.C(n_158),
.D(n_160),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_989),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_994),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_988),
.A2(n_473),
.B1(n_460),
.B2(n_165),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_987),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_SL g1019 ( 
.A1(n_1000),
.A2(n_460),
.B1(n_164),
.B2(n_166),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1001),
.B(n_994),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1015),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1006),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_1011),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_1009),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1005),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1016),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1011),
.B(n_995),
.Y(n_1028)
);

XOR2x2_ASAP7_75t_L g1029 ( 
.A(n_1008),
.B(n_996),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1030)
);

XOR2x2_ASAP7_75t_L g1031 ( 
.A(n_1010),
.B(n_997),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1020),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1016),
.Y(n_1033)
);

XOR2xp5_ASAP7_75t_L g1034 ( 
.A(n_1007),
.B(n_1003),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1013),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1024),
.Y(n_1036)
);

AO22x2_ASAP7_75t_L g1037 ( 
.A1(n_1035),
.A2(n_1007),
.B1(n_1014),
.B2(n_1012),
.Y(n_1037)
);

OA22x2_ASAP7_75t_L g1038 ( 
.A1(n_1034),
.A2(n_1017),
.B1(n_1019),
.B2(n_177),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1027),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1029),
.A2(n_162),
.B1(n_179),
.B2(n_180),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1022),
.A2(n_1025),
.B1(n_1030),
.B2(n_1023),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1033),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1021),
.Y(n_1043)
);

AOI22x1_ASAP7_75t_SL g1044 ( 
.A1(n_1022),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_1044)
);

OA22x2_ASAP7_75t_L g1045 ( 
.A1(n_1028),
.A2(n_190),
.B1(n_194),
.B2(n_199),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1031),
.A2(n_201),
.B1(n_202),
.B2(n_205),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1030),
.A2(n_1023),
.B1(n_1032),
.B2(n_1026),
.Y(n_1047)
);

OAI322xp33_ASAP7_75t_L g1048 ( 
.A1(n_1041),
.A2(n_206),
.A3(n_209),
.B1(n_210),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1036),
.Y(n_1049)
);

OAI322xp33_ASAP7_75t_L g1050 ( 
.A1(n_1047),
.A2(n_220),
.A3(n_222),
.B1(n_223),
.B2(n_224),
.C1(n_227),
.C2(n_228),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1049),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1048),
.A2(n_1038),
.B1(n_1037),
.B2(n_1040),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1050),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1051),
.Y(n_1054)
);

AND4x1_ASAP7_75t_L g1055 ( 
.A(n_1052),
.B(n_1046),
.C(n_1044),
.D(n_1042),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_1053),
.B(n_1039),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1055),
.A2(n_1045),
.B(n_1043),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_1037),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1058),
.B(n_231),
.Y(n_1060)
);

AO22x2_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_1057),
.B1(n_1059),
.B2(n_236),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_1061),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1062),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1063),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1064),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1065),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1066),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1067),
.Y(n_1068)
);

AOI221xp5_ASAP7_75t_L g1069 ( 
.A1(n_1068),
.A2(n_255),
.B1(n_259),
.B2(n_260),
.C(n_261),
.Y(n_1069)
);

AOI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1069),
.A2(n_266),
.B(n_267),
.C(n_268),
.Y(n_1070)
);


endmodule