module fake_ariane_2450_n_1667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1667;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_85),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_62),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_10),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_28),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_57),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_100),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_21),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_2),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_122),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_22),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_94),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_10),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_136),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_59),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_127),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_51),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_52),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_20),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_21),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_45),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_4),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_69),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_95),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_70),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_88),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_93),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_2),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_32),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_101),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_76),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_75),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_24),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_67),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_0),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_7),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_152),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_51),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_24),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_22),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_20),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_26),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_44),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_46),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_129),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_80),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_41),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_144),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_12),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_115),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_7),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_40),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_4),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_131),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_130),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_123),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_56),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_126),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_48),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_31),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_146),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_78),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_68),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_72),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_97),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_58),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_35),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_151),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_5),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_140),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_41),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_138),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_112),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_31),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_23),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_13),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_55),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_15),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_86),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_143),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_102),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_61),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_60),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_36),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_156),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_176),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_185),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_159),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_160),
.B(n_1),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_165),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_194),
.B(n_3),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_175),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_165),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_193),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_190),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_R g324 ( 
.A(n_238),
.B(n_108),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_172),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_172),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_260),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_234),
.B(n_9),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_295),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_174),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_189),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_215),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_203),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_211),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_215),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_223),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_191),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_196),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_197),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_224),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_198),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_305),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_228),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_222),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_206),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_234),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_202),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_231),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_235),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_208),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_232),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_255),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_253),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_256),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_275),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_214),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_226),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_246),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_222),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_290),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_227),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_246),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_316),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_249),
.C(n_239),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_171),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_313),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_326),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_325),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_351),
.B(n_154),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_219),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_308),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_312),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_312),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_327),
.B(n_241),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

CKINVDCx8_ASAP7_75t_R g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_372),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_336),
.B(n_164),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_337),
.B(n_241),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_335),
.B(n_171),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_340),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_314),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_344),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_346),
.B(n_186),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_350),
.B(n_186),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_350),
.A2(n_183),
.B(n_167),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_362),
.B(n_273),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_373),
.B(n_269),
.Y(n_438)
);

CKINVDCx8_ASAP7_75t_R g439 ( 
.A(n_328),
.Y(n_439)
);

AND3x2_ASAP7_75t_L g440 ( 
.A(n_338),
.B(n_261),
.C(n_291),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_324),
.B(n_157),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_357),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_348),
.B1(n_347),
.B2(n_359),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_415),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_345),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_395),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_381),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_395),
.A2(n_329),
.B1(n_375),
.B2(n_342),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_354),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_385),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

AND2x2_ASAP7_75t_SL g464 ( 
.A(n_438),
.B(n_187),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_403),
.B(n_356),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_383),
.A2(n_349),
.B1(n_366),
.B2(n_310),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_385),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_407),
.B(n_367),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_438),
.B(n_188),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_368),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_403),
.B(n_369),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_393),
.B(n_419),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_407),
.B(n_370),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_413),
.B(n_439),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_376),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_413),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_273),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_383),
.A2(n_309),
.B1(n_371),
.B2(n_178),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_403),
.B(n_331),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_403),
.B(n_332),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_425),
.B(n_153),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_158),
.C(n_157),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_408),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_392),
.B(n_371),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_158),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_169),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_388),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_386),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_388),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_392),
.B(n_200),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_417),
.B(n_169),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_425),
.B(n_153),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_392),
.B(n_201),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_393),
.B(n_210),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_389),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_388),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_425),
.B(n_323),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_425),
.B(n_199),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_426),
.A2(n_210),
.B1(n_243),
.B2(n_251),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_389),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_426),
.A2(n_237),
.B1(n_270),
.B2(n_268),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_425),
.B(n_204),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_389),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_419),
.A2(n_254),
.B1(n_236),
.B2(n_247),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_441),
.B(n_155),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_389),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_415),
.B(n_209),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_391),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_426),
.A2(n_427),
.B1(n_428),
.B2(n_384),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_387),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_391),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_391),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_419),
.A2(n_266),
.B1(n_263),
.B2(n_250),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_387),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_170),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_381),
.A2(n_374),
.B1(n_364),
.B2(n_361),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_411),
.B(n_155),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_419),
.A2(n_181),
.B1(n_305),
.B2(n_303),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_419),
.A2(n_170),
.B1(n_303),
.B2(n_272),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_426),
.B(n_161),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_434),
.B(n_181),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_427),
.B(n_300),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_427),
.B(n_161),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_437),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_416),
.B(n_272),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_391),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_427),
.B(n_162),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_419),
.B(n_233),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_428),
.B(n_387),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_437),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_427),
.A2(n_293),
.B1(n_284),
.B2(n_279),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_420),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_420),
.B(n_343),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_391),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_409),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_384),
.B(n_162),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_300),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_409),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_393),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_384),
.B(n_163),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_391),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_414),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_393),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_428),
.A2(n_293),
.B1(n_284),
.B2(n_279),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_384),
.B(n_163),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_391),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_437),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_440),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_434),
.B(n_154),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_410),
.B(n_422),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_404),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_416),
.B(n_244),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_404),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_484),
.B(n_410),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_484),
.B(n_410),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_SL g591 ( 
.A(n_450),
.B(n_422),
.Y(n_591)
);

BUFx6f_ASAP7_75t_SL g592 ( 
.A(n_464),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_457),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_484),
.B(n_422),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_531),
.B(n_422),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_466),
.B(n_423),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_471),
.B(n_423),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_494),
.B(n_423),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_423),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_514),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_429),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_429),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_460),
.B(n_430),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_577),
.B(n_430),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_559),
.A2(n_586),
.B1(n_548),
.B2(n_474),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_496),
.B(n_432),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_464),
.A2(n_428),
.B1(n_412),
.B2(n_418),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_494),
.B(n_413),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_494),
.B(n_501),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_461),
.B(n_432),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_442),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_444),
.B(n_442),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_564),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_501),
.B(n_439),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_SL g620 ( 
.A(n_461),
.B(n_439),
.C(n_294),
.Y(n_620)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_513),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_455),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_447),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_493),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_586),
.B(n_412),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_412),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_474),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g629 ( 
.A1(n_520),
.A2(n_298),
.B1(n_294),
.B2(n_296),
.C(n_433),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_455),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_495),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_470),
.B(n_412),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_513),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_418),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_546),
.B(n_418),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_469),
.B(n_477),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_474),
.A2(n_436),
.B1(n_435),
.B2(n_433),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_453),
.B(n_569),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_501),
.B(n_418),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_545),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_547),
.A2(n_433),
.B(n_435),
.C(n_431),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_352),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_576),
.Y(n_643)
);

BUFx8_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_498),
.B(n_360),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_453),
.B(n_431),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_565),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_454),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_474),
.A2(n_436),
.B1(n_435),
.B2(n_433),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_542),
.B(n_431),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_542),
.B(n_436),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_498),
.B(n_440),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_SL g653 ( 
.A(n_468),
.B(n_298),
.C(n_296),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_483),
.B(n_166),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_480),
.B(n_378),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_445),
.B(n_448),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_443),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_533),
.B(n_378),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_473),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_459),
.B(n_168),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_445),
.B(n_404),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_526),
.A2(n_382),
.B1(n_394),
.B2(n_380),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_483),
.B(n_380),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_445),
.B(n_404),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_448),
.B(n_404),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_473),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_459),
.B(n_173),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_528),
.B(n_382),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_443),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_508),
.B(n_394),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_446),
.B(n_398),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_567),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_499),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_468),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_448),
.B(n_404),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_508),
.B(n_396),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_518),
.B(n_428),
.C(n_396),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_500),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_446),
.B(n_398),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_541),
.B(n_428),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_578),
.A2(n_539),
.B1(n_563),
.B2(n_522),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_541),
.B(n_399),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_446),
.B(n_399),
.Y(n_683)
);

AND2x4_ASAP7_75t_SL g684 ( 
.A(n_515),
.B(n_406),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_497),
.B(n_406),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_459),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_500),
.A2(n_390),
.B(n_401),
.C(n_400),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_567),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_503),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_400),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_503),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_490),
.B(n_177),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_511),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_497),
.B(n_390),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_582),
.B(n_400),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_487),
.A2(n_177),
.B1(n_180),
.B2(n_182),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_458),
.B(n_179),
.C(n_280),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_478),
.B(n_401),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_511),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_565),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_570),
.B(n_401),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_446),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_456),
.B(n_404),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_517),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_467),
.B(n_401),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_536),
.B(n_179),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_402),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_456),
.B(n_405),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_515),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_568),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_570),
.B(n_402),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_488),
.B(n_402),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_543),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_570),
.B(n_402),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_573),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_535),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_537),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_570),
.B(n_405),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_456),
.B(n_482),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_405),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_515),
.B(n_405),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_536),
.B(n_180),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_524),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_572),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_524),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_451),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_529),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_451),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_515),
.B(n_560),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_482),
.B(n_405),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_487),
.B(n_405),
.Y(n_732)
);

BUFx8_ASAP7_75t_L g733 ( 
.A(n_487),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_487),
.B(n_405),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_487),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_482),
.B(n_182),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_536),
.B(n_271),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_536),
.B(n_537),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_549),
.A2(n_301),
.B1(n_271),
.B2(n_274),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_487),
.A2(n_552),
.B1(n_556),
.B2(n_583),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_552),
.A2(n_556),
.B1(n_583),
.B2(n_560),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_552),
.B(n_274),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_552),
.B(n_276),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_529),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_624),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_663),
.B(n_492),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_603),
.B(n_472),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_616),
.B(n_552),
.Y(n_748)
);

BUFx8_ASAP7_75t_L g749 ( 
.A(n_642),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_616),
.B(n_552),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_606),
.B(n_579),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_643),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_663),
.B(n_491),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_621),
.B(n_537),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_639),
.A2(n_544),
.B(n_550),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_621),
.B(n_537),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_621),
.B(n_537),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_681),
.A2(n_554),
.B(n_558),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_685),
.B(n_512),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_613),
.A2(n_550),
.B(n_475),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_618),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_618),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_639),
.A2(n_502),
.B(n_452),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_583),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_735),
.B(n_587),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_716),
.B(n_462),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_656),
.A2(n_720),
.B(n_597),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_623),
.B(n_585),
.Y(n_769)
);

AOI21xp33_ASAP7_75t_L g770 ( 
.A1(n_714),
.A2(n_502),
.B(n_485),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_617),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_600),
.A2(n_530),
.B(n_452),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_628),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_593),
.B(n_462),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_601),
.B(n_694),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_713),
.B(n_608),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_608),
.B(n_583),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_720),
.A2(n_475),
.B(n_476),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_600),
.A2(n_530),
.B(n_485),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_627),
.A2(n_504),
.B(n_479),
.C(n_581),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_650),
.A2(n_651),
.B(n_595),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_622),
.B(n_465),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_610),
.B(n_670),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_628),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_725),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_609),
.A2(n_504),
.B1(n_475),
.B2(n_581),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_682),
.B(n_583),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_655),
.A2(n_532),
.B(n_486),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_627),
.B(n_462),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_662),
.A2(n_619),
.B(n_612),
.C(n_598),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_657),
.B(n_476),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_738),
.A2(n_476),
.B(n_479),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_632),
.B(n_479),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_669),
.B(n_504),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_738),
.A2(n_553),
.B(n_555),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_622),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_686),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_625),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_711),
.B(n_630),
.Y(n_799)
);

OAI321xp33_ASAP7_75t_L g800 ( 
.A1(n_697),
.A2(n_258),
.A3(n_257),
.B1(n_252),
.B2(n_262),
.C(n_278),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_640),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_553),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_589),
.A2(n_553),
.B(n_555),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_589),
.A2(n_555),
.B(n_562),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_674),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_666),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_621),
.B(n_585),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_590),
.A2(n_562),
.B(n_575),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_623),
.B(n_585),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_671),
.B(n_562),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_668),
.A2(n_575),
.B(n_581),
.C(n_527),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_631),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_575),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_725),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_590),
.A2(n_510),
.B(n_486),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_648),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_594),
.A2(n_516),
.B(n_506),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_604),
.A2(n_509),
.B1(n_506),
.B2(n_580),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_621),
.B(n_585),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_659),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_695),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_668),
.A2(n_527),
.B(n_510),
.C(n_580),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_679),
.B(n_465),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_R g824 ( 
.A(n_620),
.B(n_585),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_689),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_679),
.B(n_683),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_623),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_662),
.A2(n_521),
.B(n_566),
.C(n_557),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_683),
.A2(n_525),
.B(n_574),
.C(n_566),
.Y(n_829)
);

BUFx12f_ASAP7_75t_L g830 ( 
.A(n_644),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_655),
.A2(n_507),
.B(n_574),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_654),
.A2(n_301),
.B(n_276),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_602),
.B(n_605),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_695),
.B(n_509),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_644),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_690),
.B(n_516),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_645),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_623),
.B(n_534),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_698),
.B(n_532),
.Y(n_839)
);

OAI321xp33_ASAP7_75t_L g840 ( 
.A1(n_629),
.A2(n_299),
.A3(n_292),
.B1(n_297),
.B2(n_538),
.C(n_557),
.Y(n_840)
);

OAI321xp33_ASAP7_75t_L g841 ( 
.A1(n_676),
.A2(n_154),
.A3(n_195),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_706),
.B(n_534),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_693),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_661),
.A2(n_561),
.B(n_534),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_731),
.A2(n_561),
.B(n_587),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_652),
.B(n_280),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_680),
.A2(n_561),
.B1(n_587),
.B2(n_289),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_633),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_695),
.B(n_587),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_638),
.B(n_289),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_614),
.B(n_287),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_633),
.B(n_621),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_661),
.A2(n_665),
.B(n_664),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_700),
.B(n_287),
.Y(n_854)
);

AO21x1_ASAP7_75t_L g855 ( 
.A1(n_736),
.A2(n_217),
.B(n_195),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_664),
.A2(n_286),
.B(n_283),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_633),
.B(n_286),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_633),
.B(n_283),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_673),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_739),
.B(n_282),
.C(n_264),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_736),
.A2(n_217),
.B(n_195),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_675),
.A2(n_259),
.B(n_248),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_678),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_710),
.B(n_245),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_730),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_635),
.B(n_240),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_615),
.B(n_230),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_225),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_735),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_731),
.A2(n_221),
.B(n_220),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_675),
.A2(n_704),
.B(n_709),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_699),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_710),
.B(n_9),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_658),
.A2(n_218),
.B(n_213),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_612),
.A2(n_11),
.B(n_14),
.C(n_16),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_192),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_691),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_592),
.B(n_16),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_730),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_611),
.B(n_205),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_611),
.B(n_212),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_704),
.A2(n_195),
.B(n_154),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_709),
.A2(n_217),
.B(n_195),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_684),
.B(n_17),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_619),
.A2(n_217),
.B1(n_154),
.B2(n_25),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_733),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_592),
.B(n_17),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_730),
.A2(n_217),
.B1(n_25),
.B2(n_26),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_718),
.A2(n_217),
.B(n_79),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_705),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_686),
.B(n_18),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_626),
.B(n_27),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_637),
.A2(n_28),
.B(n_33),
.C(n_34),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_588),
.B(n_33),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_634),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_722),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_596),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_SL g899 ( 
.A(n_647),
.B(n_34),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_724),
.A2(n_91),
.B(n_148),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_677),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_687),
.A2(n_98),
.B(n_147),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_726),
.A2(n_90),
.B(n_141),
.Y(n_903)
);

AO21x1_ASAP7_75t_L g904 ( 
.A1(n_701),
.A2(n_89),
.B(n_139),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_728),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_641),
.A2(n_38),
.B(n_44),
.C(n_45),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_744),
.A2(n_105),
.B(n_134),
.Y(n_907)
);

CKINVDCx11_ASAP7_75t_R g908 ( 
.A(n_686),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_599),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_649),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_107),
.B(n_132),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_729),
.A2(n_65),
.B(n_110),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_646),
.B(n_49),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_672),
.B(n_50),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_740),
.B(n_50),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_719),
.A2(n_721),
.B(n_672),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_688),
.A2(n_121),
.B(n_149),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_SL g918 ( 
.A1(n_902),
.A2(n_591),
.B(n_688),
.C(n_723),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_752),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_783),
.B(n_607),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_765),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_835),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_796),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_758),
.A2(n_692),
.B(n_741),
.C(n_740),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_790),
.A2(n_741),
.B(n_696),
.C(n_715),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_826),
.A2(n_708),
.B(n_712),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_833),
.A2(n_751),
.B1(n_748),
.B2(n_750),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_781),
.A2(n_707),
.B(n_737),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_747),
.A2(n_742),
.B(n_743),
.C(n_734),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_819),
.A2(n_667),
.B(n_660),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_771),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_886),
.B(n_732),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_761),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_837),
.A2(n_733),
.B1(n_653),
.B2(n_53),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_784),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_830),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_775),
.B(n_776),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_768),
.A2(n_756),
.B(n_754),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_801),
.B(n_762),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_846),
.B(n_854),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_901),
.A2(n_872),
.B1(n_843),
.B2(n_820),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_798),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_879),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_784),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_799),
.B(n_896),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_749),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_749),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_799),
.B(n_821),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_821),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_816),
.B(n_825),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_901),
.A2(n_812),
.B1(n_915),
.B2(n_905),
.Y(n_954)
);

OAI22x1_ASAP7_75t_L g955 ( 
.A1(n_888),
.A2(n_887),
.B1(n_878),
.B2(n_884),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_789),
.B(n_793),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_805),
.Y(n_957)
);

NAND2x1_ASAP7_75t_L g958 ( 
.A(n_797),
.B(n_827),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_746),
.B(n_897),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_897),
.B(n_851),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_757),
.B(n_756),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_884),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_915),
.A2(n_894),
.B1(n_873),
.B2(n_813),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_878),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_802),
.B(n_877),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_851),
.B(n_832),
.Y(n_966)
);

AOI222xp33_ASAP7_75t_L g967 ( 
.A1(n_899),
.A2(n_887),
.B1(n_841),
.B2(n_873),
.C1(n_840),
.C2(n_910),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_895),
.A2(n_885),
.B(n_906),
.C(n_875),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_879),
.B(n_784),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_784),
.B(n_785),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_782),
.B(n_764),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_774),
.B(n_791),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_834),
.Y(n_973)
);

OR2x2_ASAP7_75t_SL g974 ( 
.A(n_860),
.B(n_865),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_785),
.B(n_814),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_773),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_774),
.A2(n_753),
.B1(n_849),
.B2(n_791),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_807),
.A2(n_836),
.B(n_823),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_797),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_773),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_891),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_857),
.A2(n_858),
.B(n_809),
.C(n_769),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_898),
.B(n_767),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_834),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_810),
.A2(n_759),
.B1(n_913),
.B2(n_893),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_831),
.A2(n_845),
.B(n_788),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_SL g988 ( 
.A1(n_892),
.A2(n_794),
.B(n_895),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_815),
.A2(n_817),
.B(n_792),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_865),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_874),
.B(n_892),
.C(n_870),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_828),
.A2(n_800),
.B(n_767),
.C(n_794),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_797),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_850),
.A2(n_867),
.B(n_811),
.C(n_866),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_787),
.A2(n_871),
.B(n_853),
.C(n_849),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_795),
.A2(n_808),
.B(n_804),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_777),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_803),
.A2(n_760),
.B(n_778),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_814),
.B(n_797),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_824),
.B(n_857),
.C(n_858),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_859),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_863),
.B(n_890),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_839),
.B(n_898),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_869),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_824),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_842),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_864),
.A2(n_876),
.B1(n_909),
.B2(n_868),
.Y(n_1007)
);

CKINVDCx6p67_ASAP7_75t_R g1008 ( 
.A(n_914),
.Y(n_1008)
);

CKINVDCx8_ASAP7_75t_R g1009 ( 
.A(n_770),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_818),
.A2(n_829),
.B(n_822),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_856),
.B(n_848),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_755),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_852),
.A2(n_780),
.B(n_916),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_827),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_883),
.A2(n_889),
.B(n_881),
.C(n_880),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_763),
.A2(n_882),
.B(n_772),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_848),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_766),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_R g1019 ( 
.A(n_844),
.B(n_904),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_862),
.B(n_838),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_779),
.B(n_847),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_903),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_SL g1023 ( 
.A(n_766),
.B(n_907),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_917),
.A2(n_911),
.B(n_912),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_752),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_783),
.A2(n_826),
.B1(n_833),
.B2(n_751),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_783),
.A2(n_826),
.B1(n_833),
.B2(n_751),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_801),
.A2(n_468),
.B1(n_461),
.B2(n_478),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_796),
.B(n_307),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_826),
.A2(n_636),
.B(n_783),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_SL g1031 ( 
.A(n_830),
.B(n_461),
.Y(n_1031)
);

AO32x1_ASAP7_75t_L g1032 ( 
.A1(n_910),
.A2(n_681),
.A3(n_818),
.B1(n_786),
.B2(n_847),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_796),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_826),
.A2(n_636),
.B(n_783),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_752),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_783),
.B(n_833),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_830),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_752),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_765),
.B(n_879),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_835),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_745),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_SL g1042 ( 
.A1(n_878),
.A2(n_674),
.B1(n_468),
.B2(n_461),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_783),
.B(n_449),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_796),
.B(n_307),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_745),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_747),
.A2(n_681),
.B(n_783),
.C(n_489),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1046),
.A2(n_1034),
.B(n_1030),
.Y(n_1047)
);

BUFx10_ASAP7_75t_L g1048 ( 
.A(n_949),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_952),
.B(n_984),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_SL g1050 ( 
.A(n_922),
.B(n_1040),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_1015),
.A2(n_985),
.A3(n_927),
.B(n_986),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1026),
.A2(n_1027),
.B1(n_1036),
.B2(n_972),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_985),
.A2(n_927),
.A3(n_1021),
.B(n_1010),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1036),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_919),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_948),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_983),
.B(n_943),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1024),
.A2(n_918),
.B(n_1023),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_991),
.A2(n_988),
.B(n_924),
.C(n_968),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_957),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_933),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_930),
.A2(n_954),
.A3(n_978),
.B(n_996),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_939),
.Y(n_1063)
);

BUFx2_ASAP7_75t_R g1064 ( 
.A(n_950),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1028),
.A2(n_963),
.B1(n_977),
.B2(n_1043),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1029),
.B(n_1044),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_963),
.A2(n_937),
.B1(n_959),
.B2(n_935),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_973),
.B(n_971),
.Y(n_1068)
);

AO32x2_ASAP7_75t_L g1069 ( 
.A1(n_954),
.A2(n_944),
.A3(n_990),
.B1(n_1042),
.B2(n_1032),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_1033),
.Y(n_1070)
);

AOI211x1_ASAP7_75t_L g1071 ( 
.A1(n_944),
.A2(n_953),
.B(n_920),
.C(n_965),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_931),
.B(n_964),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_953),
.A2(n_956),
.B1(n_1008),
.B2(n_1007),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_956),
.A2(n_1022),
.B(n_929),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_967),
.A2(n_955),
.B1(n_960),
.B2(n_966),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_923),
.B(n_1003),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_992),
.A2(n_994),
.B(n_925),
.C(n_982),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_995),
.A2(n_989),
.A3(n_1013),
.B(n_998),
.Y(n_1078)
);

O2A1O1Ixp5_ASAP7_75t_L g1079 ( 
.A1(n_932),
.A2(n_941),
.B(n_1020),
.C(n_961),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_928),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_942),
.B(n_962),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_945),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1003),
.B(n_973),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_965),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_936),
.A2(n_1012),
.B1(n_951),
.B2(n_974),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1006),
.A2(n_1005),
.B1(n_1009),
.B2(n_1025),
.Y(n_1086)
);

AO22x2_ASAP7_75t_L g1087 ( 
.A1(n_1006),
.A2(n_1000),
.B1(n_997),
.B2(n_981),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_926),
.A2(n_1032),
.B(n_1016),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1031),
.A2(n_1035),
.B1(n_1038),
.B2(n_997),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_928),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_987),
.B(n_1001),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1032),
.A2(n_1004),
.B(n_975),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_934),
.B(n_969),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_999),
.A2(n_1011),
.B(n_958),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1014),
.A2(n_1017),
.B(n_970),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_934),
.B(n_969),
.Y(n_1096)
);

BUFx10_ASAP7_75t_L g1097 ( 
.A(n_938),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1002),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1004),
.A2(n_993),
.B(n_1018),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_976),
.A2(n_980),
.B(n_1004),
.Y(n_1100)
);

BUFx4_ASAP7_75t_SL g1101 ( 
.A(n_1037),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_979),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_921),
.A2(n_934),
.B1(n_1039),
.B2(n_946),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_921),
.A2(n_946),
.B1(n_1039),
.B2(n_979),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_979),
.A2(n_938),
.B1(n_947),
.B2(n_1041),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1045),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1019),
.A2(n_938),
.B(n_947),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_947),
.B(n_940),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1033),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1036),
.C(n_826),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1015),
.A2(n_855),
.A3(n_861),
.B(n_985),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1036),
.C(n_826),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_922),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1046),
.A2(n_826),
.B(n_1030),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_940),
.B(n_1036),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_928),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_940),
.B(n_1036),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_964),
.A2(n_478),
.B1(n_899),
.B2(n_654),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_967),
.B(n_1046),
.C(n_968),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1046),
.A2(n_826),
.B(n_1030),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_SL g1121 ( 
.A(n_964),
.B(n_478),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_919),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_949),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1026),
.A2(n_826),
.B1(n_1027),
.B2(n_1036),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_928),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_968),
.A2(n_518),
.B(n_988),
.C(n_1027),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_919),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_922),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_967),
.A2(n_470),
.B(n_464),
.Y(n_1129)
);

OAI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_964),
.A2(n_478),
.B1(n_899),
.B2(n_654),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_940),
.B(n_1036),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_943),
.B(n_593),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1036),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_940),
.B(n_1036),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_949),
.B(n_457),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_940),
.B(n_1036),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_943),
.B(n_593),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1046),
.A2(n_758),
.B(n_616),
.C(n_991),
.Y(n_1138)
);

OAI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_523),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1015),
.A2(n_855),
.A3(n_861),
.B(n_985),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_941),
.A2(n_1013),
.B(n_989),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_928),
.Y(n_1142)
);

BUFx4_ASAP7_75t_R g1143 ( 
.A(n_1037),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_919),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1018),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_943),
.B(n_593),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_963),
.A2(n_985),
.B(n_954),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_922),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_922),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_919),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1029),
.B(n_461),
.Y(n_1151)
);

AOI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_967),
.A2(n_470),
.B(n_464),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_SL g1153 ( 
.A1(n_963),
.A2(n_906),
.B1(n_681),
.B2(n_910),
.C(n_1026),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_984),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1027),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1046),
.A2(n_758),
.B(n_616),
.C(n_991),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1033),
.B(n_796),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1046),
.A2(n_758),
.B(n_616),
.C(n_991),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1046),
.A2(n_826),
.B(n_1030),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1029),
.B(n_461),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1026),
.A2(n_826),
.B1(n_1027),
.B2(n_1036),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_957),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_L g1163 ( 
.A1(n_968),
.A2(n_902),
.B(n_758),
.C(n_963),
.Y(n_1163)
);

NAND3x1_ASAP7_75t_L g1164 ( 
.A(n_1028),
.B(n_887),
.C(n_878),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_967),
.A2(n_470),
.B(n_464),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_919),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_940),
.B(n_1036),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1026),
.B(n_1027),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_943),
.B(n_593),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_922),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_957),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_1119),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1101),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1097),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1168),
.B(n_1124),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1072),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1091),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1060),
.Y(n_1178)
);

INVx6_ASAP7_75t_L g1179 ( 
.A(n_1097),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1055),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1119),
.A2(n_1147),
.B1(n_1075),
.B2(n_1139),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1113),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1070),
.Y(n_1184)
);

BUFx4f_ASAP7_75t_SL g1185 ( 
.A(n_1048),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1162),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1171),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1075),
.A2(n_1139),
.B1(n_1065),
.B2(n_1161),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1157),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1052),
.A2(n_1073),
.B1(n_1054),
.B2(n_1130),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1135),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1082),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1149),
.Y(n_1193)
);

BUFx8_ASAP7_75t_L g1194 ( 
.A(n_1143),
.Y(n_1194)
);

INVx4_ASAP7_75t_SL g1195 ( 
.A(n_1093),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_1063),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1121),
.A2(n_1057),
.B1(n_1066),
.B2(n_1115),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1109),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1123),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1118),
.A2(n_1085),
.B1(n_1136),
.B2(n_1167),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1081),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1123),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1117),
.A2(n_1134),
.B1(n_1131),
.B2(n_1169),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1132),
.A2(n_1137),
.B1(n_1146),
.B2(n_1056),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1121),
.A2(n_1164),
.B1(n_1086),
.B2(n_1089),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_1080),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1090),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1076),
.B(n_1084),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1128),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1148),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1067),
.A2(n_1068),
.B1(n_1087),
.B2(n_1083),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1125),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1122),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1170),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1087),
.A2(n_1133),
.B1(n_1159),
.B2(n_1120),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1108),
.B(n_1127),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1144),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1089),
.A2(n_1166),
.B1(n_1150),
.B2(n_1049),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1153),
.A2(n_1158),
.B1(n_1156),
.B2(n_1138),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1154),
.Y(n_1220)
);

AO22x1_ASAP7_75t_L g1221 ( 
.A1(n_1049),
.A2(n_1142),
.B1(n_1116),
.B2(n_1100),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1153),
.A2(n_1059),
.B1(n_1103),
.B2(n_1077),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1098),
.B(n_1071),
.Y(n_1223)
);

INVx5_ASAP7_75t_L g1224 ( 
.A(n_1096),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1114),
.A2(n_1047),
.B1(n_1069),
.B2(n_1155),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1053),
.B(n_1106),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1116),
.Y(n_1227)
);

BUFx8_ASAP7_75t_SL g1228 ( 
.A(n_1154),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1154),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1064),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1069),
.A2(n_1096),
.B1(n_1092),
.B2(n_1088),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1069),
.A2(n_1096),
.B1(n_1163),
.B2(n_1095),
.Y(n_1232)
);

BUFx2_ASAP7_75t_SL g1233 ( 
.A(n_1145),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1094),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1050),
.A2(n_1053),
.B1(n_1105),
.B2(n_1112),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1104),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1102),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1078),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1099),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1110),
.A2(n_1074),
.B1(n_1058),
.B2(n_1053),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1079),
.Y(n_1242)
);

BUFx2_ASAP7_75t_R g1243 ( 
.A(n_1051),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1111),
.A2(n_1140),
.B1(n_1062),
.B2(n_1141),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1062),
.A2(n_1111),
.B(n_1140),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1062),
.A2(n_1119),
.B1(n_1075),
.B2(n_1129),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1078),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1078),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_967),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1115),
.B(n_1117),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1060),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1055),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_967),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1147),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1151),
.A2(n_1160),
.B(n_1126),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1132),
.B(n_1137),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1048),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1143),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1091),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1060),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1060),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1063),
.Y(n_1262)
);

NAND2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1068),
.B(n_821),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1151),
.A2(n_964),
.B1(n_955),
.B2(n_1160),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1143),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1139),
.A2(n_1163),
.B(n_1126),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1078),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1060),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1057),
.B(n_1070),
.Y(n_1269)
);

OAI22x1_ASAP7_75t_L g1270 ( 
.A1(n_1075),
.A2(n_1089),
.B1(n_1119),
.B2(n_964),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1143),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1101),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1055),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_967),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_967),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1101),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1119),
.A2(n_1168),
.B1(n_1151),
.B2(n_1160),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1147),
.Y(n_1278)
);

BUFx8_ASAP7_75t_L g1279 ( 
.A(n_1072),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1165),
.B2(n_967),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1132),
.B(n_1137),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1113),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1226),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1223),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1249),
.A2(n_1280),
.B1(n_1275),
.B2(n_1274),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1254),
.B(n_1278),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1245),
.A2(n_1266),
.B(n_1241),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1254),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1208),
.B(n_1278),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1225),
.B(n_1180),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1248),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1182),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1192),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1188),
.A2(n_1181),
.B1(n_1190),
.B2(n_1277),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1184),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1269),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1234),
.B(n_1235),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1213),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1248),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1234),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1239),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1225),
.B(n_1217),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1252),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1274),
.B2(n_1280),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1188),
.B(n_1181),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1273),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1267),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1247),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1247),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1264),
.A2(n_1237),
.B1(n_1275),
.B2(n_1253),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_SL g1311 ( 
.A(n_1255),
.B(n_1265),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1189),
.B(n_1246),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1216),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1237),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1231),
.B(n_1215),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1238),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1242),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1246),
.B(n_1211),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1220),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1265),
.B(n_1262),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1178),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1250),
.B(n_1197),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1231),
.B(n_1215),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1240),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1244),
.B(n_1190),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1211),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1232),
.A2(n_1219),
.B(n_1172),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1251),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1175),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1197),
.B(n_1200),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1218),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1262),
.B(n_1176),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1177),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1222),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1200),
.B(n_1203),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1259),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1260),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1232),
.B(n_1281),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1256),
.B(n_1261),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1198),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1205),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1236),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1236),
.B(n_1204),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1220),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1172),
.A2(n_1174),
.B(n_1263),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1183),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1270),
.A2(n_1221),
.B(n_1199),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1220),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1233),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1179),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1179),
.Y(n_1352)
);

BUFx5_ASAP7_75t_L g1353 ( 
.A(n_1229),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1268),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1212),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1224),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1195),
.A2(n_1224),
.B(n_1204),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1292),
.Y(n_1358)
);

AOI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1285),
.A2(n_1186),
.B1(n_1187),
.B2(n_1201),
.C(n_1191),
.Y(n_1359)
);

AOI21xp33_ASAP7_75t_L g1360 ( 
.A1(n_1304),
.A2(n_1279),
.B(n_1202),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1287),
.B(n_1257),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1294),
.A2(n_1194),
.B1(n_1183),
.B2(n_1282),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1294),
.A2(n_1271),
.B(n_1258),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1292),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1331),
.A2(n_1310),
.B(n_1305),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1340),
.B(n_1230),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1305),
.A2(n_1193),
.B(n_1227),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1330),
.A2(n_1173),
.B(n_1276),
.C(n_1272),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1325),
.B(n_1194),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1330),
.B(n_1279),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1293),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1347),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1296),
.B(n_1295),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1323),
.B(n_1318),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1287),
.B(n_1207),
.Y(n_1375)
);

AO32x2_ASAP7_75t_L g1376 ( 
.A1(n_1315),
.A2(n_1206),
.A3(n_1228),
.B1(n_1185),
.B2(n_1282),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1343),
.A2(n_1206),
.B(n_1185),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1338),
.B(n_1196),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1338),
.B(n_1214),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1335),
.A2(n_1209),
.B(n_1210),
.C(n_1336),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1316),
.A2(n_1324),
.B(n_1319),
.C(n_1326),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1288),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1343),
.A2(n_1318),
.B(n_1289),
.Y(n_1383)
);

AO32x2_ASAP7_75t_L g1384 ( 
.A1(n_1354),
.A2(n_1320),
.A3(n_1345),
.B1(n_1349),
.B2(n_1356),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1329),
.B(n_1290),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1290),
.B(n_1302),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1287),
.B(n_1302),
.Y(n_1387)
);

NAND4xp25_ASAP7_75t_SL g1388 ( 
.A(n_1319),
.B(n_1311),
.C(n_1313),
.D(n_1335),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1313),
.A2(n_1344),
.B(n_1342),
.C(n_1311),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1298),
.B(n_1303),
.Y(n_1390)
);

AND2x2_ASAP7_75t_SL g1391 ( 
.A(n_1328),
.B(n_1286),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1350),
.A2(n_1321),
.B(n_1341),
.C(n_1354),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1350),
.B(n_1284),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1328),
.A2(n_1346),
.B(n_1342),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1314),
.B(n_1284),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1300),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1314),
.B(n_1322),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1344),
.A2(n_1286),
.B(n_1327),
.C(n_1317),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_1339),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1328),
.A2(n_1355),
.B(n_1333),
.C(n_1349),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1357),
.B(n_1306),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1308),
.A2(n_1309),
.B(n_1332),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1387),
.B(n_1382),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1387),
.B(n_1300),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1382),
.B(n_1309),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1395),
.B(n_1308),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1358),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1364),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1399),
.B(n_1300),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1372),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1391),
.B(n_1300),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1371),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1391),
.B(n_1297),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1328),
.B1(n_1312),
.B2(n_1332),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1381),
.A2(n_1312),
.B1(n_1348),
.B2(n_1352),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1372),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1388),
.A2(n_1337),
.B1(n_1283),
.B2(n_1334),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1390),
.B(n_1307),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1392),
.B(n_1351),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1385),
.B(n_1291),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1402),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1402),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1393),
.B(n_1301),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1402),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1396),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1384),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1427),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1424),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1404),
.B(n_1401),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1429),
.B(n_1386),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.Y(n_1434)
);

OAI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1414),
.A2(n_1389),
.B1(n_1381),
.B2(n_1398),
.C(n_1362),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1425),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1429),
.B(n_1373),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1403),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1429),
.B(n_1397),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1427),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1415),
.A2(n_1394),
.B(n_1398),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1403),
.B(n_1383),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1384),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1415),
.B(n_1362),
.C(n_1380),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1405),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1407),
.Y(n_1450)
);

OAI211xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1416),
.A2(n_1368),
.B(n_1363),
.C(n_1370),
.Y(n_1451)
);

AOI211xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1410),
.A2(n_1360),
.B(n_1392),
.C(n_1375),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1406),
.Y(n_1453)
);

AOI211xp5_ASAP7_75t_L g1454 ( 
.A1(n_1416),
.A2(n_1375),
.B(n_1400),
.C(n_1367),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1407),
.Y(n_1455)
);

INVx5_ASAP7_75t_L g1456 ( 
.A(n_1428),
.Y(n_1456)
);

NAND2x1_ASAP7_75t_SL g1457 ( 
.A(n_1446),
.B(n_1413),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1440),
.B(n_1421),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1450),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1433),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1453),
.B(n_1406),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1439),
.B(n_1443),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1453),
.B(n_1408),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1450),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1456),
.B(n_1413),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1421),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1447),
.A2(n_1414),
.B1(n_1420),
.B2(n_1374),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1448),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1436),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1440),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1450),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1436),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1454),
.B(n_1422),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1433),
.B(n_1426),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1432),
.B(n_1419),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1432),
.B(n_1419),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1408),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1455),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1455),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1456),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1456),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1442),
.B(n_1412),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1456),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1474),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1460),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1449),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1460),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1465),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1463),
.B(n_1484),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1462),
.B(n_1483),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1462),
.B(n_1433),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1468),
.B(n_1442),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1465),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1468),
.B(n_1418),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1477),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1463),
.B(n_1449),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1477),
.Y(n_1507)
);

CKINVDCx16_ASAP7_75t_R g1508 ( 
.A(n_1466),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1484),
.B(n_1485),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1474),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1492),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1474),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1482),
.A2(n_1447),
.B1(n_1435),
.B2(n_1454),
.C(n_1430),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1469),
.B(n_1442),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1487),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1469),
.B(n_1438),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1438),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1488),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1458),
.B(n_1449),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1492),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1483),
.B(n_1433),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1458),
.B(n_1455),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1457),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1464),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1464),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1458),
.B(n_1454),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1486),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1466),
.B(n_1456),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1479),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1466),
.B(n_1447),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1486),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1470),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1502),
.B(n_1461),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1513),
.A2(n_1534),
.B(n_1504),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_SL g1539 ( 
.A(n_1526),
.B(n_1435),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1470),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1530),
.A2(n_1435),
.B(n_1452),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

NAND2x1_ASAP7_75t_L g1543 ( 
.A(n_1526),
.B(n_1491),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1535),
.B(n_1511),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

NAND4xp25_ASAP7_75t_SL g1548 ( 
.A(n_1509),
.B(n_1481),
.C(n_1478),
.D(n_1480),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1494),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1518),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1528),
.A2(n_1441),
.B(n_1430),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1498),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1495),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1506),
.B(n_1471),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1472),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1498),
.Y(n_1560)
);

OAI21xp33_ASAP7_75t_L g1561 ( 
.A1(n_1529),
.A2(n_1457),
.B(n_1452),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1506),
.B(n_1509),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1503),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1478),
.Y(n_1564)
);

NAND2x1_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1491),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1516),
.B(n_1478),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1418),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1529),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1524),
.B(n_1459),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1524),
.B(n_1459),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1554),
.B(n_1472),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1531),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_SL g1573 ( 
.A(n_1538),
.B(n_1451),
.C(n_1515),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1542),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1575)
);

AOI211xp5_ASAP7_75t_L g1576 ( 
.A1(n_1561),
.A2(n_1451),
.B(n_1531),
.C(n_1527),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1537),
.A2(n_1452),
.B(n_1527),
.C(n_1359),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

AOI21xp33_ASAP7_75t_L g1580 ( 
.A1(n_1537),
.A2(n_1444),
.B(n_1503),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1543),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1480),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1568),
.B(n_1480),
.Y(n_1583)
);

OAI32xp33_ASAP7_75t_L g1584 ( 
.A1(n_1554),
.A2(n_1501),
.A3(n_1521),
.B1(n_1445),
.B2(n_1525),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1560),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1563),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1555),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1481),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1501),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1567),
.B(n_1418),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1481),
.Y(n_1591)
);

OAI32xp33_ASAP7_75t_L g1592 ( 
.A1(n_1550),
.A2(n_1445),
.A3(n_1437),
.B1(n_1490),
.B2(n_1479),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1548),
.A2(n_1445),
.B(n_1505),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1577),
.A2(n_1562),
.B1(n_1546),
.B2(n_1536),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1572),
.A2(n_1570),
.B1(n_1569),
.B2(n_1565),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1575),
.B(n_1410),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1577),
.A2(n_1562),
.B1(n_1536),
.B2(n_1540),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1589),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1581),
.B(n_1540),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1573),
.A2(n_1549),
.B(n_1569),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1573),
.A2(n_1559),
.B1(n_1570),
.B2(n_1565),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1587),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1576),
.A2(n_1558),
.B1(n_1557),
.B2(n_1556),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1556),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

AOI221x1_ASAP7_75t_L g1611 ( 
.A1(n_1580),
.A2(n_1549),
.B1(n_1523),
.B2(n_1520),
.C(n_1514),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1592),
.A2(n_1430),
.B1(n_1441),
.B2(n_1512),
.C1(n_1510),
.C2(n_1533),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

AOI211xp5_ASAP7_75t_L g1615 ( 
.A1(n_1596),
.A2(n_1584),
.B(n_1595),
.C(n_1590),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1605),
.B(n_1590),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1601),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1585),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_R g1619 ( 
.A(n_1603),
.B(n_1586),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1609),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1604),
.B(n_1582),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1613),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1588),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1605),
.A2(n_1600),
.B(n_1611),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1614),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1608),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1599),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_SL g1628 ( 
.A(n_1624),
.B(n_1612),
.C(n_1602),
.Y(n_1628)
);

AOI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1624),
.A2(n_1598),
.B(n_1607),
.C(n_1606),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1620),
.B(n_1610),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1621),
.A2(n_1612),
.B(n_1583),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1617),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1623),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1622),
.B(n_1510),
.C(n_1494),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1630),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1628),
.A2(n_1626),
.B(n_1625),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_L g1638 ( 
.A(n_1632),
.B(n_1558),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1629),
.A2(n_1615),
.B(n_1619),
.C(n_1566),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1633),
.A2(n_1552),
.B(n_1512),
.C(n_1533),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_L g1641 ( 
.A1(n_1637),
.A2(n_1627),
.B(n_1631),
.C(n_1634),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1638),
.Y(n_1642)
);

AOI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1640),
.A2(n_1635),
.B(n_1566),
.C(n_1564),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1636),
.A2(n_1552),
.B1(n_1441),
.B2(n_1479),
.C(n_1490),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1552),
.Y(n_1645)
);

AOI322xp5_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1564),
.A3(n_1490),
.B1(n_1436),
.B2(n_1420),
.C1(n_1517),
.C2(n_1514),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1642),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1645),
.A2(n_1491),
.B1(n_1523),
.B2(n_1520),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1641),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1643),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1644),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1647),
.B(n_1379),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1648),
.A2(n_1646),
.B1(n_1491),
.B2(n_1489),
.C(n_1493),
.Y(n_1653)
);

AOI222xp33_ASAP7_75t_L g1654 ( 
.A1(n_1651),
.A2(n_1517),
.B1(n_1507),
.B2(n_1505),
.C1(n_1436),
.C2(n_1434),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1652),
.Y(n_1655)
);

AO22x2_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1649),
.B1(n_1650),
.B2(n_1651),
.Y(n_1656)
);

AOI22x1_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1654),
.B1(n_1653),
.B2(n_1507),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1532),
.B1(n_1491),
.B2(n_1370),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1491),
.B1(n_1532),
.B2(n_1493),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1659),
.A2(n_1366),
.B(n_1493),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1659),
.Y(n_1661)
);

OAI21xp33_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1489),
.B(n_1378),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1660),
.A2(n_1473),
.B(n_1472),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1489),
.B1(n_1467),
.B2(n_1459),
.Y(n_1664)
);

XNOR2xp5_ASAP7_75t_L g1665 ( 
.A(n_1662),
.B(n_1376),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1664),
.A2(n_1665),
.B1(n_1434),
.B2(n_1431),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1377),
.B1(n_1369),
.B2(n_1476),
.Y(n_1667)
);


endmodule