module fake_netlist_5_1293_n_1451 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1451);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1451;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_317),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_57),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_203),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_88),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_24),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_217),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_252),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_13),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_114),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_178),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_22),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_327),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_156),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_12),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_111),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_142),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_105),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_2),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_151),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_277),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_179),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_207),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_353),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_265),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_183),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_248),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_110),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_204),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_60),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_219),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_275),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_271),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_19),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_154),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_79),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_196),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_345),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_262),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_162),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_184),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_113),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_34),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_309),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_27),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_116),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_123),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_9),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_59),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_75),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_133),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_92),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_6),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_246),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_190),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_325),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_322),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_284),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_34),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_242),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_126),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_20),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_231),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_318),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_281),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_104),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_100),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_233),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_50),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_291),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_65),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_109),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_238),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_26),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_119),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_19),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_191),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_57),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_108),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_59),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_297),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_13),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_43),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_256),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_72),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_192),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_296),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_276),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_295),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_141),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_76),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_170),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_323),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_215),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_28),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_27),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_93),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_115),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_266),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_44),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_38),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_332),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_42),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_143),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_65),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_99),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_272),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_11),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_10),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_350),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_26),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_240),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_55),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_351),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_362),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_164),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_225),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_340),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_2),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_346),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_85),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_274),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_168),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_319),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_118),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_166),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_132),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_198),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_68),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_152),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_51),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_165),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_42),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_226),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_344),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_316),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_83),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_359),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_106),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_53),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_282),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_159),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_347),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_321),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_343),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_349),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_239),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_122),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_12),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_280),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_313),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_14),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_241),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_247),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_209),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_176),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_169),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_117),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_91),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_18),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_158),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_80),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_283),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_11),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_16),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_155),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_315),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_15),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_365),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_188),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_254),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_97),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_357),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_352),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_485),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_386),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_419),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_386),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_381),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_475),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_539),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_376),
.B(n_0),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_503),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_376),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_539),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_419),
.B(n_0),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_539),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_384),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_1),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_383),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_432),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_432),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_418),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_421),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_385),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_396),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_404),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_411),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_445),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_460),
.B(n_1),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_459),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_372),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_414),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_502),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_3),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_379),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_371),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_415),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_417),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_477),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_487),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_391),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_402),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_375),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_377),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_374),
.B(n_3),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_416),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_389),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_423),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_410),
.B(n_4),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_424),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_444),
.B(n_393),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_505),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_401),
.B(n_496),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_378),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_380),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_382),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_388),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_390),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_392),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_422),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_426),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_435),
.B(n_443),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_427),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_413),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_428),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_450),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_397),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_452),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_398),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_429),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_394),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_425),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_399),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_454),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_430),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_400),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_403),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_456),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_457),
.B(n_4),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_434),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_436),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_408),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_394),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_409),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_441),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_438),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_439),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_442),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_394),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_446),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_458),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_462),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_447),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_474),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_554),
.B(n_387),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_623),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_556),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_596),
.B(n_612),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_564),
.B(n_412),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_549),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_614),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_585),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_561),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_549),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_598),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_616),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_571),
.B(n_420),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_624),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_572),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_578),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_635),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_626),
.B(n_406),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_593),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_635),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_594),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_578),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_573),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_574),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_581),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_642),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_586),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_647),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_607),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_580),
.B(n_406),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_587),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_595),
.B(n_431),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_584),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_609),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_642),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_610),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_611),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_619),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_599),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_584),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_649),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_621),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_625),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_601),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_628),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_629),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_636),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_639),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_640),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_590),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_590),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_615),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_644),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_617),
.B(n_461),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_566),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_645),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_622),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_R g712 ( 
.A(n_627),
.B(n_437),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_602),
.B(n_431),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_646),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_591),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_591),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_569),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_632),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_494),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_633),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_608),
.B(n_497),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_637),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_570),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_597),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_634),
.A2(n_480),
.B(n_476),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_575),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_577),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_597),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_588),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_589),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_592),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_712),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_727),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_709),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_709),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_709),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_683),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_672),
.B(n_551),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_662),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_653),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_730),
.B(n_550),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_672),
.B(n_582),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_709),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_729),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_725),
.B(n_500),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_685),
.B(n_719),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_713),
.A2(n_567),
.B1(n_600),
.B2(n_631),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_670),
.B(n_641),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_705),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_SL g757 ( 
.A(n_681),
.B(n_613),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_671),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_732),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_731),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_650),
.B(n_643),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_674),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_692),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_652),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_654),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_682),
.Y(n_768)
);

BUFx6f_ASAP7_75t_SL g769 ( 
.A(n_692),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_655),
.B(n_648),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_664),
.B(n_562),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_718),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_687),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_708),
.B(n_613),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_689),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_666),
.B(n_565),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_721),
.B(n_603),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_690),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_660),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_721),
.B(n_604),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_679),
.B(n_654),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_552),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_695),
.B(n_553),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_691),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_668),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_667),
.Y(n_787)
);

BUFx4f_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_696),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_656),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_701),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_666),
.B(n_576),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

AND2x6_ASAP7_75t_L g794 ( 
.A(n_702),
.B(n_373),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_707),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_669),
.B(n_583),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_676),
.B(n_677),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_658),
.B(n_555),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_669),
.B(n_394),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_714),
.B(n_557),
.Y(n_800)
);

INVx4_ASAP7_75t_SL g801 ( 
.A(n_725),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_691),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_698),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_698),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_692),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_698),
.B(n_373),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_669),
.B(n_394),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_699),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_662),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_656),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_677),
.B(n_618),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_699),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_700),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_678),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_678),
.B(n_618),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_717),
.B(n_440),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_688),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_688),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_700),
.Y(n_819)
);

INVx6_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_688),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_680),
.B(n_373),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_710),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_710),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_703),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_703),
.B(n_531),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_771),
.B(n_703),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_771),
.B(n_680),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_761),
.B(n_684),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_761),
.B(n_684),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_770),
.B(n_697),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_737),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_751),
.B(n_697),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_825),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_785),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_803),
.B(n_706),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_744),
.B(n_816),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_816),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_774),
.B(n_706),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_788),
.A2(n_509),
.B1(n_533),
.B2(n_508),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_765),
.B(n_776),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_803),
.B(n_711),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_804),
.B(n_711),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_826),
.B(n_720),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_826),
.B(n_720),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_722),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_796),
.B(n_722),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_749),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_735),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_798),
.B(n_620),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_796),
.B(n_733),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_741),
.B(n_620),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_735),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_820),
.B(n_693),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_741),
.B(n_659),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_742),
.B(n_733),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_742),
.B(n_733),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_752),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_786),
.B(n_694),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_752),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_746),
.B(n_481),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_746),
.A2(n_723),
.B(n_728),
.C(n_717),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_767),
.B(n_780),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_767),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_777),
.B(n_659),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_754),
.A2(n_478),
.B1(n_513),
.B2(n_465),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_781),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_785),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_780),
.B(n_488),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_759),
.Y(n_870)
);

AND2x6_ASAP7_75t_SL g871 ( 
.A(n_815),
.B(n_657),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_755),
.B(n_630),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_762),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_817),
.B(n_492),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_745),
.Y(n_875)
);

OAI21xp33_ASAP7_75t_L g876 ( 
.A1(n_783),
.A2(n_482),
.B(n_479),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_764),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_788),
.A2(n_750),
.B1(n_754),
.B2(n_768),
.Y(n_878)
);

AND2x4_ASAP7_75t_SL g879 ( 
.A(n_793),
.B(n_657),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_817),
.B(n_498),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_743),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_818),
.B(n_504),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_818),
.B(n_506),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_792),
.B(n_630),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_750),
.A2(n_535),
.B1(n_515),
.B2(n_520),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_754),
.A2(n_517),
.B1(n_543),
.B2(n_522),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_773),
.Y(n_888)
);

NAND2x1_ASAP7_75t_L g889 ( 
.A(n_821),
.B(n_373),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_758),
.B(n_723),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_821),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_768),
.B(n_559),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_775),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_801),
.A2(n_510),
.B1(n_527),
.B2(n_525),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_748),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_800),
.B(n_663),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_822),
.B(n_493),
.C(n_483),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_778),
.B(n_789),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_791),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_784),
.A2(n_548),
.B1(n_568),
.B2(n_560),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_802),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_808),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_784),
.A2(n_560),
.B1(n_568),
.B2(n_559),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_801),
.A2(n_536),
.B1(n_547),
.B2(n_545),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_786),
.B(n_716),
.Y(n_906)
);

INVx8_ASAP7_75t_L g907 ( 
.A(n_769),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_785),
.B(n_728),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_736),
.B(n_663),
.Y(n_909)
);

BUFx8_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_795),
.B(n_665),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_819),
.B(n_734),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_756),
.B(n_726),
.Y(n_913)
);

BUFx6f_ASAP7_75t_SL g914 ( 
.A(n_793),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_812),
.B(n_734),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_745),
.B(n_665),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_812),
.B(n_813),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_763),
.B(n_668),
.Y(n_918)
);

OR2x6_ASAP7_75t_L g919 ( 
.A(n_820),
.B(n_395),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_748),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_812),
.B(n_449),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_878),
.A2(n_824),
.B(n_823),
.C(n_799),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_835),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_887),
.B(n_757),
.C(n_811),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_881),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_854),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_917),
.A2(n_740),
.B(n_738),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_828),
.B(n_814),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_838),
.B(n_805),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_867),
.B(n_756),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_827),
.B(n_801),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_839),
.B(n_760),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_R g933 ( 
.A(n_913),
.B(n_809),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_835),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_832),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_892),
.B(n_523),
.C(n_514),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_R g937 ( 
.A(n_859),
.B(n_772),
.Y(n_937)
);

INVx6_ASAP7_75t_L g938 ( 
.A(n_854),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_914),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_851),
.B(n_782),
.Y(n_940)
);

BUFx12f_ASAP7_75t_SL g941 ( 
.A(n_854),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_835),
.Y(n_942)
);

AOI211xp5_ASAP7_75t_L g943 ( 
.A1(n_885),
.A2(n_760),
.B(n_797),
.C(n_534),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_848),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_866),
.A2(n_820),
.B1(n_715),
.B2(n_724),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_906),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_856),
.B(n_782),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_902),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_857),
.B(n_813),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_870),
.Y(n_950)
);

AND3x2_ASAP7_75t_SL g951 ( 
.A(n_901),
.B(n_661),
.C(n_766),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_914),
.Y(n_952)
);

AND2x2_ASAP7_75t_SL g953 ( 
.A(n_879),
.B(n_829),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_847),
.A2(n_807),
.B(n_799),
.C(n_787),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_871),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_873),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_834),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_877),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_SL g959 ( 
.A(n_830),
.B(n_715),
.C(n_675),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_SL g960 ( 
.A(n_831),
.B(n_724),
.C(n_675),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_834),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_834),
.B(n_779),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_916),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_844),
.B(n_661),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_845),
.B(n_813),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_861),
.B(n_790),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_SL g967 ( 
.A(n_852),
.B(n_538),
.C(n_526),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_919),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_868),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_836),
.B(n_810),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_833),
.B(n_738),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_890),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_888),
.A2(n_740),
.B1(n_747),
.B2(n_739),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_907),
.B(n_739),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_903),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_911),
.B(n_542),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_R g977 ( 
.A(n_841),
.B(n_907),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_893),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_868),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_900),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_842),
.B(n_843),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_908),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_919),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_SL g984 ( 
.A(n_846),
.B(n_451),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_895),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_897),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_899),
.B(n_747),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_849),
.B(n_853),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_875),
.B(n_739),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_923),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_971),
.B(n_890),
.Y(n_991)
);

OAI21x1_ASAP7_75t_SL g992 ( 
.A1(n_954),
.A2(n_862),
.B(n_869),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_981),
.B(n_883),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_981),
.B(n_872),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_946),
.B(n_918),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_928),
.B(n_837),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_935),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_SL g998 ( 
.A1(n_964),
.A2(n_850),
.B(n_901),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_932),
.B(n_909),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_931),
.A2(n_874),
.B(n_882),
.C(n_880),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_940),
.B(n_886),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_987),
.A2(n_905),
.B1(n_894),
.B2(n_840),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_931),
.A2(n_863),
.B(n_884),
.Y(n_1003)
);

OAI22x1_ASAP7_75t_L g1004 ( 
.A1(n_951),
.A2(n_904),
.B1(n_855),
.B2(n_865),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_930),
.B(n_904),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_987),
.A2(n_920),
.B1(n_858),
.B2(n_864),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_941),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_944),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_947),
.A2(n_940),
.B(n_949),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_982),
.B(n_947),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_922),
.A2(n_915),
.B(n_891),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_949),
.A2(n_921),
.B(n_860),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_927),
.A2(n_807),
.B(n_889),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_970),
.A2(n_912),
.B(n_898),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_934),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_SL g1016 ( 
.A(n_923),
.B(n_919),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_988),
.A2(n_912),
.B(n_896),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_950),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_956),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_938),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_958),
.B(n_876),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_970),
.A2(n_463),
.B1(n_464),
.B2(n_455),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_988),
.A2(n_394),
.B(n_806),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_924),
.A2(n_907),
.B(n_405),
.C(n_491),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_959),
.B(n_960),
.C(n_945),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_SL g1026 ( 
.A1(n_966),
.A2(n_78),
.B(n_77),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_969),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_978),
.B(n_466),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_980),
.B(n_467),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_969),
.A2(n_806),
.B(n_794),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_979),
.A2(n_986),
.B(n_985),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_948),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_966),
.A2(n_753),
.B(n_405),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_975),
.A2(n_753),
.B(n_806),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_965),
.A2(n_806),
.B(n_753),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_985),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_986),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_938),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_963),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_942),
.A2(n_753),
.B(n_405),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_943),
.A2(n_405),
.B(n_491),
.C(n_395),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_937),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_973),
.A2(n_989),
.B(n_976),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_972),
.A2(n_468),
.B1(n_472),
.B2(n_471),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_967),
.A2(n_499),
.B(n_433),
.C(n_7),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_962),
.B(n_484),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_997),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_1026),
.A2(n_961),
.B(n_945),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1008),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_990),
.B(n_961),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_1025),
.A2(n_953),
.B1(n_962),
.B2(n_984),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_1038),
.B(n_974),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_1041),
.A2(n_983),
.A3(n_951),
.B(n_936),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1010),
.B(n_979),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_1039),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_998),
.A2(n_933),
.B1(n_955),
.B2(n_929),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_1031),
.A2(n_934),
.B(n_968),
.Y(n_1058)
);

BUFx2_ASAP7_75t_R g1059 ( 
.A(n_1042),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_990),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1009),
.A2(n_929),
.B(n_794),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_1024),
.A2(n_977),
.B(n_974),
.C(n_82),
.Y(n_1062)
);

AND2x2_ASAP7_75t_SL g1063 ( 
.A(n_1025),
.B(n_994),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1001),
.A2(n_993),
.B1(n_996),
.B2(n_1018),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1031),
.A2(n_974),
.B(n_957),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_991),
.A2(n_957),
.B(n_926),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_1038),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_1023),
.A2(n_489),
.B(n_486),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1019),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1013),
.A2(n_957),
.B(n_491),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1043),
.A2(n_925),
.B(n_490),
.C(n_511),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_1012),
.A2(n_491),
.B(n_395),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_995),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1002),
.A2(n_952),
.B1(n_939),
.B2(n_501),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1020),
.B(n_81),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_1024),
.A2(n_910),
.B(n_499),
.C(n_433),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1007),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1034),
.A2(n_794),
.B(n_501),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1032),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_1000),
.A2(n_794),
.B(n_512),
.C(n_516),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1023),
.A2(n_501),
.B(n_395),
.Y(n_1081)
);

AND2x4_ASAP7_75t_SL g1082 ( 
.A(n_1027),
.B(n_910),
.Y(n_1082)
);

CKINVDCx11_ASAP7_75t_R g1083 ( 
.A(n_1042),
.Y(n_1083)
);

CKINVDCx11_ASAP7_75t_R g1084 ( 
.A(n_1044),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1036),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_992),
.A2(n_518),
.B(n_501),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1037),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_L g1088 ( 
.A(n_999),
.B(n_495),
.Y(n_1088)
);

INVxp33_ASAP7_75t_L g1089 ( 
.A(n_1005),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1015),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1046),
.B(n_519),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1003),
.A2(n_537),
.B(n_518),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1015),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1011),
.A2(n_1000),
.B(n_1017),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1006),
.A2(n_537),
.B(n_518),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1027),
.B(n_84),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1021),
.B(n_521),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1014),
.A2(n_524),
.B(n_529),
.C(n_528),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1004),
.A2(n_530),
.B1(n_540),
.B2(n_532),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1041),
.A2(n_537),
.B1(n_546),
.B2(n_518),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_1045),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_1035),
.A2(n_1033),
.B(n_1040),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_1028),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1073),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1048),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1064),
.A2(n_1016),
.B(n_1029),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1060),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_SL g1109 ( 
.A(n_1057),
.B(n_1022),
.C(n_544),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_1083),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1074),
.A2(n_1064),
.B1(n_1099),
.B2(n_1089),
.C(n_1076),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1063),
.A2(n_546),
.B1(n_537),
.B2(n_1030),
.Y(n_1112)
);

AOI222xp33_ASAP7_75t_L g1113 ( 
.A1(n_1084),
.A2(n_546),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_1113)
);

INVx4_ASAP7_75t_SL g1114 ( 
.A(n_1067),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1057),
.A2(n_546),
.B1(n_1030),
.B2(n_10),
.Y(n_1115)
);

OAI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1074),
.A2(n_14),
.B(n_5),
.C(n_8),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1073),
.B(n_5),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1069),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_1103),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1079),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1059),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_SL g1122 ( 
.A(n_1052),
.B(n_15),
.C(n_16),
.Y(n_1122)
);

AND2x4_ASAP7_75t_SL g1123 ( 
.A(n_1067),
.B(n_86),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1060),
.B(n_87),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1055),
.B(n_17),
.Y(n_1125)
);

NOR3xp33_ASAP7_75t_SL g1126 ( 
.A(n_1066),
.B(n_17),
.C(n_18),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1085),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1047),
.B(n_20),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1053),
.B(n_89),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1059),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1087),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_SL g1132 ( 
.A(n_1071),
.B(n_21),
.C(n_22),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1093),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1056),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1067),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1077),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1090),
.Y(n_1137)
);

OAI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1091),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1053),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1101),
.A2(n_28),
.B1(n_23),
.B2(n_25),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1097),
.B(n_90),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1082),
.Y(n_1142)
);

AOI221xp5_ASAP7_75t_L g1143 ( 
.A1(n_1100),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1060),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_1053),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1100),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_1146)
);

OAI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1088),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_SL g1148 ( 
.A(n_1075),
.B(n_1055),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1058),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1101),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_1096),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1075),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1096),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1098),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.C(n_40),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1054),
.B(n_39),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1051),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1051),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_1068),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1049),
.Y(n_1161)
);

CKINVDCx8_ASAP7_75t_R g1162 ( 
.A(n_1068),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1054),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_SL g1164 ( 
.A(n_1061),
.B(n_41),
.Y(n_1164)
);

NAND2xp33_ASAP7_75t_R g1165 ( 
.A(n_1061),
.B(n_94),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1080),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1102),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1102),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1168)
);

AOI21xp33_ASAP7_75t_L g1169 ( 
.A1(n_1086),
.A2(n_48),
.B(n_49),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1086),
.B(n_50),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1062),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_1095),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1070),
.B(n_95),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1094),
.B(n_96),
.Y(n_1174)
);

AO21x2_ASAP7_75t_L g1175 ( 
.A1(n_1092),
.A2(n_101),
.B(n_98),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1072),
.B1(n_1081),
.B2(n_53),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1117),
.B(n_102),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1127),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1104),
.B(n_51),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1110),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1147),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1138),
.A2(n_1078),
.B1(n_54),
.B2(n_56),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1151),
.B(n_103),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1122),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1151),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1125),
.B(n_1134),
.Y(n_1186)
);

OAI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1111),
.A2(n_1132),
.B1(n_1113),
.B2(n_1141),
.C(n_1140),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1148),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1107),
.A2(n_1169),
.B(n_1149),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1105),
.B(n_62),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1151),
.A2(n_112),
.B(n_107),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1152),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1143),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1146),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1129),
.B(n_120),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1136),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1119),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1137),
.B(n_70),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1150),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1131),
.B(n_73),
.Y(n_1200)
);

OAI21xp33_ASAP7_75t_L g1201 ( 
.A1(n_1167),
.A2(n_74),
.B(n_121),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1168),
.A2(n_74),
.B1(n_124),
.B2(n_125),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1153),
.B(n_127),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1129),
.A2(n_128),
.B(n_129),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1155),
.B(n_1106),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1164),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1139),
.B(n_135),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1119),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1139),
.B(n_139),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1115),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1118),
.B(n_146),
.Y(n_1211)
);

AOI222xp33_ASAP7_75t_L g1212 ( 
.A1(n_1116),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.C1(n_150),
.C2(n_153),
.Y(n_1212)
);

AOI221xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1157),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.C(n_163),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1121),
.B(n_167),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1120),
.B(n_171),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1161),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1145),
.A2(n_175),
.B1(n_177),
.B2(n_180),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1165),
.A2(n_1139),
.B1(n_1130),
.B2(n_1142),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1171),
.A2(n_181),
.B(n_182),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1133),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1170),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1124),
.A2(n_189),
.B1(n_193),
.B2(n_194),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1163),
.A2(n_195),
.B1(n_197),
.B2(n_199),
.Y(n_1223)
);

NAND2x1_ASAP7_75t_L g1224 ( 
.A(n_1108),
.B(n_200),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1158),
.B(n_201),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1126),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_1226)
);

AOI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1144),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1154),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1135),
.Y(n_1229)
);

AOI32xp33_ASAP7_75t_L g1230 ( 
.A1(n_1112),
.A2(n_216),
.A3(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1159),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1108),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1114),
.B(n_227),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1128),
.B(n_1154),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1174),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1114),
.B(n_232),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1166),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1162),
.A2(n_237),
.B1(n_243),
.B2(n_244),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1173),
.A2(n_245),
.B(n_249),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1156),
.A2(n_250),
.B1(n_253),
.B2(n_255),
.C(n_257),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1220),
.B(n_1173),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1205),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1178),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1186),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1189),
.B(n_1160),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1189),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1234),
.B(n_1175),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1198),
.B(n_1175),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1232),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1190),
.B(n_1123),
.Y(n_1250)
);

NOR2x1_ASAP7_75t_L g1251 ( 
.A(n_1218),
.B(n_1172),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1200),
.B(n_1172),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1215),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1197),
.B(n_1177),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1213),
.A2(n_258),
.B(n_259),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_1183),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1211),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1179),
.B(n_260),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1228),
.B(n_261),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1229),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1203),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1176),
.B(n_263),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1180),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1225),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1181),
.B(n_264),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1214),
.B(n_267),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1213),
.B(n_268),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1227),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1207),
.B(n_269),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_270),
.Y(n_1270)
);

AO22x1_ASAP7_75t_L g1271 ( 
.A1(n_1183),
.A2(n_1233),
.B1(n_1185),
.B2(n_1196),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1188),
.B(n_1207),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1209),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1209),
.B(n_273),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1224),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1212),
.B(n_278),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1233),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1236),
.Y(n_1278)
);

OAI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1187),
.A2(n_279),
.B1(n_285),
.B2(n_286),
.C(n_287),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1237),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1212),
.B(n_288),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1195),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1235),
.B(n_289),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1191),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1219),
.Y(n_1285)
);

OAI211xp5_ASAP7_75t_L g1286 ( 
.A1(n_1193),
.A2(n_290),
.B(n_292),
.C(n_293),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1192),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1194),
.A2(n_294),
.B1(n_298),
.B2(n_299),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1239),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1276),
.A2(n_1199),
.B1(n_1202),
.B2(n_1206),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1276),
.A2(n_1238),
.B1(n_1208),
.B2(n_1201),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1243),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1290),
.B(n_1222),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1243),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1242),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1242),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1260),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1245),
.B(n_1221),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1244),
.B(n_1204),
.Y(n_1300)
);

NAND5xp2_ASAP7_75t_SL g1301 ( 
.A(n_1281),
.B(n_1210),
.C(n_1240),
.D(n_1231),
.E(n_1216),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1246),
.B(n_1245),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1247),
.B(n_1223),
.Y(n_1303)
);

AOI331xp33_ASAP7_75t_L g1304 ( 
.A1(n_1287),
.A2(n_1217),
.A3(n_1182),
.B1(n_1230),
.B2(n_303),
.B3(n_304),
.C1(n_305),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1246),
.B(n_300),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_R g1306 ( 
.A(n_1263),
.B(n_301),
.Y(n_1306)
);

OAI33xp33_ASAP7_75t_L g1307 ( 
.A1(n_1253),
.A2(n_302),
.A3(n_306),
.B1(n_307),
.B2(n_308),
.B3(n_310),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1247),
.Y(n_1308)
);

OAI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1287),
.A2(n_311),
.B1(n_312),
.B2(n_314),
.C(n_320),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1281),
.A2(n_324),
.B1(n_328),
.B2(n_330),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1279),
.A2(n_1259),
.B1(n_1280),
.B2(n_1283),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1259),
.A2(n_331),
.B1(n_333),
.B2(n_334),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1248),
.B(n_336),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1241),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1280),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1288),
.A2(n_341),
.B1(n_348),
.B2(n_354),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1241),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1241),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1283),
.A2(n_355),
.B1(n_356),
.B2(n_358),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1256),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1265),
.A2(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1257),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1257),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1249),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1297),
.B(n_1248),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1308),
.B(n_1253),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1317),
.B(n_1241),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_R g1328 ( 
.A(n_1306),
.B(n_1263),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1302),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1308),
.B(n_1278),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1302),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1317),
.B(n_1254),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1318),
.B(n_1254),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1318),
.B(n_1278),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1293),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1296),
.B(n_1252),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1314),
.B(n_1256),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1293),
.Y(n_1338)
);

NOR2x1_ASAP7_75t_L g1339 ( 
.A(n_1298),
.B(n_1251),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1314),
.B(n_1251),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1296),
.B(n_1282),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1295),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1311),
.B(n_1267),
.C(n_1262),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1295),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1322),
.B(n_1282),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1323),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1324),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1320),
.B(n_1261),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1348),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1335),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1348),
.B(n_1320),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1335),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1342),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1325),
.B(n_1299),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1342),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1327),
.B(n_1320),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1337),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1344),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1343),
.A2(n_1292),
.B1(n_1310),
.B2(n_1291),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1347),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1327),
.B(n_1320),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1344),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1360),
.B(n_1340),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1351),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1350),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1360),
.B(n_1354),
.Y(n_1366)
);

OAI31xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1359),
.A2(n_1339),
.A3(n_1300),
.B(n_1294),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1349),
.B(n_1340),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1351),
.B(n_1333),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1352),
.B(n_1329),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1357),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1357),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1349),
.B(n_1336),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1356),
.B(n_1298),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1353),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1355),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1358),
.B(n_1336),
.Y(n_1377)
);

OAI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1367),
.A2(n_1328),
.B1(n_1312),
.B2(n_1319),
.C(n_1262),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1367),
.A2(n_1326),
.B(n_1330),
.C(n_1346),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1371),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1364),
.A2(n_1303),
.B1(n_1299),
.B2(n_1356),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1365),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1369),
.Y(n_1385)
);

OAI21xp33_ASAP7_75t_L g1386 ( 
.A1(n_1366),
.A2(n_1303),
.B(n_1313),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1378),
.A2(n_1363),
.B1(n_1368),
.B2(n_1373),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1384),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1385),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1379),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1379),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1381),
.B(n_1377),
.Y(n_1392)
);

NOR3xp33_ASAP7_75t_SL g1393 ( 
.A(n_1387),
.B(n_1386),
.C(n_1309),
.Y(n_1393)
);

OAI211xp5_ASAP7_75t_L g1394 ( 
.A1(n_1390),
.A2(n_1380),
.B(n_1382),
.C(n_1383),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1391),
.B(n_1361),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1392),
.B(n_1389),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1388),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1390),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1394),
.A2(n_1301),
.B(n_1375),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1393),
.A2(n_1376),
.B(n_1370),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1398),
.Y(n_1401)
);

NOR3x1_ASAP7_75t_L g1402 ( 
.A(n_1396),
.B(n_1271),
.C(n_1258),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1398),
.B(n_1267),
.C(n_1321),
.Y(n_1403)
);

NOR3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1397),
.B(n_1266),
.C(n_1307),
.Y(n_1404)
);

NOR3xp33_ASAP7_75t_L g1405 ( 
.A(n_1395),
.B(n_1250),
.C(n_1270),
.Y(n_1405)
);

AOI322xp5_ASAP7_75t_L g1406 ( 
.A1(n_1400),
.A2(n_1272),
.A3(n_1313),
.B1(n_1370),
.B2(n_1333),
.C1(n_1332),
.C2(n_1331),
.Y(n_1406)
);

NAND4xp25_ASAP7_75t_SL g1407 ( 
.A(n_1399),
.B(n_1286),
.C(n_1332),
.D(n_1290),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1401),
.B(n_1362),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1403),
.B(n_1346),
.Y(n_1409)
);

OAI211xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1404),
.A2(n_1405),
.B(n_1402),
.C(n_1315),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1399),
.A2(n_1301),
.B1(n_1255),
.B2(n_1320),
.Y(n_1411)
);

AO22x2_ASAP7_75t_L g1412 ( 
.A1(n_1408),
.A2(n_1409),
.B1(n_1410),
.B2(n_1407),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1411),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1406),
.Y(n_1414)
);

OAI21xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1406),
.A2(n_1329),
.B(n_1331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1406),
.B(n_1334),
.Y(n_1416)
);

AOI321xp33_ASAP7_75t_L g1417 ( 
.A1(n_1407),
.A2(n_1304),
.A3(n_1289),
.B1(n_1316),
.B2(n_1274),
.C(n_1269),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1414),
.B(n_1334),
.Y(n_1418)
);

NOR2x1_ASAP7_75t_L g1419 ( 
.A(n_1413),
.B(n_1274),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1416),
.B(n_1269),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1412),
.B(n_1337),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1415),
.B(n_1338),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1417),
.B(n_1275),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1412),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_SL g1425 ( 
.A(n_1424),
.B(n_1418),
.C(n_1423),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1419),
.B(n_1337),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1421),
.B(n_1269),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1420),
.B(n_1341),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1422),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1424),
.A2(n_1305),
.B(n_1268),
.C(n_1284),
.Y(n_1430)
);

NOR3x1_ASAP7_75t_SL g1431 ( 
.A(n_1424),
.B(n_1271),
.C(n_1269),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1427),
.B(n_1305),
.Y(n_1432)
);

NAND4xp25_ASAP7_75t_L g1433 ( 
.A(n_1429),
.B(n_1274),
.C(n_1277),
.D(n_1272),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1425),
.B(n_1341),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1426),
.B(n_1345),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1428),
.Y(n_1436)
);

NAND4xp75_ASAP7_75t_L g1437 ( 
.A(n_1431),
.B(n_1255),
.C(n_1275),
.D(n_1284),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1430),
.B(n_1345),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_R g1439 ( 
.A1(n_1431),
.A2(n_1268),
.B1(n_1285),
.B2(n_1264),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1436),
.Y(n_1440)
);

AND4x1_ASAP7_75t_L g1441 ( 
.A(n_1434),
.B(n_1273),
.C(n_1274),
.D(n_1285),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1440),
.A2(n_1437),
.B1(n_1432),
.B2(n_1435),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1441),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1442),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1443),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1444),
.A2(n_1438),
.B(n_1439),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1445),
.B(n_1433),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_R g1448 ( 
.A(n_1447),
.B(n_364),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1448),
.A2(n_1446),
.B1(n_1277),
.B2(n_1255),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1449),
.A2(n_1273),
.B1(n_1256),
.B2(n_368),
.C(n_369),
.Y(n_1450)
);

AOI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1450),
.A2(n_366),
.B(n_367),
.C(n_370),
.Y(n_1451)
);


endmodule