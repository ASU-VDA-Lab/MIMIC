module fake_jpeg_12668_n_509 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_54),
.B(n_57),
.Y(n_145)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_16),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_81),
.Y(n_123)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_16),
.B(n_13),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_13),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_24),
.B(n_13),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_33),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_49),
.Y(n_139)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_33),
.B(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_40),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_22),
.C(n_41),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_41),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_131),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_22),
.B1(n_47),
.B2(n_46),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_118),
.A2(n_134),
.B1(n_136),
.B2(n_143),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_21),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_77),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_42),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_63),
.A2(n_22),
.B1(n_47),
.B2(n_46),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_64),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_45),
.B1(n_31),
.B2(n_41),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_75),
.B(n_23),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_53),
.A2(n_41),
.B1(n_21),
.B2(n_49),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_25),
.B1(n_29),
.B2(n_36),
.Y(n_195)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_20),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_29),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_160),
.B(n_203),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_188),
.Y(n_211)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_170),
.Y(n_214)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_108),
.A2(n_74),
.B1(n_84),
.B2(n_45),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_177),
.Y(n_226)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_175),
.A2(n_180),
.B1(n_190),
.B2(n_199),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_104),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

NOR2x1_ASAP7_75t_R g210 ( 
.A(n_178),
.B(n_87),
.Y(n_210)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_183),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_103),
.B(n_96),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_182),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_95),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_185),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_186),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_78),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_192),
.Y(n_213)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_116),
.A2(n_45),
.B1(n_49),
.B2(n_39),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_113),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_200),
.C(n_89),
.Y(n_220)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_44),
.B1(n_38),
.B2(n_25),
.Y(n_225)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_197),
.Y(n_245)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_120),
.B(n_122),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_201),
.Y(n_221)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_92),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_37),
.B1(n_20),
.B2(n_39),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_132),
.B1(n_44),
.B2(n_29),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_56),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_129),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_205),
.Y(n_231)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_115),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_138),
.B1(n_149),
.B2(n_135),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_174),
.B(n_162),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_209),
.A2(n_179),
.B(n_164),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_37),
.B(n_39),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_212),
.A2(n_38),
.B(n_18),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_160),
.B(n_117),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_216),
.B(n_218),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_163),
.B(n_182),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_141),
.A3(n_128),
.B1(n_117),
.B2(n_132),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_119),
.B1(n_86),
.B2(n_62),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_224),
.B1(n_140),
.B2(n_114),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_167),
.A2(n_119),
.B1(n_149),
.B2(n_135),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_38),
.B1(n_18),
.B2(n_25),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_158),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_157),
.C(n_68),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_72),
.C(n_142),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_142),
.C(n_69),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_128),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_193),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_211),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_258),
.C(n_265),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_224),
.B1(n_36),
.B2(n_18),
.Y(n_283)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_256),
.Y(n_304)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_266),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_226),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_169),
.B1(n_170),
.B2(n_166),
.Y(n_257)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_261),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_200),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_200),
.C(n_188),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_267),
.A2(n_276),
.B1(n_227),
.B2(n_180),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_213),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_214),
.Y(n_306)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_281),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_213),
.A2(n_194),
.B1(n_205),
.B2(n_171),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_274),
.B(n_230),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_159),
.B1(n_173),
.B2(n_196),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_222),
.A2(n_199),
.B1(n_184),
.B2(n_197),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_221),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_283),
.A2(n_312),
.B1(n_183),
.B2(n_191),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_246),
.A2(n_215),
.B1(n_207),
.B2(n_216),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_284),
.A2(n_302),
.B1(n_309),
.B2(n_278),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_287),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_262),
.B(n_277),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_211),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_280),
.B1(n_281),
.B2(n_259),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_249),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_292),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_242),
.B(n_232),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_245),
.B(n_236),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_223),
.B1(n_210),
.B2(n_234),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_310),
.B(n_311),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_242),
.B1(n_239),
.B2(n_211),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_223),
.CI(n_229),
.CON(n_303),
.SN(n_303)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_303),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_255),
.Y(n_332)
);

OAI22x1_ASAP7_75t_SL g309 ( 
.A1(n_254),
.A2(n_219),
.B1(n_225),
.B2(n_214),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_248),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_260),
.A2(n_220),
.B1(n_241),
.B2(n_217),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_236),
.B1(n_245),
.B2(n_227),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_250),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g334 ( 
.A1(n_315),
.A2(n_273),
.B(n_264),
.Y(n_334)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_321),
.B1(n_329),
.B2(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_279),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_340),
.Y(n_362)
);

AO22x1_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_257),
.B1(n_254),
.B2(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_271),
.B1(n_265),
.B2(n_247),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_333),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_258),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_335),
.C(n_343),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_314),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_266),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_290),
.A2(n_254),
.B1(n_263),
.B2(n_267),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_338),
.B1(n_285),
.B2(n_286),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_294),
.B(n_284),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_331),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_257),
.B1(n_254),
.B2(n_261),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_274),
.B1(n_253),
.B2(n_245),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_342),
.B1(n_282),
.B2(n_290),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_314),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_237),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_300),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_238),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_347),
.C(n_349),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_295),
.B1(n_121),
.B2(n_125),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_243),
.C(n_238),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_302),
.B(n_238),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_356),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_354),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_363),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_291),
.B1(n_301),
.B2(n_282),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_301),
.B1(n_282),
.B2(n_288),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_359),
.A2(n_360),
.B1(n_367),
.B2(n_371),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_292),
.B1(n_306),
.B2(n_308),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_304),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_303),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_377),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_318),
.A2(n_286),
.B1(n_298),
.B2(n_312),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_308),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_338),
.A2(n_314),
.B(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_372),
.B(n_375),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_303),
.C(n_297),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_358),
.C(n_355),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_315),
.B1(n_310),
.B2(n_313),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_313),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_313),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_238),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_283),
.B1(n_295),
.B2(n_227),
.Y(n_379)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_393),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_345),
.C(n_349),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_386),
.C(n_395),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_366),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_404),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_324),
.C(n_326),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_324),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_391),
.B(n_396),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_327),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_377),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_400),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_316),
.C(n_341),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_362),
.B(n_327),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_341),
.C(n_238),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_401),
.C(n_402),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_319),
.C(n_161),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_319),
.C(n_175),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_299),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_299),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_409),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_121),
.C(n_125),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_375),
.C(n_381),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_299),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_398),
.A2(n_367),
.B1(n_369),
.B2(n_380),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_411),
.A2(n_422),
.B1(n_429),
.B2(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_372),
.B(n_359),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_414),
.A2(n_427),
.B(n_431),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_360),
.B1(n_356),
.B2(n_352),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_34),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_398),
.A2(n_368),
.B1(n_353),
.B2(n_364),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_374),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_424),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_361),
.C(n_140),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_428),
.C(n_430),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_60),
.C(n_99),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_59),
.C(n_80),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_390),
.A2(n_37),
.B(n_44),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_432),
.A2(n_26),
.B1(n_23),
.B2(n_2),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_382),
.C(n_386),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_450),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_416),
.A2(n_397),
.B1(n_395),
.B2(n_406),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_435),
.A2(n_437),
.B1(n_443),
.B2(n_444),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_416),
.A2(n_389),
.B1(n_399),
.B2(n_394),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_399),
.Y(n_439)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_441),
.Y(n_456)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_440),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_413),
.B(n_400),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_421),
.A2(n_66),
.B1(n_71),
.B2(n_36),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_423),
.A2(n_206),
.B1(n_34),
.B2(n_2),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_422),
.A2(n_206),
.B1(n_26),
.B2(n_23),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_447),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_34),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_426),
.C(n_410),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_449),
.B(n_418),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_417),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_462),
.Y(n_473)
);

BUFx4f_ASAP7_75t_SL g454 ( 
.A(n_438),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_457),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_436),
.A2(n_423),
.B1(n_411),
.B2(n_431),
.Y(n_459)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_419),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_461),
.B(n_5),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_451),
.A2(n_430),
.B(n_428),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_435),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_466),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_0),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_34),
.C(n_26),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_26),
.C(n_3),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_26),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_442),
.C(n_441),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_442),
.C(n_446),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_443),
.C(n_433),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_475),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_455),
.A2(n_444),
.B(n_3),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_477),
.B(n_6),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_0),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_482),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_460),
.A2(n_0),
.B(n_3),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_0),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_465),
.C(n_459),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_469),
.B(n_454),
.Y(n_484)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_473),
.C(n_454),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_486),
.A2(n_477),
.B(n_492),
.Y(n_497)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_488),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_478),
.C(n_475),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_468),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_490),
.A2(n_491),
.B(n_480),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_470),
.A2(n_467),
.B(n_466),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_494),
.A2(n_496),
.B(n_483),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_SL g501 ( 
.A1(n_497),
.A2(n_498),
.B(n_485),
.C(n_7),
.Y(n_501)
);

AOI321xp33_ASAP7_75t_SL g498 ( 
.A1(n_486),
.A2(n_456),
.A3(n_479),
.B1(n_476),
.B2(n_9),
.C(n_6),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_500),
.A2(n_501),
.B(n_502),
.Y(n_505)
);

O2A1O1Ixp33_ASAP7_75t_SL g502 ( 
.A1(n_498),
.A2(n_490),
.B(n_7),
.C(n_8),
.Y(n_502)
);

OAI321xp33_ASAP7_75t_L g503 ( 
.A1(n_493),
.A2(n_495),
.A3(n_499),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_6),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_6),
.B(n_7),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_505),
.B(n_9),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_10),
.C(n_497),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_10),
.Y(n_509)
);


endmodule