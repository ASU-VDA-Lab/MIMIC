module fake_jpeg_6663_n_306 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_286;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_38),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_6),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_40),
.A2(n_45),
.B(n_20),
.C(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_43),
.B(n_23),
.Y(n_94)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_52),
.Y(n_108)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_92),
.B1(n_23),
.B2(n_25),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_57),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_58),
.B(n_76),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_86),
.B1(n_91),
.B2(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_24),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_16),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_87),
.B(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_36),
.A2(n_34),
.B1(n_19),
.B2(n_16),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_19),
.B1(n_31),
.B2(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_90),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_40),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_127),
.B1(n_83),
.B2(n_18),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_20),
.B1(n_18),
.B2(n_15),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_15),
.B1(n_32),
.B2(n_14),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_123),
.B1(n_110),
.B2(n_99),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_28),
.B1(n_31),
.B2(n_18),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_31),
.B1(n_18),
.B2(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_128),
.B(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_55),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_131),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_59),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_137),
.Y(n_175)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_60),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_51),
.B1(n_96),
.B2(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_138),
.B(n_139),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_98),
.B1(n_90),
.B2(n_63),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_60),
.C(n_71),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_118),
.B(n_107),
.Y(n_192)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_156),
.B1(n_162),
.B2(n_101),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_66),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

OAI22x1_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_93),
.B1(n_95),
.B2(n_77),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_157),
.B(n_159),
.Y(n_191)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_32),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_10),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_114),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_121),
.B(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_32),
.B(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_32),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_126),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_15),
.B1(n_32),
.B2(n_14),
.Y(n_162)
);

NOR4xp25_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_137),
.C(n_131),
.D(n_144),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_152),
.B(n_149),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_127),
.B1(n_73),
.B2(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_174),
.B1(n_163),
.B2(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_189),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_124),
.B(n_111),
.C(n_107),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_171),
.A2(n_172),
.B(n_5),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_157),
.B(n_159),
.Y(n_172)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_125),
.B1(n_14),
.B2(n_122),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_187),
.B1(n_140),
.B2(n_136),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_122),
.B1(n_118),
.B2(n_126),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_9),
.C(n_12),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_1),
.C(n_2),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_130),
.B(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_10),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_199),
.CI(n_201),
.CON(n_231),
.SN(n_231)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_160),
.B(n_133),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_204),
.B1(n_206),
.B2(n_166),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_139),
.B(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_203),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_179),
.B1(n_185),
.B2(n_166),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_8),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_1),
.C(n_2),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_1),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_3),
.B(n_4),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_8),
.Y(n_215)
);

OAI322xp33_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_173),
.A3(n_182),
.B1(n_184),
.B2(n_178),
.C1(n_174),
.C2(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_3),
.B(n_4),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_220),
.B1(n_181),
.B2(n_9),
.C(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

HAxp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_221),
.CON(n_229),
.SN(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

AO32x1_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_174),
.A3(n_166),
.B1(n_171),
.B2(n_177),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_238),
.B(n_219),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_207),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_196),
.B1(n_222),
.B2(n_169),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_195),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_217),
.B(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_197),
.C(n_199),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_251),
.C(n_258),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_225),
.A2(n_241),
.B1(n_212),
.B2(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_225),
.B1(n_222),
.B2(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_235),
.C(n_201),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_259),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_195),
.C(n_209),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_223),
.C(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_231),
.C(n_228),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_229),
.B1(n_214),
.B2(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_269),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_246),
.B(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_243),
.C(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_246),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_276),
.B(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_169),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_242),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_283),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_249),
.C(n_244),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_264),
.A3(n_257),
.B1(n_261),
.B2(n_263),
.C1(n_260),
.C2(n_259),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_279),
.C(n_278),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_196),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_236),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_262),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_290),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_260),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_186),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_293),
.B(n_289),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_254),
.B(n_193),
.C(n_285),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_279),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_298),
.B(n_288),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_300),
.B(n_302),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_230),
.B1(n_234),
.B2(n_226),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_295),
.A3(n_254),
.B1(n_232),
.B2(n_185),
.C1(n_253),
.C2(n_164),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_256),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_304),
.Y(n_306)
);


endmodule