module fake_jpeg_25320_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_27),
.B1(n_22),
.B2(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_16),
.B1(n_10),
.B2(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_9),
.C(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_28),
.B1(n_9),
.B2(n_31),
.Y(n_50)
);

NOR2x1p5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_15),
.Y(n_41)
);

NAND2x1p5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_15),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_8),
.C(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_39),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_51),
.B1(n_41),
.B2(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_59),
.C(n_60),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_41),
.B(n_31),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_47),
.B1(n_38),
.B2(n_42),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_46),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_51),
.B(n_53),
.C(n_50),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_55),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_43),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_59),
.CI(n_43),
.CON(n_67),
.SN(n_67)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_62),
.A3(n_61),
.B1(n_64),
.B2(n_42),
.C(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_3),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_70),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_67),
.B1(n_66),
.B2(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_71),
.B1(n_3),
.B2(n_5),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_5),
.Y(n_74)
);


endmodule