module fake_jpeg_31753_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_25),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_42),
.B(n_9),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_22),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_40),
.B1(n_9),
.B2(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_26),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_25),
.B1(n_14),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_75),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_82),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_14),
.B1(n_29),
.B2(n_24),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_40),
.C(n_38),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_74),
.C(n_53),
.Y(n_87)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

XOR2x2_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_13),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_41),
.B1(n_16),
.B2(n_21),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_13),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_21),
.B1(n_29),
.B2(n_13),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_11),
.B1(n_13),
.B2(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_50),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_93),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_48),
.B(n_61),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_99),
.B(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_61),
.Y(n_95)
);

AND2x4_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_54),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_71),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_72),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.C(n_109),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_77),
.C(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_86),
.B1(n_90),
.B2(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_92),
.B1(n_91),
.B2(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_96),
.B(n_99),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_96),
.B(n_88),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_105),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_125),
.C(n_127),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_109),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_91),
.C(n_102),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_103),
.C(n_84),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_114),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_119),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_129),
.B1(n_132),
.B2(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_134),
.B1(n_132),
.B2(n_135),
.C(n_54),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_69),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_84),
.Y(n_143)
);


endmodule