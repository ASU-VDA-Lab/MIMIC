module fake_netlist_6_3482_n_1754 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1754);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1754;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_76),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_23),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_22),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_52),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_0),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_37),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_44),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_47),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_81),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_45),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_20),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_112),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_67),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_2),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_57),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_24),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_96),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_27),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_48),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_50),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_46),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_57),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_32),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_29),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_77),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_25),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_92),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_13),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_31),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_116),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_45),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_73),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_24),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_119),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_22),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_93),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_0),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_16),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_99),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_100),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_65),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_71),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_7),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_90),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_41),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_26),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_140),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_6),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_65),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_86),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_130),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_155),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_126),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_87),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_61),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_70),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_5),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_79),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_143),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_115),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_98),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_63),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_134),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_54),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_15),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_78),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_23),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_62),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_137),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_72),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_53),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_1),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_19),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_56),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_103),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_41),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_153),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_39),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_1),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_26),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_192),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_161),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_195),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_192),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_192),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_184),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_192),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_192),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_199),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_171),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_3),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_192),
.B(n_4),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_191),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_252),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_192),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_202),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_175),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_283),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_4),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_169),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_175),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_167),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_205),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_167),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_167),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_222),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_167),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_211),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_218),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_227),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_232),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_209),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_244),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_177),
.B(n_8),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_209),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_209),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_178),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_173),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_255),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_258),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_177),
.B(n_9),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_249),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_264),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_273),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_156),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_193),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_173),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_196),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_156),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_197),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_200),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_208),
.B(n_9),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_203),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_157),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_279),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_157),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_160),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_210),
.B(n_10),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_249),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_279),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_189),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_214),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_208),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_210),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_323),
.B(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_226),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_331),
.B(n_217),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_358),
.A2(n_261),
.B(n_226),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_376),
.B(n_181),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_316),
.B(n_261),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_318),
.B(n_284),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_186),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_318),
.B(n_284),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_357),
.B(n_217),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_193),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_319),
.B(n_322),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_369),
.B(n_277),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_367),
.B(n_277),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_350),
.B(n_159),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_324),
.B(n_224),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

OA21x2_ASAP7_75t_L g435 ( 
.A1(n_324),
.A2(n_198),
.B(n_194),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_353),
.B(n_354),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_224),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_354),
.Y(n_438)
);

BUFx8_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_163),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_364),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_404),
.A2(n_339),
.B1(n_225),
.B2(n_295),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_404),
.B(n_413),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_314),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_391),
.B(n_224),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_399),
.B(n_320),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_328),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_415),
.A2(n_344),
.B1(n_235),
.B2(n_201),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_412),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_391),
.B(n_406),
.Y(n_457)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_289),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_404),
.B(n_380),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_415),
.B(n_224),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_390),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_332),
.Y(n_464)
);

INVx8_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_352),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_387),
.A2(n_204),
.B1(n_254),
.B2(n_253),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_398),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_429),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_436),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g474 ( 
.A1(n_406),
.A2(n_313),
.B1(n_325),
.B2(n_317),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_429),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_387),
.A2(n_355),
.B1(n_346),
.B2(n_348),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_401),
.A2(n_341),
.B1(n_356),
.B2(n_374),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_401),
.B(n_326),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_311),
.C(n_335),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_R g483 ( 
.A(n_442),
.B(n_342),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_361),
.B1(n_375),
.B2(n_372),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_391),
.B(n_224),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

AND3x2_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_248),
.C(n_180),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_423),
.B(n_343),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_442),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_359),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_384),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_435),
.A2(n_259),
.B1(n_213),
.B2(n_309),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_373),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_427),
.A2(n_366),
.B1(n_360),
.B2(n_330),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_441),
.B(n_373),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_378),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_422),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_435),
.A2(n_256),
.B1(n_228),
.B2(n_303),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_420),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_379),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_428),
.B(n_176),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_441),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_410),
.B(n_229),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_385),
.B(n_310),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_428),
.B(n_188),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_410),
.B(n_229),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_385),
.B(n_160),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_410),
.B(n_229),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_389),
.Y(n_529)
);

AO22x2_ASAP7_75t_L g530 ( 
.A1(n_410),
.A2(n_207),
.B1(n_242),
.B2(n_281),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_435),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_393),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_393),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_393),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_229),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_383),
.B(n_206),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_439),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_422),
.A2(n_246),
.B1(n_269),
.B2(n_266),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_430),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_439),
.B(n_229),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_382),
.B(n_378),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_383),
.B(n_212),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_439),
.B(n_294),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_439),
.B(n_294),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_437),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_439),
.B(n_294),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_394),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_439),
.B(n_294),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_383),
.B(n_215),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_438),
.B(n_162),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_394),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_382),
.B(n_294),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_431),
.A2(n_297),
.B1(n_282),
.B2(n_267),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_424),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_383),
.B(n_220),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_438),
.B(n_162),
.Y(n_571)
);

AND2x2_ASAP7_75t_SL g572 ( 
.A(n_431),
.B(n_297),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_430),
.A2(n_304),
.B1(n_301),
.B2(n_292),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_424),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_382),
.B(n_297),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_389),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_381),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_438),
.B(n_164),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_411),
.B(n_245),
.C(n_216),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_381),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_440),
.B(n_164),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_381),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_388),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_388),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_425),
.B(n_297),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_388),
.B(n_233),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_392),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_440),
.B(n_277),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_402),
.A2(n_297),
.B1(n_237),
.B2(n_262),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_392),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_440),
.B(n_165),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_511),
.B(n_425),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_500),
.B(n_165),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_510),
.B(n_250),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_520),
.B(n_443),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_479),
.B(n_243),
.C(n_241),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_425),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_447),
.A2(n_179),
.B1(n_182),
.B2(n_301),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_447),
.A2(n_179),
.B1(n_182),
.B2(n_292),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_580),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_465),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_448),
.B(n_185),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_497),
.B(n_185),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_514),
.B(n_190),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_514),
.B(n_190),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_425),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_580),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_465),
.B(n_425),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_543),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_452),
.B(n_238),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_465),
.B(n_260),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_446),
.C(n_460),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_501),
.A2(n_414),
.B1(n_411),
.B2(n_268),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_453),
.B(n_238),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_SL g616 ( 
.A(n_486),
.B(n_166),
.C(n_168),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_449),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_582),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_582),
.Y(n_619)
);

NOR2x1_ASAP7_75t_L g620 ( 
.A(n_481),
.B(n_579),
.Y(n_620)
);

BUFx8_ASAP7_75t_L g621 ( 
.A(n_463),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_531),
.A2(n_286),
.B1(n_304),
.B2(n_276),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_472),
.B(n_425),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_585),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_460),
.B(n_286),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_472),
.B(n_425),
.Y(n_626)
);

NAND2x1p5_ASAP7_75t_L g627 ( 
.A(n_501),
.B(n_403),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_457),
.B(n_270),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_517),
.A2(n_414),
.B1(n_411),
.B2(n_272),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_517),
.A2(n_414),
.B1(n_274),
.B2(n_271),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_472),
.B(n_426),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_522),
.B(n_554),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_490),
.B(n_426),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_496),
.B(n_219),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_490),
.B(n_426),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_589),
.B(n_402),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_459),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_531),
.A2(n_402),
.B1(n_426),
.B2(n_249),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_590),
.B(n_249),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_426),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_572),
.B(n_426),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_496),
.B(n_221),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_572),
.B(n_426),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_544),
.B(n_443),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_463),
.B(n_223),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_504),
.B(n_443),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_552),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_469),
.B(n_230),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_589),
.B(n_527),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_566),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_588),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_467),
.B(n_426),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_469),
.B(n_231),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_591),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_473),
.B(n_426),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_477),
.B(n_402),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_483),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_503),
.B(n_249),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_553),
.B(n_426),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_389),
.Y(n_664)
);

BUFx8_ASAP7_75t_L g665 ( 
.A(n_504),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_591),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_455),
.B(n_240),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_509),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_577),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_456),
.B(n_471),
.Y(n_670)
);

OAI221xp5_ASAP7_75t_L g671 ( 
.A1(n_454),
.A2(n_251),
.B1(n_257),
.B2(n_263),
.C(n_265),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_461),
.B(n_389),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_461),
.B(n_389),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_583),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_482),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_509),
.B(n_444),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_499),
.B(n_464),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_547),
.B(n_444),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_547),
.B(n_516),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_482),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_389),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_464),
.B(n_166),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_516),
.B(n_389),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_516),
.B(n_408),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_505),
.B(n_402),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_488),
.A2(n_392),
.B(n_400),
.C(n_434),
.Y(n_686)
);

BUFx8_ASAP7_75t_L g687 ( 
.A(n_510),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_510),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_492),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_506),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_512),
.B(n_408),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_488),
.B(n_444),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_458),
.A2(n_402),
.B1(n_249),
.B2(n_434),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_573),
.B(n_402),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_515),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_530),
.B(n_403),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_508),
.B(n_408),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_515),
.A2(n_395),
.B1(n_405),
.B2(n_434),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_566),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_464),
.B(n_168),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_530),
.B(n_444),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_464),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_515),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_466),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_492),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_530),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_530),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_524),
.B(n_408),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_466),
.B(n_170),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_560),
.B(n_249),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_466),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_494),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_494),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_450),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_466),
.B(n_444),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_408),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_578),
.B(n_249),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_581),
.B(n_408),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_408),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_451),
.B(n_408),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_450),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_540),
.B(n_170),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_540),
.B(n_172),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_541),
.B(n_172),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_518),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_475),
.B(n_174),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_451),
.B(n_408),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_518),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_451),
.B(n_408),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_462),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_462),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_458),
.A2(n_416),
.B1(n_400),
.B2(n_395),
.Y(n_733)
);

AOI221xp5_ASAP7_75t_L g734 ( 
.A1(n_480),
.A2(n_305),
.B1(n_183),
.B2(n_187),
.C(n_236),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_470),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_451),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_475),
.B(n_174),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_532),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_458),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_451),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_458),
.A2(n_416),
.B1(n_400),
.B2(n_395),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_566),
.B(n_444),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_451),
.B(n_407),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_584),
.B(n_407),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_532),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_474),
.B(n_183),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_523),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_470),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_584),
.B(n_407),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_476),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_584),
.B(n_407),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_537),
.B(n_187),
.Y(n_752)
);

BUFx6f_ASAP7_75t_SL g753 ( 
.A(n_521),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_533),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_533),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_534),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_534),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_491),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_587),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_545),
.A2(n_396),
.B1(n_397),
.B2(n_405),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_476),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_548),
.B(n_407),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_559),
.B(n_305),
.C(n_239),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_688),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_601),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_653),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_679),
.B(n_523),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_593),
.A2(n_485),
.B(n_529),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_642),
.A2(n_570),
.B(n_525),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_645),
.A2(n_519),
.B(n_549),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_607),
.A2(n_529),
.B(n_485),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_609),
.A2(n_529),
.B(n_485),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_602),
.A2(n_558),
.B(n_545),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_567),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_610),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_691),
.A2(n_549),
.B(n_550),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_602),
.A2(n_626),
.B(n_623),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_631),
.A2(n_550),
.B(n_556),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_632),
.B(n_568),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_605),
.B(n_574),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_L g781 ( 
.A1(n_647),
.A2(n_288),
.B(n_291),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_633),
.A2(n_556),
.B(n_558),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_635),
.A2(n_564),
.B(n_575),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_653),
.B(n_523),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_641),
.A2(n_564),
.B(n_575),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_613),
.A2(n_651),
.B(n_628),
.C(n_707),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_759),
.B(n_535),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_617),
.A2(n_638),
.B(n_678),
.C(n_707),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_606),
.B(n_535),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_630),
.A2(n_546),
.B1(n_565),
.B2(n_478),
.Y(n_790)
);

CKINVDCx8_ASAP7_75t_R g791 ( 
.A(n_661),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_681),
.A2(n_495),
.B(n_493),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_678),
.B(n_538),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_688),
.A2(n_546),
.B1(n_487),
.B2(n_484),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_746),
.B(n_538),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_683),
.A2(n_498),
.B(n_489),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_616),
.B(n_291),
.C(n_236),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_708),
.A2(n_403),
.B(n_239),
.C(n_275),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_601),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_746),
.B(n_557),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_684),
.A2(n_502),
.B(n_576),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_596),
.B(n_648),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_661),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_670),
.B(n_275),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_708),
.A2(n_403),
.B(n_290),
.C(n_308),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_608),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_608),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_717),
.A2(n_507),
.B(n_576),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_614),
.A2(n_569),
.B1(n_563),
.B2(n_562),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_618),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_687),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_627),
.A2(n_562),
.B(n_569),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_596),
.B(n_278),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_648),
.B(n_557),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_594),
.A2(n_563),
.B(n_405),
.C(n_397),
.Y(n_816)
);

AO21x1_ASAP7_75t_L g817 ( 
.A1(n_685),
.A2(n_421),
.B(n_397),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_676),
.B(n_669),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_620),
.A2(n_521),
.B1(n_528),
.B2(n_526),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_719),
.A2(n_576),
.B(n_507),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_627),
.A2(n_521),
.B(n_526),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_720),
.A2(n_576),
.B(n_507),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_695),
.B(n_539),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_676),
.B(n_539),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_716),
.A2(n_521),
.B1(n_528),
.B2(n_526),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_669),
.B(n_555),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_629),
.A2(n_555),
.B1(n_396),
.B2(n_409),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_762),
.A2(n_598),
.B(n_652),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_627),
.A2(n_528),
.B(n_521),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_652),
.A2(n_576),
.B(n_507),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_652),
.A2(n_507),
.B(n_418),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_742),
.A2(n_407),
.B(n_418),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_674),
.B(n_555),
.Y(n_833)
);

BUFx12f_ASAP7_75t_L g834 ( 
.A(n_665),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_742),
.A2(n_418),
.B(n_555),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_664),
.A2(n_418),
.B(n_409),
.Y(n_836)
);

O2A1O1Ixp5_ASAP7_75t_L g837 ( 
.A1(n_694),
.A2(n_421),
.B(n_409),
.C(n_416),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_747),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_747),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_618),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_644),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_656),
.A2(n_418),
.B(n_417),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_649),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_649),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_619),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_687),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_659),
.A2(n_528),
.B(n_526),
.Y(n_847)
);

NOR2x1_ASAP7_75t_L g848 ( 
.A(n_763),
.B(n_396),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_677),
.B(n_278),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_536),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_695),
.B(n_418),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_646),
.B(n_536),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_699),
.A2(n_417),
.B(n_419),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_634),
.B(n_280),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_699),
.A2(n_417),
.B(n_419),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_704),
.B(n_433),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_646),
.B(n_536),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_L g858 ( 
.A(n_668),
.B(n_280),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_739),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_699),
.A2(n_419),
.B(n_421),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_650),
.B(n_657),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_599),
.B(n_144),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_704),
.A2(n_445),
.B(n_433),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_595),
.B(n_536),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_716),
.A2(n_528),
.B1(n_526),
.B2(n_521),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_663),
.A2(n_445),
.B(n_433),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_595),
.B(n_536),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_727),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_758),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_696),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_692),
.B(n_433),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_739),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_721),
.A2(n_445),
.B(n_433),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_728),
.A2(n_445),
.B(n_433),
.Y(n_874)
);

CKINVDCx10_ASAP7_75t_R g875 ( 
.A(n_665),
.Y(n_875)
);

BUFx2_ASAP7_75t_SL g876 ( 
.A(n_753),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_433),
.B(n_528),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_744),
.A2(n_433),
.B(n_526),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_692),
.B(n_433),
.Y(n_879)
);

NOR2x1_ASAP7_75t_L g880 ( 
.A(n_660),
.B(n_433),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_595),
.B(n_536),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_687),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_749),
.A2(n_586),
.B(n_308),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_702),
.B(n_148),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_747),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_665),
.B(n_298),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_751),
.A2(n_586),
.B(n_306),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_690),
.B(n_586),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_737),
.Y(n_889)
);

AOI21xp33_ASAP7_75t_L g890 ( 
.A1(n_622),
.A2(n_306),
.B(n_302),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_690),
.B(n_703),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_698),
.A2(n_586),
.B(n_302),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_639),
.A2(n_586),
.B(n_300),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_703),
.B(n_586),
.Y(n_894)
);

O2A1O1Ixp5_ASAP7_75t_L g895 ( 
.A1(n_636),
.A2(n_129),
.B(n_88),
.C(n_94),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_672),
.A2(n_132),
.B(n_97),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_752),
.B(n_300),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_725),
.A2(n_299),
.B(n_298),
.C(n_296),
.Y(n_898)
);

BUFx5_ASAP7_75t_L g899 ( 
.A(n_715),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_643),
.B(n_299),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_619),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_752),
.B(n_296),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_736),
.B(n_138),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_701),
.B(n_290),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_701),
.B(n_288),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_736),
.A2(n_285),
.B(n_127),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_673),
.B(n_285),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_624),
.B(n_11),
.Y(n_908)
);

AOI21xp33_ASAP7_75t_L g909 ( 
.A1(n_625),
.A2(n_11),
.B(n_12),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_740),
.A2(n_125),
.B(n_122),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_696),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_667),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_624),
.B(n_14),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_640),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_740),
.A2(n_118),
.B(n_113),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_662),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_734),
.A2(n_18),
.B(n_21),
.C(n_27),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_743),
.A2(n_709),
.B(n_697),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_758),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_637),
.B(n_654),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_637),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_712),
.B(n_28),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_654),
.A2(n_80),
.B(n_30),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_655),
.B(n_28),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_655),
.A2(n_33),
.B(n_34),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_658),
.B(n_33),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_705),
.B(n_34),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_658),
.A2(n_35),
.B(n_36),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_666),
.B(n_35),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_666),
.A2(n_36),
.B(n_37),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_38),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_711),
.A2(n_38),
.B(n_39),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_600),
.B(n_40),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_718),
.A2(n_42),
.B(n_43),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_682),
.B(n_42),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_662),
.A2(n_51),
.B(n_52),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_700),
.B(n_53),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_715),
.A2(n_54),
.B(n_55),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_611),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_675),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_612),
.A2(n_58),
.B(n_59),
.Y(n_941)
);

O2A1O1Ixp5_ASAP7_75t_L g942 ( 
.A1(n_604),
.A2(n_59),
.B(n_60),
.C(n_64),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_733),
.B(n_64),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_741),
.B(n_66),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_675),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_761),
.B(n_66),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_803),
.B(n_791),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_802),
.B(n_732),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_861),
.B(n_615),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_777),
.A2(n_748),
.B(n_735),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_916),
.A2(n_696),
.B1(n_760),
.B2(n_739),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_814),
.B(n_710),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_870),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_854),
.A2(n_597),
.B1(n_739),
.B2(n_723),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_766),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_870),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_780),
.B(n_724),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_854),
.B(n_696),
.Y(n_958)
);

NOR2x1_ASAP7_75t_L g959 ( 
.A(n_872),
.B(n_612),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_935),
.A2(n_671),
.B(n_640),
.C(n_686),
.Y(n_960)
);

INVxp33_ASAP7_75t_SL g961 ( 
.A(n_886),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_869),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_766),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_780),
.B(n_732),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_919),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_788),
.A2(n_693),
.B(n_750),
.C(n_748),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_788),
.A2(n_731),
.B(n_750),
.C(n_735),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_SL g968 ( 
.A1(n_916),
.A2(n_937),
.B1(n_935),
.B2(n_912),
.Y(n_968)
);

INVx3_ASAP7_75t_SL g969 ( 
.A(n_927),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_872),
.B(n_612),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_834),
.B(n_612),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_900),
.B(n_731),
.Y(n_972)
);

NOR2xp67_ASAP7_75t_SL g973 ( 
.A(n_876),
.B(n_753),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_868),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_775),
.Y(n_975)
);

AO21x1_ASAP7_75t_L g976 ( 
.A1(n_937),
.A2(n_722),
.B(n_680),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_900),
.B(n_804),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_786),
.A2(n_738),
.B(n_680),
.C(n_689),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_870),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_795),
.A2(n_738),
.B(n_689),
.C(n_706),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_795),
.B(n_745),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_828),
.A2(n_760),
.B(n_706),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_818),
.A2(n_760),
.B1(n_753),
.B2(n_714),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_884),
.B(n_745),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_813),
.A2(n_760),
.B(n_713),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_897),
.B(n_729),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_870),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_902),
.B(n_729),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_773),
.A2(n_754),
.B(n_713),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_800),
.B(n_714),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_800),
.B(n_787),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_812),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_927),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_889),
.A2(n_621),
.B1(n_726),
.B2(n_754),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_849),
.B(n_621),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_875),
.Y(n_996)
);

CKINVDCx16_ASAP7_75t_R g997 ( 
.A(n_846),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_806),
.B(n_726),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_922),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_764),
.B(n_621),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_781),
.B(n_797),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_824),
.A2(n_755),
.B(n_756),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_771),
.A2(n_755),
.B(n_756),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_905),
.B(n_904),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_890),
.B(n_757),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_841),
.A2(n_757),
.B1(n_844),
.B2(n_843),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_921),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_943),
.A2(n_944),
.B1(n_891),
.B2(n_911),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_789),
.A2(n_779),
.B(n_898),
.C(n_776),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_859),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_922),
.A2(n_917),
.B(n_939),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_882),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_764),
.B(n_838),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_779),
.B(n_904),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_768),
.A2(n_782),
.B(n_778),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_808),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_884),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_808),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_838),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_L g1020 ( 
.A(n_903),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_943),
.A2(n_944),
.B1(n_911),
.B2(n_907),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_789),
.A2(n_933),
.B(n_909),
.C(n_938),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_811),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_774),
.B(n_815),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_SL g1025 ( 
.A1(n_903),
.A2(n_893),
.B1(n_892),
.B2(n_917),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_858),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_907),
.B(n_848),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_772),
.A2(n_829),
.B(n_821),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_862),
.B(n_765),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_914),
.B(n_936),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_931),
.A2(n_946),
.B(n_942),
.C(n_929),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_769),
.A2(n_918),
.B(n_793),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_811),
.B(n_901),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_901),
.B(n_899),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_799),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_852),
.B(n_857),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_807),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_908),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_SL g1039 ( 
.A1(n_770),
.A2(n_906),
.B(n_847),
.C(n_783),
.Y(n_1039)
);

AO22x1_ASAP7_75t_L g1040 ( 
.A1(n_880),
.A2(n_864),
.B1(n_881),
.B2(n_867),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_840),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_767),
.A2(n_871),
.B1(n_879),
.B2(n_850),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_767),
.A2(n_871),
.B1(n_879),
.B2(n_851),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_798),
.A2(n_805),
.B1(n_826),
.B2(n_833),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_784),
.A2(n_835),
.B(n_790),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_845),
.B(n_945),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_823),
.B(n_839),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_913),
.A2(n_924),
.B1(n_926),
.B2(n_941),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_895),
.A2(n_792),
.B(n_796),
.C(n_832),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_798),
.A2(n_805),
.B(n_934),
.C(n_932),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_851),
.A2(n_940),
.B1(n_817),
.B2(n_899),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_784),
.A2(n_785),
.B(n_823),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_856),
.A2(n_801),
.B(n_809),
.Y(n_1053)
);

OAI22x1_ASAP7_75t_L g1054 ( 
.A1(n_819),
.A2(n_825),
.B1(n_865),
.B2(n_856),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_940),
.B(n_839),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_920),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_SL g1057 ( 
.A(n_925),
.B(n_930),
.C(n_928),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_923),
.A2(n_860),
.B(n_855),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_820),
.A2(n_822),
.B(n_794),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_899),
.B(n_885),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_899),
.B(n_885),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_899),
.A2(n_894),
.B1(n_888),
.B2(n_883),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_910),
.B(n_915),
.C(n_887),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_L g1064 ( 
.A(n_896),
.B(n_836),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_899),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_810),
.A2(n_827),
.B1(n_842),
.B2(n_853),
.Y(n_1066)
);

AO32x1_ASAP7_75t_L g1067 ( 
.A1(n_837),
.A2(n_816),
.A3(n_866),
.B1(n_863),
.B2(n_873),
.Y(n_1067)
);

BUFx5_ASAP7_75t_L g1068 ( 
.A(n_830),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_874),
.B(n_877),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_831),
.A2(n_490),
.B(n_472),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_878),
.A2(n_490),
.B(n_472),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_775),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_897),
.B(n_456),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_802),
.B(n_542),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_861),
.A2(n_613),
.B1(n_900),
.B2(n_854),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_854),
.A2(n_900),
.B(n_786),
.C(n_613),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_854),
.B(n_479),
.C(n_900),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_854),
.A2(n_900),
.B(n_786),
.C(n_613),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_922),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_766),
.Y(n_1080)
);

INVx3_ASAP7_75t_SL g1081 ( 
.A(n_803),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_788),
.A2(n_515),
.B(n_776),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_828),
.A2(n_490),
.B(n_472),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_802),
.A2(n_916),
.B1(n_531),
.B2(n_542),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_SL g1085 ( 
.A1(n_854),
.A2(n_500),
.B(n_900),
.C(n_935),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_1085),
.B(n_1078),
.C(n_1076),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_993),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1032),
.A2(n_1015),
.B(n_1028),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_974),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1083),
.A2(n_1069),
.B(n_1039),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1069),
.A2(n_1024),
.B(n_1045),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1071),
.A2(n_964),
.B(n_1030),
.Y(n_1093)
);

BUFx4f_ASAP7_75t_L g1094 ( 
.A(n_1081),
.Y(n_1094)
);

INVx6_ASAP7_75t_SL g1095 ( 
.A(n_971),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_969),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_977),
.B(n_991),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1030),
.A2(n_1049),
.B(n_1063),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1074),
.B(n_1004),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_1022),
.B(n_1011),
.C(n_957),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_975),
.Y(n_1101)
);

AO31x2_ASAP7_75t_L g1102 ( 
.A1(n_976),
.A2(n_983),
.A3(n_1044),
.B(n_1058),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1014),
.B(n_948),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1084),
.A2(n_968),
.B1(n_1025),
.B2(n_951),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1082),
.A2(n_982),
.B(n_985),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_974),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_972),
.A2(n_1082),
.B(n_1052),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_966),
.A2(n_1009),
.B(n_1053),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_952),
.B(n_988),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1031),
.A2(n_1059),
.B(n_1066),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_1084),
.A2(n_1040),
.B(n_1020),
.C(n_1044),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1066),
.A2(n_1070),
.B(n_990),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_981),
.A2(n_1036),
.B(n_1048),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1050),
.A2(n_983),
.B(n_1002),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_954),
.A2(n_1001),
.B(n_949),
.C(n_1005),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_953),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_958),
.A2(n_1027),
.B(n_1038),
.C(n_1021),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1056),
.B(n_999),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1012),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1073),
.B(n_986),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1079),
.B(n_961),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1017),
.B(n_1026),
.Y(n_1123)
);

AND2x6_ASAP7_75t_L g1124 ( 
.A(n_959),
.B(n_970),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1034),
.A2(n_1067),
.B(n_1060),
.Y(n_1125)
);

AOI221x1_ASAP7_75t_L g1126 ( 
.A1(n_951),
.A2(n_1008),
.B1(n_1054),
.B2(n_978),
.C(n_980),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_995),
.B(n_962),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_948),
.B(n_1008),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1072),
.A2(n_1020),
.B1(n_1065),
.B2(n_984),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1051),
.A2(n_1061),
.B(n_1062),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_947),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_994),
.A2(n_984),
.B1(n_1029),
.B2(n_1000),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_SL g1133 ( 
.A(n_971),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1033),
.A2(n_1006),
.B(n_1064),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1046),
.B(n_1007),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1057),
.B(n_1043),
.C(n_1006),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_965),
.B(n_1012),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_SL g1138 ( 
.A1(n_1042),
.A2(n_1010),
.B(n_998),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_970),
.A2(n_971),
.B1(n_997),
.B2(n_1010),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_R g1140 ( 
.A(n_996),
.B(n_987),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1047),
.A2(n_1067),
.A3(n_1033),
.B(n_1016),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1067),
.A2(n_1018),
.A3(n_1019),
.B(n_1035),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_992),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1037),
.B(n_1041),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_967),
.A2(n_1080),
.B(n_1055),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_955),
.B(n_963),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_973),
.A2(n_1080),
.B(n_987),
.C(n_956),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1013),
.B(n_955),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_992),
.A2(n_953),
.B1(n_956),
.B2(n_979),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_953),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1019),
.A2(n_987),
.B(n_963),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_956),
.B(n_979),
.C(n_987),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1068),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1068),
.A2(n_1077),
.B(n_1075),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1068),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1068),
.A2(n_652),
.B(n_1032),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_977),
.B(n_313),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_977),
.B(n_313),
.Y(n_1159)
);

AO32x2_ASAP7_75t_L g1160 ( 
.A1(n_968),
.A2(n_983),
.A3(n_1025),
.B1(n_1084),
.B2(n_1044),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1077),
.A2(n_1075),
.B(n_977),
.C(n_1076),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_977),
.B(n_1084),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_996),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1010),
.B(n_987),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1077),
.A2(n_1085),
.B(n_1076),
.C(n_1078),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1077),
.A2(n_1075),
.B1(n_977),
.B2(n_446),
.C(n_613),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_974),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_977),
.B(n_1075),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1077),
.A2(n_1085),
.B(n_1076),
.C(n_1078),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1075),
.B(n_861),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_993),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1078),
.C(n_1022),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1017),
.B(n_1010),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1075),
.B(n_861),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_977),
.B(n_313),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1077),
.A2(n_1085),
.B(n_1076),
.C(n_1078),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1075),
.B(n_861),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_977),
.B(n_313),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_953),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1010),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_974),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1003),
.A2(n_950),
.B(n_989),
.Y(n_1192)
);

AO21x2_ASAP7_75t_L g1193 ( 
.A1(n_1082),
.A2(n_976),
.B(n_1015),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1075),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_976),
.A2(n_817),
.A3(n_983),
.B(n_1044),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1078),
.C(n_1022),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1075),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_977),
.B(n_313),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_975),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1204)
);

AOI211x1_ASAP7_75t_L g1205 ( 
.A1(n_1011),
.A2(n_938),
.B(n_909),
.C(n_957),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1078),
.C(n_1022),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1078),
.C(n_1022),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1077),
.B(n_1075),
.C(n_977),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1075),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_976),
.A2(n_817),
.A3(n_983),
.B(n_1044),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_SL g1213 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1078),
.C(n_1022),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1023),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_976),
.A2(n_817),
.A3(n_983),
.B(n_1044),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1017),
.B(n_1010),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1032),
.A2(n_652),
.B(n_602),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1169),
.A2(n_1097),
.B1(n_1209),
.B2(n_1171),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1090),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1209),
.A2(n_1164),
.B1(n_1210),
.B2(n_1194),
.Y(n_1222)
);

CKINVDCx8_ASAP7_75t_R g1223 ( 
.A(n_1131),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1164),
.A2(n_1210),
.B1(n_1194),
.B2(n_1200),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1165),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1162),
.A2(n_1184),
.B1(n_1181),
.B2(n_1174),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1146),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1170),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1105),
.A2(n_1200),
.B1(n_1158),
.B2(n_1182),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1120),
.Y(n_1230)
);

BUFx8_ASAP7_75t_L g1231 ( 
.A(n_1133),
.Y(n_1231)
);

OAI21xp33_ASAP7_75t_L g1232 ( 
.A1(n_1116),
.A2(n_1088),
.B(n_1204),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1146),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1202),
.Y(n_1234)
);

INVx6_ASAP7_75t_L g1235 ( 
.A(n_1150),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1107),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1105),
.A2(n_1198),
.B1(n_1088),
.B2(n_1204),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1159),
.A2(n_1201),
.B1(n_1187),
.B2(n_1198),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1136),
.A2(n_1128),
.B1(n_1099),
.B2(n_1110),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1150),
.B(n_1188),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1150),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1098),
.A2(n_1156),
.B(n_1092),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1136),
.A2(n_1099),
.B1(n_1121),
.B2(n_1103),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1103),
.A2(n_1114),
.B1(n_1106),
.B2(n_1115),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_1133),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1144),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1165),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1107),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1106),
.A2(n_1115),
.B1(n_1111),
.B2(n_1190),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1190),
.A2(n_1108),
.B1(n_1119),
.B2(n_1109),
.Y(n_1250)
);

BUFx4_ASAP7_75t_SL g1251 ( 
.A(n_1087),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1132),
.A2(n_1154),
.B1(n_1139),
.B2(n_1094),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_SL g1253 ( 
.A(n_1095),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1138),
.A2(n_1127),
.B1(n_1135),
.B2(n_1093),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1122),
.A2(n_1094),
.B1(n_1129),
.B2(n_1124),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1129),
.A2(n_1124),
.B1(n_1175),
.B2(n_1137),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1096),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1117),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1095),
.A2(n_1193),
.B1(n_1113),
.B2(n_1216),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1142),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1142),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1150),
.Y(n_1262)
);

BUFx4f_ASAP7_75t_L g1263 ( 
.A(n_1166),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1123),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1124),
.A2(n_1160),
.B1(n_1213),
.B2(n_1208),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1193),
.A2(n_1124),
.B1(n_1205),
.B2(n_1100),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1117),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1141),
.Y(n_1268)
);

BUFx4f_ASAP7_75t_SL g1269 ( 
.A(n_1177),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1143),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1117),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1188),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1177),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1118),
.A2(n_1148),
.B1(n_1154),
.B2(n_1167),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1160),
.A2(n_1176),
.B1(n_1207),
.B2(n_1199),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1188),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1152),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1152),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1141),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1086),
.B1(n_1173),
.B2(n_1183),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1188),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1189),
.A2(n_1091),
.B1(n_1218),
.B2(n_1130),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1149),
.A2(n_1126),
.B1(n_1189),
.B2(n_1146),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1166),
.B(n_1147),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1089),
.A2(n_1125),
.B1(n_1145),
.B2(n_1153),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1151),
.B(n_1134),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1140),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1155),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1112),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1197),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1197),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1197),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1212),
.Y(n_1293)
);

CKINVDCx14_ASAP7_75t_R g1294 ( 
.A(n_1102),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1157),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1161),
.A2(n_1219),
.B1(n_1215),
.B2(n_1214),
.Y(n_1296)
);

CKINVDCx16_ASAP7_75t_R g1297 ( 
.A(n_1102),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1172),
.A2(n_1206),
.B1(n_1203),
.B2(n_1196),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1178),
.A2(n_1186),
.B1(n_1211),
.B2(n_1195),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1102),
.B(n_1217),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1104),
.A2(n_1163),
.B1(n_1168),
.B2(n_1179),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1212),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1180),
.A2(n_1185),
.B1(n_1191),
.B2(n_1192),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1217),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1217),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1170),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1165),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1170),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1090),
.Y(n_1309)
);

INVx8_ASAP7_75t_L g1310 ( 
.A(n_1150),
.Y(n_1310)
);

BUFx8_ASAP7_75t_L g1311 ( 
.A(n_1133),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1164),
.A2(n_1075),
.B1(n_977),
.B2(n_1169),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1313)
);

NAND2x1p5_ASAP7_75t_L g1314 ( 
.A(n_1150),
.B(n_1188),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1170),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1094),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1101),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1169),
.A2(n_1077),
.B1(n_977),
.B2(n_1075),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1101),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1101),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

INVx5_ASAP7_75t_L g1322 ( 
.A(n_1146),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1101),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1164),
.A2(n_1075),
.B1(n_977),
.B2(n_1169),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1171),
.A2(n_1077),
.B1(n_1169),
.B2(n_1209),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1162),
.A2(n_977),
.B(n_1077),
.Y(n_1326)
);

AOI21xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1158),
.A2(n_480),
.B(n_977),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1170),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1150),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1150),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1150),
.Y(n_1331)
);

INVx3_ASAP7_75t_SL g1332 ( 
.A(n_1107),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1164),
.A2(n_1075),
.B1(n_977),
.B2(n_1169),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1169),
.A2(n_977),
.B1(n_1164),
.B2(n_968),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1090),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1286),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1290),
.Y(n_1337)
);

BUFx2_ASAP7_75t_SL g1338 ( 
.A(n_1227),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1292),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1260),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1293),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1260),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1268),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1242),
.A2(n_1303),
.B(n_1301),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1299),
.A2(n_1326),
.B(n_1261),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1224),
.A2(n_1325),
.B(n_1222),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1286),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1300),
.B(n_1294),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1227),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1294),
.B(n_1297),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1302),
.B(n_1279),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1304),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1304),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1332),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1244),
.B(n_1224),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1325),
.A2(n_1222),
.B(n_1318),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1234),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1228),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1301),
.A2(n_1303),
.B(n_1298),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1227),
.B(n_1233),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1227),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1317),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1319),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1320),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1323),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1332),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_1308),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1233),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1306),
.Y(n_1371)
);

AOI21xp33_ASAP7_75t_L g1372 ( 
.A1(n_1312),
.A2(n_1333),
.B(n_1324),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1316),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1315),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1249),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1233),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1295),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1274),
.A2(n_1226),
.B(n_1220),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1305),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1296),
.A2(n_1298),
.B(n_1285),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1334),
.A2(n_1229),
.B1(n_1238),
.B2(n_1232),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1277),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1278),
.A2(n_1288),
.B(n_1313),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1236),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1305),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1291),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1322),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1322),
.B(n_1282),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1322),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1259),
.A2(n_1282),
.B(n_1266),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1266),
.A2(n_1250),
.B(n_1275),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1322),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1284),
.A2(n_1246),
.B(n_1267),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1231),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1309),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1271),
.A2(n_1289),
.B(n_1280),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1275),
.A2(n_1254),
.B(n_1280),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1265),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1289),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1239),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1239),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1254),
.B(n_1252),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1329),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1327),
.A2(n_1264),
.B1(n_1328),
.B2(n_1335),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1348),
.B(n_1221),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1354),
.B(n_1273),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1344),
.A2(n_1380),
.B(n_1360),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1348),
.B(n_1221),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1357),
.A2(n_1255),
.B(n_1256),
.C(n_1263),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1373),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1357),
.A2(n_1263),
.B(n_1314),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1346),
.A2(n_1310),
.B(n_1314),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_SL g1416 ( 
.A(n_1338),
.B(n_1331),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1359),
.B(n_1384),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1348),
.B(n_1230),
.Y(n_1418)
);

AO32x2_ASAP7_75t_L g1419 ( 
.A1(n_1362),
.A2(n_1394),
.A3(n_1376),
.B1(n_1370),
.B2(n_1382),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_SL g1420 ( 
.A1(n_1378),
.A2(n_1329),
.B(n_1245),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1358),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1372),
.A2(n_1230),
.B(n_1310),
.C(n_1331),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1337),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1381),
.A2(n_1307),
.B1(n_1270),
.B2(n_1310),
.C(n_1331),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1371),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1345),
.B(n_1276),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1381),
.A2(n_1223),
.B1(n_1269),
.B2(n_1253),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1351),
.B(n_1258),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1346),
.A2(n_1331),
.B1(n_1240),
.B2(n_1251),
.C(n_1231),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1354),
.B(n_1245),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1345),
.B(n_1240),
.Y(n_1431)
);

NAND2x1_ASAP7_75t_L g1432 ( 
.A(n_1361),
.B(n_1262),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1339),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1351),
.B(n_1330),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1372),
.A2(n_1231),
.B(n_1311),
.C(n_1245),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1351),
.B(n_1366),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1371),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1366),
.B(n_1272),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1377),
.A2(n_1287),
.B1(n_1330),
.B2(n_1241),
.Y(n_1439)
);

AND2x4_ASAP7_75t_SL g1440 ( 
.A(n_1384),
.B(n_1311),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1272),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1406),
.A2(n_1311),
.B1(n_1225),
.B2(n_1247),
.C(n_1257),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1359),
.B(n_1225),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1387),
.B(n_1247),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1339),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1377),
.B(n_1407),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1366),
.B(n_1235),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1353),
.B(n_1241),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1349),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_1358),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1353),
.B(n_1281),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1377),
.A2(n_1287),
.B1(n_1281),
.B2(n_1321),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1361),
.B(n_1257),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1358),
.B(n_1363),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1404),
.A2(n_1399),
.B(n_1386),
.C(n_1350),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_R g1458 ( 
.A(n_1378),
.B(n_1396),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1392),
.A2(n_1344),
.B(n_1360),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1360),
.A2(n_1378),
.B(n_1383),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1392),
.A2(n_1393),
.B(n_1399),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1341),
.Y(n_1462)
);

NOR2xp67_ASAP7_75t_L g1463 ( 
.A(n_1347),
.B(n_1395),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1404),
.A2(n_1350),
.B(n_1386),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1355),
.B(n_1368),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1382),
.Y(n_1466)
);

OAI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1406),
.A2(n_1403),
.B(n_1402),
.C(n_1401),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_SL g1468 ( 
.A(n_1338),
.B(n_1383),
.Y(n_1468)
);

CKINVDCx14_ASAP7_75t_R g1469 ( 
.A(n_1396),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_SL g1470 ( 
.A1(n_1398),
.A2(n_1388),
.B(n_1395),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1336),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1423),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1423),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1433),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1461),
.B(n_1345),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1461),
.B(n_1345),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1425),
.B(n_1382),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1461),
.B(n_1345),
.Y(n_1480)
);

NAND2x1_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1361),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1340),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1450),
.B(n_1340),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1340),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1446),
.A2(n_1401),
.B1(n_1356),
.B2(n_1403),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1466),
.B(n_1342),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1436),
.B(n_1375),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1436),
.B(n_1375),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1456),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1421),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1412),
.A2(n_1400),
.B1(n_1401),
.B2(n_1388),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1437),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1437),
.B(n_1365),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1456),
.B(n_1365),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1457),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1445),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1455),
.A2(n_1400),
.B1(n_1388),
.B2(n_1356),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1445),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1462),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1429),
.B(n_1407),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1463),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1464),
.A2(n_1402),
.B(n_1399),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1459),
.B(n_1343),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1459),
.B(n_1343),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1467),
.B(n_1347),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1471),
.B(n_1367),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1482),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1498),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1490),
.Y(n_1509)
);

INVx5_ASAP7_75t_SL g1510 ( 
.A(n_1472),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1495),
.B(n_1419),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1498),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1473),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1473),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1487),
.B(n_1417),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1491),
.A2(n_1427),
.B1(n_1458),
.B2(n_1388),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1482),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1482),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1474),
.Y(n_1519)
);

NAND4xp25_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1442),
.C(n_1424),
.D(n_1435),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1488),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1495),
.B(n_1489),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1495),
.B(n_1419),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1503),
.B(n_1504),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1492),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1474),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1492),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1489),
.B(n_1419),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1479),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1483),
.B(n_1419),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1490),
.Y(n_1531)
);

NAND4xp25_ASAP7_75t_L g1532 ( 
.A(n_1502),
.B(n_1465),
.C(n_1444),
.D(n_1443),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1475),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1481),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1419),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_1460),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1479),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1485),
.A2(n_1398),
.B1(n_1379),
.B2(n_1385),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1460),
.Y(n_1539)
);

OAI322xp33_ASAP7_75t_L g1540 ( 
.A1(n_1497),
.A2(n_1379),
.A3(n_1385),
.B1(n_1397),
.B2(n_1374),
.C1(n_1355),
.C2(n_1368),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1505),
.A2(n_1398),
.B1(n_1422),
.B2(n_1469),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1476),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1490),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1483),
.B(n_1459),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1476),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1524),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1524),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1477),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1477),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1477),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1513),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1513),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1516),
.B(n_1505),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1536),
.B(n_1506),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1534),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1514),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1523),
.B(n_1478),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1478),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1537),
.B(n_1502),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1497),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1496),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1508),
.B(n_1496),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_R g1567 ( 
.A(n_1515),
.B(n_1413),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1430),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_L g1569 ( 
.A(n_1540),
.B(n_1453),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1510),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1535),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1530),
.B(n_1484),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1539),
.B(n_1493),
.Y(n_1573)
);

NAND4xp25_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1500),
.C(n_1428),
.D(n_1397),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1508),
.B(n_1499),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1539),
.B(n_1493),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1519),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1521),
.B(n_1486),
.Y(n_1578)
);

AND2x2_ASAP7_75t_SL g1579 ( 
.A(n_1523),
.B(n_1453),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1512),
.B(n_1499),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1530),
.B(n_1478),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1480),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1551),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1562),
.B(n_1532),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1554),
.Y(n_1585)
);

AOI21xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1567),
.A2(n_1568),
.B(n_1516),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1562),
.A2(n_1532),
.A3(n_1541),
.B(n_1538),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1574),
.A2(n_1541),
.B(n_1538),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1574),
.B(n_1534),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1515),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1566),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1551),
.Y(n_1593)
);

AND2x4_ASAP7_75t_SL g1594 ( 
.A(n_1570),
.B(n_1428),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1566),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

AOI31xp33_ASAP7_75t_L g1598 ( 
.A1(n_1569),
.A2(n_1453),
.A3(n_1430),
.B(n_1439),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1569),
.B(n_1522),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1552),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1512),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1534),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1452),
.B1(n_1481),
.B2(n_1448),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1553),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1558),
.B(n_1507),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1563),
.B(n_1522),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1528),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.B(n_1528),
.Y(n_1612)
);

NAND2x1_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1528),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1553),
.Y(n_1614)
);

INVxp33_ASAP7_75t_L g1615 ( 
.A(n_1563),
.Y(n_1615)
);

NAND2x1_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_1546),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1578),
.B(n_1413),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1557),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1557),
.B(n_1426),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1547),
.B(n_1510),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1564),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1564),
.Y(n_1623)
);

AOI32xp33_ASAP7_75t_L g1624 ( 
.A1(n_1547),
.A2(n_1480),
.A3(n_1440),
.B1(n_1418),
.B2(n_1544),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1584),
.B(n_1572),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.B(n_1581),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1617),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1586),
.B(n_1555),
.Y(n_1635)
);

OAI322xp33_ASAP7_75t_L g1636 ( 
.A1(n_1599),
.A2(n_1573),
.A3(n_1576),
.B1(n_1555),
.B2(n_1575),
.C1(n_1580),
.C2(n_1565),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1581),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1581),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1588),
.A2(n_1451),
.B1(n_1448),
.B2(n_1480),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1590),
.B(n_1576),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1583),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1594),
.B(n_1430),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1594),
.B(n_1577),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_L g1645 ( 
.A(n_1589),
.B(n_1415),
.C(n_1414),
.D(n_1396),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1577),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1598),
.B(n_1615),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1593),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1600),
.Y(n_1651)
);

NAND5xp2_ASAP7_75t_L g1652 ( 
.A(n_1624),
.B(n_1434),
.C(n_1447),
.D(n_1438),
.E(n_1418),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1601),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1602),
.B(n_1575),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1507),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1606),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1619),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1604),
.A2(n_1448),
.B1(n_1451),
.B2(n_1409),
.Y(n_1659)
);

OAI322xp33_ASAP7_75t_L g1660 ( 
.A1(n_1631),
.A2(n_1613),
.A3(n_1621),
.B1(n_1616),
.B2(n_1608),
.C1(n_1619),
.C2(n_1623),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1635),
.A2(n_1613),
.B(n_1616),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1649),
.A2(n_1611),
.B1(n_1620),
.B2(n_1597),
.C(n_1596),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1625),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1626),
.B(n_1607),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1627),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1645),
.A2(n_1607),
.B1(n_1620),
.B2(n_1611),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1642),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1633),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1641),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1651),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1634),
.B(n_1607),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1657),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1639),
.A2(n_1623),
.B(n_1612),
.Y(n_1676)
);

OAI32xp33_ASAP7_75t_L g1677 ( 
.A1(n_1628),
.A2(n_1619),
.A3(n_1612),
.B1(n_1618),
.B2(n_1614),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1630),
.B(n_1622),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1659),
.A2(n_1621),
.B1(n_1510),
.B2(n_1440),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1632),
.B(n_1646),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1648),
.A2(n_1597),
.B(n_1517),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1625),
.A2(n_1510),
.B1(n_1582),
.B2(n_1501),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1644),
.A2(n_1426),
.B1(n_1396),
.B2(n_1431),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1661),
.A2(n_1658),
.B(n_1643),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1667),
.B(n_1673),
.Y(n_1686)
);

OA22x2_ASAP7_75t_L g1687 ( 
.A1(n_1665),
.A2(n_1658),
.B1(n_1637),
.B2(n_1630),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1673),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1676),
.A2(n_1629),
.B1(n_1640),
.B2(n_1654),
.C(n_1655),
.Y(n_1689)
);

AOI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1667),
.A2(n_1674),
.B(n_1681),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1674),
.A2(n_1637),
.B1(n_1638),
.B2(n_1647),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1664),
.B(n_1629),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1668),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1647),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1663),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1666),
.A2(n_1640),
.B1(n_1655),
.B2(n_1656),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1671),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1678),
.B(n_1656),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1662),
.A2(n_1517),
.B1(n_1525),
.B2(n_1510),
.Y(n_1701)
);

OAI32xp33_ASAP7_75t_L g1702 ( 
.A1(n_1660),
.A2(n_1636),
.A3(n_1525),
.B1(n_1549),
.B2(n_1559),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1672),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1675),
.B(n_1582),
.Y(n_1704)
);

NOR2xp67_ASAP7_75t_SL g1705 ( 
.A(n_1686),
.B(n_1682),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1694),
.B(n_1652),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1690),
.A2(n_1680),
.B1(n_1679),
.B2(n_1683),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1685),
.A2(n_1702),
.B(n_1677),
.C(n_1701),
.Y(n_1708)
);

XNOR2x2_ASAP7_75t_L g1709 ( 
.A(n_1687),
.B(n_1684),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1685),
.A2(n_1525),
.B(n_1684),
.C(n_1410),
.Y(n_1710)
);

OAI321xp33_ASAP7_75t_L g1711 ( 
.A1(n_1697),
.A2(n_1560),
.A3(n_1559),
.B1(n_1550),
.B2(n_1549),
.C(n_1548),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1560),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1688),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1691),
.B(n_1560),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1700),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1708),
.A2(n_1692),
.B(n_1701),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1715),
.B(n_1687),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1713),
.B(n_1693),
.Y(n_1718)
);

O2A1O1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1709),
.A2(n_1703),
.B(n_1699),
.C(n_1698),
.Y(n_1719)
);

INVxp33_ASAP7_75t_L g1720 ( 
.A(n_1705),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1707),
.A2(n_1689),
.B(n_1695),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1712),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1714),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1706),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1719),
.A2(n_1711),
.B1(n_1710),
.B2(n_1704),
.C(n_1369),
.Y(n_1725)
);

AOI322xp5_ASAP7_75t_L g1726 ( 
.A1(n_1717),
.A2(n_1711),
.A3(n_1559),
.B1(n_1550),
.B2(n_1548),
.C1(n_1549),
.C2(n_1527),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_L g1727 ( 
.A1(n_1719),
.A2(n_1716),
.B(n_1721),
.C(n_1718),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1723),
.A2(n_1724),
.B1(n_1720),
.B2(n_1722),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_R g1729 ( 
.A(n_1724),
.B(n_1387),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1729),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1727),
.A2(n_1369),
.B(n_1501),
.C(n_1550),
.Y(n_1731)
);

NOR5xp2_ASAP7_75t_L g1732 ( 
.A(n_1726),
.B(n_1531),
.C(n_1374),
.D(n_1545),
.E(n_1526),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1728),
.A2(n_1725),
.B1(n_1510),
.B2(n_1548),
.Y(n_1733)
);

OAI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1727),
.A2(n_1409),
.B(n_1408),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1727),
.B(n_1451),
.C(n_1408),
.D(n_1411),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1735),
.B(n_1507),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1733),
.B(n_1432),
.C(n_1411),
.Y(n_1737)
);

XOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1730),
.B(n_1409),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1518),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1731),
.B(n_1420),
.Y(n_1740)
);

OAI21xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1736),
.A2(n_1732),
.B(n_1518),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1739),
.B(n_1518),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1738),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1743),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1744),
.A2(n_1740),
.B1(n_1737),
.B2(n_1741),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1745),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1742),
.B(n_1420),
.Y(n_1748)
);

AO221x1_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1470),
.B1(n_1405),
.B2(n_1449),
.C(n_1543),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1545),
.B1(n_1526),
.B2(n_1542),
.C(n_1533),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1524),
.B1(n_1544),
.B2(n_1509),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1750),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_R g1753 ( 
.A1(n_1751),
.A2(n_1470),
.B1(n_1524),
.B2(n_1468),
.C(n_1416),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1752),
.B(n_1391),
.C(n_1389),
.Y(n_1754)
);


endmodule