module fake_ariane_1378_n_2021 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2021);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2021;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_80),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_109),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_55),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_114),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_67),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_143),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_117),
.Y(n_223)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_158),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_52),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_27),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_111),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_51),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_19),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_62),
.Y(n_236)
);

INVx4_ASAP7_75t_R g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_65),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_99),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_66),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_77),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_39),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_122),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_145),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_16),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_41),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_184),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_178),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_102),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_85),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_28),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_123),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_35),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_106),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_74),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_72),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_19),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_130),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_91),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_98),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_36),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_120),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_110),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_142),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_164),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_185),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_58),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_144),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_198),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_40),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_149),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_31),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_166),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_43),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_128),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_81),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_44),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_32),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_127),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_104),
.Y(n_311)
);

BUFx8_ASAP7_75t_SL g312 ( 
.A(n_96),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_139),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_167),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_112),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_196),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_194),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_87),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_169),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_118),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_30),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_68),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_78),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_24),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_86),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_31),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_26),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_161),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_50),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_36),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_125),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_64),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_17),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_129),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_64),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_103),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_177),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_75),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_70),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_62),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_49),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_69),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_165),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_188),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_95),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_20),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_53),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_42),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_25),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_56),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_197),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_82),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_54),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_65),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_24),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_50),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_55),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_199),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_195),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_92),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_101),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_191),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_33),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_180),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_57),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_13),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_12),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_89),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_107),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_72),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_173),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_26),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_135),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_28),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_181),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_84),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_108),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_0),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_6),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_53),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_121),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_51),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_38),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_152),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_63),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_90),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_76),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_2),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_131),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_137),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_88),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_23),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_146),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_56),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_14),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_8),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_10),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_1),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_27),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_6),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_244),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_308),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_207),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_229),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_308),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_223),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_346),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_244),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_274),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_207),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_274),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_292),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_292),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_308),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_275),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_308),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_308),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_360),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_368),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_284),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_299),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_205),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_234),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_239),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_273),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_218),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_226),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_234),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_233),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_236),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_242),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_276),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_271),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_276),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_293),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_218),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_250),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_261),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_324),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_297),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_302),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_309),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_272),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_322),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_208),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_327),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_324),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_328),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_334),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_336),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_357),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_358),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_318),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_225),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_250),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_267),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_324),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_267),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_304),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_207),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_280),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_304),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_208),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_391),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_225),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_225),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_287),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_295),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_287),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_319),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_313),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_231),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_214),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_316),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_319),
.Y(n_503)
);

INVxp33_ASAP7_75t_SL g504 ( 
.A(n_214),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_231),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_335),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_220),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_231),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_266),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_266),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_352),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_326),
.B1(n_401),
.B2(n_256),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_425),
.Y(n_514)
);

BUFx12f_ASAP7_75t_L g515 ( 
.A(n_403),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_209),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_467),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_436),
.B(n_352),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_460),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_469),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_434),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_405),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_417),
.B(n_211),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_460),
.B(n_337),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_424),
.B(n_213),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_458),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_467),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_410),
.A2(n_227),
.B(n_221),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_464),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_406),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_488),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_405),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_325),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_408),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_243),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_408),
.B(n_337),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_448),
.B(n_452),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_418),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_420),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_496),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_457),
.B(n_377),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_499),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_405),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_245),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_421),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_423),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_502),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_454),
.B(n_353),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_402),
.B(n_266),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_506),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_454),
.B(n_246),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_429),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_412),
.B(n_220),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_414),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_431),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_409),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_465),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_413),
.B(n_228),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_437),
.A2(n_400),
.B1(n_396),
.B2(n_395),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_433),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_414),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_435),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_435),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_503),
.B(n_353),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_447),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_438),
.A2(n_331),
.B1(n_393),
.B2(n_340),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_438),
.Y(n_596)
);

CKINVDCx8_ASAP7_75t_R g597 ( 
.A(n_484),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_521),
.B(n_432),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_465),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_522),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_522),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_557),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_411),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_564),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_518),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_518),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_523),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_554),
.B(n_479),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

CKINVDCx12_ASAP7_75t_R g615 ( 
.A(n_581),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_577),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_520),
.B(n_411),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_563),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_520),
.B(n_479),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_576),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_493),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_539),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_594),
.A2(n_475),
.B1(n_426),
.B2(n_419),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_577),
.B(n_422),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_576),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_532),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_513),
.A2(n_426),
.B1(n_419),
.B2(n_475),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_567),
.B(n_415),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_528),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_517),
.A2(n_504),
.B1(n_422),
.B2(n_501),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_539),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_567),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_590),
.B(n_493),
.Y(n_640)
);

INVx11_ASAP7_75t_L g641 ( 
.A(n_540),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_530),
.B(n_500),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_583),
.A2(n_504),
.B1(n_459),
.B2(n_490),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_579),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_590),
.B(n_500),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_571),
.B(n_505),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_548),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_525),
.B(n_505),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_582),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_545),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_584),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_512),
.B(n_508),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_548),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_597),
.B(n_508),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_545),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_550),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_526),
.A2(n_510),
.B1(n_509),
.B2(n_495),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_512),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_545),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_586),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_512),
.B(n_509),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_587),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_550),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_551),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_588),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_519),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_571),
.B(n_510),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_551),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_532),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_545),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_519),
.A2(n_444),
.B1(n_440),
.B2(n_495),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_588),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_580),
.A2(n_491),
.B1(n_235),
.B2(n_238),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_578),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_589),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_519),
.B(n_497),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_526),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_553),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_545),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_541),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_553),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_580),
.B(n_538),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_559),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_560),
.B(n_204),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_515),
.B(n_416),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_560),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_538),
.B(n_204),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_515),
.B(n_443),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_593),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_527),
.B(n_445),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

BUFx6f_ASAP7_75t_SL g704 ( 
.A(n_526),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_561),
.A2(n_498),
.B(n_497),
.Y(n_705)
);

INVx8_ASAP7_75t_L g706 ( 
.A(n_545),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_591),
.B(n_206),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_562),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_516),
.B(n_446),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_596),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_562),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_578),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_593),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_546),
.B(n_498),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_552),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_511),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_592),
.A2(n_449),
.B1(n_451),
.B2(n_450),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_511),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_544),
.B(n_453),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_591),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_514),
.Y(n_721)
);

INVx6_ASAP7_75t_L g722 ( 
.A(n_572),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_545),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_514),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_566),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_529),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_529),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_533),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_536),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_455),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_569),
.B(n_461),
.Y(n_731)
);

AO21x2_ASAP7_75t_L g732 ( 
.A1(n_531),
.A2(n_252),
.B(n_248),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_524),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_597),
.B(n_462),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_533),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_535),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_535),
.B(n_556),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_556),
.B(n_489),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_524),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_573),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_573),
.B(n_463),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_574),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_574),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_540),
.B(n_206),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_595),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_531),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_536),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_566),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_566),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_634),
.A2(n_566),
.B1(n_540),
.B2(n_468),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_654),
.B(n_659),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_604),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_652),
.B(n_566),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_599),
.B(n_566),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_599),
.B(n_566),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_620),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_598),
.B(n_555),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_654),
.B(n_212),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_677),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_609),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_702),
.B(n_210),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_620),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_642),
.B(n_607),
.C(n_612),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_709),
.B(n_259),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_663),
.B(n_392),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_628),
.B(n_257),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_654),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_608),
.Y(n_768)
);

BUFx6f_ASAP7_75t_SL g769 ( 
.A(n_616),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_640),
.B(n_258),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_608),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_654),
.B(n_212),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_648),
.B(n_264),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_720),
.A2(n_235),
.B1(n_238),
.B2(n_228),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_610),
.A2(n_232),
.B(n_254),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_621),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_659),
.Y(n_777)
);

NAND2x1_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_524),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_677),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_720),
.B(n_598),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_611),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_659),
.B(n_215),
.Y(n_782)
);

NAND3x1_ASAP7_75t_L g783 ( 
.A(n_734),
.B(n_565),
.C(n_555),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_639),
.A2(n_343),
.B1(n_347),
.B2(n_240),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_673),
.B(n_215),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_621),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_677),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_639),
.B(n_216),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_656),
.B(n_265),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_625),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_617),
.B(n_343),
.C(n_240),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_636),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_710),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_693),
.A2(n_216),
.B1(n_219),
.B2(n_217),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_613),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_613),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_685),
.B(n_217),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_625),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_616),
.B(n_568),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_630),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_644),
.B(n_568),
.C(n_349),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_619),
.B(n_219),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_710),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_222),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_681),
.B(n_222),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_270),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_712),
.B(n_230),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_690),
.B(n_279),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_719),
.B(n_230),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_241),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_731),
.B(n_241),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_635),
.B(n_249),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_677),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_635),
.B(n_249),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_738),
.B(n_251),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_649),
.A2(n_251),
.B1(n_394),
.B2(n_344),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_738),
.B(n_622),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_714),
.B(n_344),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_684),
.B(n_359),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_619),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_603),
.B(n_359),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_626),
.B(n_361),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_603),
.B(n_361),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_601),
.B(n_369),
.Y(n_825)
);

AOI22x1_ASAP7_75t_L g826 ( 
.A1(n_626),
.A2(n_366),
.B1(n_371),
.B2(n_367),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_627),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_629),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_601),
.B(n_369),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_674),
.B(n_282),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_602),
.B(n_374),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_637),
.B(n_350),
.C(n_348),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_R g833 ( 
.A(n_600),
.B(n_350),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_746),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_710),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_627),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_602),
.B(n_374),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_629),
.A2(n_466),
.B1(n_470),
.B2(n_471),
.Y(n_838)
);

NAND2x1_ASAP7_75t_L g839 ( 
.A(n_725),
.B(n_547),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_632),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_616),
.B(n_710),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_638),
.B(n_376),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_631),
.B(n_472),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_638),
.B(n_376),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_632),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_645),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_473),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_643),
.A2(n_481),
.B1(n_474),
.B2(n_478),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_643),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_646),
.B(n_388),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_646),
.B(n_388),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_651),
.B(n_390),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_651),
.B(n_390),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_657),
.B(n_394),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_704),
.B(n_286),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_705),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_645),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_636),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_657),
.B(n_281),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_660),
.B(n_294),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_660),
.B(n_296),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_670),
.B(n_288),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_704),
.B(n_300),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_678),
.A2(n_224),
.B1(n_289),
.B2(n_291),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_670),
.B(n_298),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_671),
.B(n_303),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_704),
.B(n_305),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_647),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_658),
.B(n_476),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_675),
.B(n_306),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_686),
.B(n_321),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_707),
.B(n_330),
.Y(n_872)
);

OAI221xp5_ASAP7_75t_L g873 ( 
.A1(n_662),
.A2(n_373),
.B1(n_351),
.B2(n_354),
.C(n_355),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_686),
.B(n_307),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_689),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_689),
.B(n_314),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_691),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_677),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_647),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_691),
.B(n_333),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_692),
.B(n_320),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_692),
.A2(n_363),
.B(n_362),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_678),
.B(n_477),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_695),
.B(n_699),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_650),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_695),
.A2(n_480),
.B(n_485),
.C(n_483),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_696),
.B(n_351),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_600),
.Y(n_888)
);

OAI22xp33_ASAP7_75t_SL g889 ( 
.A1(n_744),
.A2(n_396),
.B1(n_354),
.B2(n_400),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_678),
.A2(n_365),
.B1(n_370),
.B2(n_372),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_678),
.B(n_482),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_699),
.B(n_355),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_708),
.B(n_356),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_708),
.B(n_356),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_711),
.B(n_378),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_605),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_711),
.A2(n_387),
.B(n_572),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_650),
.B(n_364),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_694),
.B(n_486),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_716),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_653),
.A2(n_371),
.B1(n_367),
.B2(n_366),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_605),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_653),
.B(n_364),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_655),
.A2(n_310),
.B1(n_253),
.B2(n_255),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_687),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_661),
.B(n_664),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_661),
.B(n_664),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_666),
.B(n_381),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_725),
.B(n_311),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_606),
.B(n_381),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_716),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_666),
.B(n_383),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_762),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_752),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_763),
.A2(n_807),
.B1(n_790),
.B2(n_766),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_833),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_833),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_761),
.B(n_680),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_790),
.A2(n_615),
.B1(n_747),
.B2(n_633),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_818),
.B(n_668),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_878),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_834),
.A2(n_746),
.B(n_669),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_764),
.B(n_668),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_847),
.B(n_694),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_768),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_767),
.B(n_725),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_767),
.B(n_725),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_858),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_766),
.B(n_669),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_756),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_771),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_776),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_770),
.B(n_773),
.Y(n_933)
);

INVx5_ASAP7_75t_L g934 ( 
.A(n_759),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_906),
.A2(n_713),
.B1(n_701),
.B2(n_682),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_770),
.B(n_773),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_777),
.B(n_907),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_843),
.B(n_694),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_786),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_791),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_891),
.A2(n_721),
.B1(n_724),
.B2(n_726),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_799),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_807),
.B(n_700),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_869),
.B(n_700),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_810),
.B(n_672),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_777),
.B(n_672),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_811),
.B(n_679),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_878),
.B(n_665),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_759),
.B(n_679),
.Y(n_949)
);

NOR2x2_ASAP7_75t_L g950 ( 
.A(n_774),
.B(n_700),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_796),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_812),
.B(n_682),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_827),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_836),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_765),
.B(n_683),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_793),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_780),
.B(n_633),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_888),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_888),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_796),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_896),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_700),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_840),
.B(n_683),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_845),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_800),
.B(n_676),
.Y(n_965)
);

AND2x6_ASAP7_75t_SL g966 ( 
.A(n_887),
.B(n_700),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_757),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_846),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_857),
.B(n_701),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_868),
.Y(n_970)
);

AND2x6_ASAP7_75t_SL g971 ( 
.A(n_887),
.B(n_676),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_902),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_879),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_841),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_885),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_750),
.A2(n_726),
.B1(n_724),
.B2(n_736),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_794),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_788),
.B(n_615),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_828),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_828),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_884),
.A2(n_713),
.B(n_614),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_759),
.B(n_749),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_899),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_783),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_SL g985 ( 
.A1(n_750),
.A2(n_715),
.B1(n_729),
.B2(n_747),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_875),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_816),
.B(n_741),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_899),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_875),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_819),
.B(n_883),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_801),
.A2(n_729),
.B1(n_748),
.B2(n_749),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_L g992 ( 
.A(n_872),
.B(n_614),
.C(n_606),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_855),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_898),
.B(n_721),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_788),
.B(n_614),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_760),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_804),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_769),
.Y(n_998)
);

NOR2x2_ASAP7_75t_L g999 ( 
.A(n_774),
.B(n_641),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_835),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_813),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_792),
.B(n_623),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_900),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_759),
.B(n_748),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_815),
.B(n_623),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_903),
.B(n_736),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_SL g1007 ( 
.A1(n_873),
.A2(n_641),
.B1(n_383),
.B2(n_389),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_779),
.B(n_623),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_908),
.B(n_745),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_801),
.A2(n_687),
.B1(n_706),
.B2(n_745),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_784),
.A2(n_737),
.B(n_688),
.C(n_697),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_779),
.B(n_733),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_779),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_781),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_912),
.B(n_718),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_787),
.B(n_687),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_779),
.B(n_733),
.Y(n_1017)
);

BUFx2_ASAP7_75t_SL g1018 ( 
.A(n_769),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_809),
.B(n_718),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_911),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_754),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_789),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_797),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_814),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_832),
.B(n_395),
.C(n_389),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_821),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_849),
.Y(n_1027)
);

NAND2x1_ASAP7_75t_SL g1028 ( 
.A(n_863),
.B(n_705),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_877),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_872),
.A2(n_687),
.B1(n_706),
.B2(n_717),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_755),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_814),
.B(n_905),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_814),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_910),
.B(n_743),
.Y(n_1034)
);

INVx8_ASAP7_75t_L g1035 ( 
.A(n_905),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_867),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_867),
.B(n_624),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_910),
.B(n_743),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_802),
.A2(n_830),
.B1(n_809),
.B2(n_890),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_820),
.B(n_727),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_856),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_905),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_905),
.B(n_624),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_886),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_787),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_830),
.B(n_727),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_859),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_753),
.B(n_733),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_856),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_778),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_892),
.B(n_728),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_889),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_859),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_893),
.B(n_728),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_894),
.B(n_742),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_860),
.B(n_742),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_861),
.B(n_735),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_758),
.A2(n_739),
.B(n_732),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_862),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_862),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_839),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_871),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_880),
.B(n_740),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_826),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_817),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_798),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_909),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_805),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_901),
.B(n_703),
.C(n_697),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_909),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_751),
.B(n_739),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_751),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_865),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_758),
.B(n_772),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_785),
.B(n_739),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_865),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_866),
.Y(n_1077)
);

AND2x6_ASAP7_75t_SL g1078 ( 
.A(n_806),
.B(n_442),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_838),
.B(n_848),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_808),
.B(n_717),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_825),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_838),
.B(n_442),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_866),
.Y(n_1083)
);

XOR2xp5_ASAP7_75t_L g1084 ( 
.A(n_864),
.B(n_717),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_829),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_803),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_772),
.B(n_723),
.Y(n_1087)
);

INVx5_ASAP7_75t_L g1088 ( 
.A(n_782),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_870),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_782),
.B(n_723),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_803),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_848),
.B(n_624),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_823),
.B(n_688),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_842),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1035),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_922),
.A2(n_850),
.B(n_823),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_929),
.A2(n_852),
.B(n_850),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_956),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_933),
.A2(n_824),
.B(n_822),
.C(n_795),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_915),
.A2(n_775),
.B(n_882),
.C(n_844),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_988),
.B(n_456),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_936),
.B(n_993),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_913),
.B(n_904),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1039),
.A2(n_851),
.B1(n_853),
.B2(n_854),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1035),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_935),
.A2(n_852),
.B(n_837),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_924),
.B(n_687),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_965),
.B(n_456),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_916),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1001),
.B(n_870),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_918),
.A2(n_831),
.B(n_895),
.C(n_881),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_943),
.B(n_874),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_943),
.B(n_1079),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_917),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_919),
.B(n_723),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_937),
.A2(n_897),
.B(n_895),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_937),
.A2(n_881),
.B(n_876),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_920),
.B(n_874),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_924),
.B(n_876),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1058),
.A2(n_703),
.B(n_688),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_923),
.B(n_987),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_914),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_963),
.A2(n_706),
.B1(n_698),
.B2(n_618),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_945),
.A2(n_732),
.B(n_237),
.C(n_3),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1036),
.B(n_938),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1065),
.A2(n_706),
.B1(n_723),
.B2(n_665),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_944),
.B(n_1036),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_SL g1128 ( 
.A(n_978),
.B(n_706),
.Y(n_1128)
);

BUFx4f_ASAP7_75t_L g1129 ( 
.A(n_959),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_947),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1074),
.A2(n_698),
.B(n_618),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_952),
.A2(n_618),
.B(n_698),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_969),
.A2(n_698),
.B1(n_618),
.B2(n_665),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1048),
.A2(n_618),
.B(n_698),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_951),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_985),
.A2(n_665),
.B1(n_332),
.B2(n_260),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_998),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1002),
.A2(n_1075),
.B(n_995),
.C(n_1069),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_SL g1139 ( 
.A(n_1052),
.B(n_262),
.C(n_263),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_944),
.B(n_1085),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1019),
.A2(n_278),
.B(n_277),
.C(n_269),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_930),
.B(n_5),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1019),
.A2(n_268),
.B(n_339),
.C(n_329),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_930),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_938),
.B(n_5),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_990),
.B(n_7),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1094),
.B(n_7),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_951),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_978),
.A2(n_317),
.B1(n_283),
.B2(n_285),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_955),
.B(n_8),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_958),
.Y(n_1151)
);

BUFx12f_ASAP7_75t_L g1152 ( 
.A(n_983),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1074),
.A2(n_549),
.B(n_585),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1035),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1068),
.B(n_9),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_957),
.B(n_290),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_979),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_934),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_961),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_925),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_981),
.A2(n_1038),
.B(n_1034),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_926),
.A2(n_315),
.B(n_323),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1046),
.A2(n_301),
.B(n_247),
.C(n_207),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1046),
.B(n_931),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_928),
.B(n_962),
.Y(n_1165)
);

O2A1O1Ixp5_ASAP7_75t_SL g1166 ( 
.A1(n_1087),
.A2(n_311),
.B(n_575),
.C(n_585),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1041),
.A2(n_311),
.B(n_722),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_962),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_972),
.Y(n_1169)
);

BUFx4f_ASAP7_75t_L g1170 ( 
.A(n_1000),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_926),
.A2(n_572),
.B(n_345),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1042),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1013),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_977),
.B(n_1062),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_995),
.A2(n_207),
.B(n_247),
.C(n_345),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_994),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1066),
.B(n_312),
.Y(n_1177)
);

CKINVDCx8_ASAP7_75t_R g1178 ( 
.A(n_1018),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_958),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_974),
.B(n_13),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_927),
.A2(n_572),
.B(n_338),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1087),
.A2(n_549),
.B(n_585),
.Y(n_1182)
);

AOI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1064),
.A2(n_247),
.B1(n_338),
.B2(n_345),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_SL g1184 ( 
.A1(n_946),
.A2(n_15),
.B(n_18),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_979),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1080),
.A2(n_572),
.B(n_311),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_932),
.B(n_18),
.Y(n_1187)
);

AOI222xp33_ASAP7_75t_L g1188 ( 
.A1(n_984),
.A2(n_975),
.B1(n_940),
.B2(n_942),
.C1(n_953),
.C2(n_954),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_974),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_939),
.A2(n_722),
.B1(n_345),
.B2(n_338),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_964),
.A2(n_722),
.B1(n_345),
.B2(n_338),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_968),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_1002),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_970),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_973),
.B(n_21),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1066),
.B(n_23),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1084),
.B(n_29),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_SL g1198 ( 
.A1(n_946),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_986),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1006),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1200)
);

AND2x2_ASAP7_75t_SL g1201 ( 
.A(n_976),
.B(n_247),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_997),
.B(n_34),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1009),
.A2(n_247),
.B1(n_338),
.B2(n_42),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1025),
.A2(n_37),
.B(n_40),
.C(n_43),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_977),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_927),
.A2(n_572),
.B(n_585),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1078),
.B(n_37),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_967),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_934),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1081),
.B(n_45),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_949),
.A2(n_585),
.B(n_575),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_996),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1042),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_934),
.B(n_575),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1042),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1007),
.A2(n_46),
.B(n_47),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_986),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_949),
.A2(n_575),
.B(n_549),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1005),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1067),
.A2(n_311),
.A3(n_487),
.B(n_414),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1008),
.A2(n_575),
.B(n_549),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1081),
.A2(n_52),
.B(n_54),
.C(n_57),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1028),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1086),
.B(n_59),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_1012),
.A2(n_60),
.B(n_61),
.C(n_63),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_941),
.B(n_60),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1091),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_971),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1008),
.A2(n_549),
.B(n_547),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_941),
.B(n_1082),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1075),
.A2(n_547),
.B(n_414),
.C(n_487),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_991),
.B(n_61),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_966),
.B(n_66),
.Y(n_1233)
);

AOI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1049),
.A2(n_1041),
.B1(n_1061),
.B2(n_1050),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1014),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1071),
.A2(n_547),
.B(n_487),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_989),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_976),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1071),
.A2(n_547),
.B(n_487),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_SL g1240 ( 
.A(n_1093),
.B(n_71),
.C(n_311),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1092),
.B(n_71),
.Y(n_1241)
);

OAI21xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1045),
.A2(n_311),
.B(n_83),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1042),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1092),
.B(n_722),
.Y(n_1244)
);

AOI22x1_ASAP7_75t_L g1245 ( 
.A1(n_1061),
.A2(n_487),
.B1(n_113),
.B2(n_115),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1030),
.A2(n_79),
.B1(n_119),
.B2(n_124),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1022),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1015),
.A2(n_133),
.B(n_136),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1040),
.A2(n_140),
.B(n_141),
.Y(n_1249)
);

AOI22x1_ASAP7_75t_L g1250 ( 
.A1(n_1050),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1033),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1102),
.B(n_1023),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1161),
.A2(n_1090),
.B(n_1012),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1125),
.B(n_1037),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1097),
.A2(n_992),
.B(n_1056),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_1201),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1121),
.B(n_1140),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1144),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1232),
.B(n_999),
.C(n_1093),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1127),
.B(n_1027),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1164),
.B(n_1029),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1099),
.A2(n_1011),
.B(n_1051),
.C(n_1054),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1159),
.B(n_1076),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1109),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1170),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1113),
.A2(n_1010),
.B1(n_921),
.B2(n_1047),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1159),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1161),
.A2(n_1090),
.B(n_1057),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1153),
.A2(n_1032),
.B(n_1017),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1145),
.A2(n_1060),
.B1(n_1059),
.B2(n_1077),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1238),
.A2(n_950),
.B(n_1044),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1216),
.A2(n_1073),
.B(n_1053),
.C(n_1055),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1241),
.A2(n_1088),
.B1(n_1089),
.B2(n_1083),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1175),
.A2(n_1096),
.A3(n_1246),
.B(n_1231),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1114),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1123),
.A2(n_1017),
.B(n_1032),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1131),
.A2(n_1004),
.B(n_982),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_L g1278 ( 
.A1(n_1104),
.A2(n_1004),
.B(n_982),
.C(n_1070),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1197),
.B(n_1089),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_1026),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1212),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1241),
.A2(n_1088),
.B1(n_1083),
.B2(n_1016),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1178),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1111),
.A2(n_1063),
.B(n_1088),
.C(n_1070),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1251),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1168),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1188),
.B(n_1101),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1100),
.A2(n_1031),
.B(n_1021),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1122),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1138),
.A2(n_1016),
.B(n_1088),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1238),
.A2(n_1021),
.B(n_1031),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_R g1292 ( 
.A(n_1137),
.B(n_1033),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1129),
.B(n_1033),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1188),
.B(n_1026),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1107),
.B(n_1033),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1133),
.A2(n_1106),
.B(n_1132),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_L g1297 ( 
.A(n_1251),
.B(n_1072),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1230),
.A2(n_1020),
.B1(n_1003),
.B2(n_960),
.Y(n_1298)
);

AOI31xp67_ASAP7_75t_L g1299 ( 
.A1(n_1112),
.A2(n_1067),
.A3(n_989),
.B(n_1020),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1117),
.A2(n_980),
.B(n_1043),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1118),
.A2(n_1043),
.B(n_1024),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1142),
.B(n_1003),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1098),
.B(n_1072),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1167),
.A2(n_948),
.B(n_1072),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1072),
.A3(n_1013),
.B1(n_948),
.B2(n_171),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1210),
.A2(n_156),
.B(n_160),
.C(n_163),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1180),
.B(n_201),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1166),
.A2(n_176),
.B(n_182),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1234),
.A2(n_183),
.B(n_193),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_1158),
.B(n_1209),
.Y(n_1310)
);

AOI211x1_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_1195),
.B(n_1160),
.C(n_1192),
.Y(n_1311)
);

AND2x2_ASAP7_75t_SL g1312 ( 
.A(n_1233),
.B(n_1180),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1152),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1110),
.B(n_1169),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1119),
.B(n_1194),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1129),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1119),
.B(n_1165),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1251),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1228),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1235),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1150),
.A2(n_1143),
.B1(n_1141),
.B2(n_1226),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1146),
.A2(n_1242),
.B(n_1116),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1120),
.A2(n_1134),
.B(n_1236),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1124),
.A2(n_1149),
.B(n_1203),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1246),
.A2(n_1223),
.A3(n_1163),
.B(n_1133),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1177),
.B(n_1189),
.Y(n_1326)
);

O2A1O1Ixp5_ASAP7_75t_SL g1327 ( 
.A1(n_1120),
.A2(n_1249),
.B(n_1248),
.C(n_1247),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1186),
.A2(n_1239),
.B(n_1249),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1135),
.A2(n_1148),
.A3(n_1199),
.B(n_1217),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1221),
.A2(n_1229),
.B(n_1211),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1186),
.A2(n_1248),
.B(n_1218),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1103),
.B(n_1227),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1157),
.Y(n_1333)
);

AO22x2_ASAP7_75t_L g1334 ( 
.A1(n_1185),
.A2(n_1237),
.B1(n_1196),
.B2(n_1147),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_L g1335 ( 
.A(n_1107),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1172),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1107),
.A2(n_1244),
.B(n_1115),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1128),
.A2(n_1206),
.B(n_1171),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1181),
.A2(n_1245),
.B(n_1183),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1151),
.B(n_1179),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1154),
.B(n_1095),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1224),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1155),
.Y(n_1344)
);

BUFx4f_ASAP7_75t_L g1345 ( 
.A(n_1172),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1154),
.B(n_1095),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_1191),
.B(n_1193),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1204),
.A2(n_1240),
.B(n_1219),
.C(n_1130),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1126),
.A2(n_1162),
.B(n_1220),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1225),
.A2(n_1184),
.B(n_1200),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1158),
.A2(n_1209),
.B(n_1176),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1222),
.A2(n_1136),
.B(n_1250),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1220),
.A2(n_1207),
.A3(n_1198),
.B(n_1139),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1156),
.A2(n_1174),
.B(n_1173),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1220),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1173),
.A2(n_1214),
.B(n_1172),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1214),
.A2(n_1213),
.B(n_1215),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1202),
.B(n_1105),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1213),
.A2(n_1215),
.B(n_1243),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1243),
.A2(n_1105),
.B(n_1208),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_936),
.B(n_933),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1102),
.B(n_600),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1097),
.A2(n_936),
.B(n_933),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1153),
.A2(n_1131),
.B(n_1182),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1144),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1097),
.A2(n_936),
.B(n_933),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1201),
.A2(n_915),
.B1(n_936),
.B2(n_933),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1251),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1161),
.A2(n_1186),
.B(n_1231),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1161),
.A2(n_936),
.B(n_933),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1153),
.A2(n_1131),
.B(n_1182),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1251),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1232),
.B(n_936),
.C(n_933),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1175),
.A2(n_1096),
.A3(n_1058),
.B(n_1246),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1232),
.B(n_936),
.C(n_933),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1175),
.A2(n_1096),
.A3(n_1058),
.B(n_1246),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1109),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1161),
.A2(n_936),
.B(n_933),
.Y(n_1380)
);

AOI211x1_ASAP7_75t_L g1381 ( 
.A1(n_1216),
.A2(n_801),
.B(n_1238),
.C(n_873),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1097),
.A2(n_936),
.B(n_933),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1098),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1152),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1114),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1201),
.A2(n_915),
.B1(n_936),
.B2(n_933),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1161),
.A2(n_936),
.B(n_933),
.Y(n_1389)
);

AO32x2_ASAP7_75t_L g1390 ( 
.A1(n_1238),
.A2(n_1203),
.A3(n_1104),
.B1(n_1246),
.B2(n_985),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1391)
);

CKINVDCx16_ASAP7_75t_R g1392 ( 
.A(n_1152),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1140),
.B(n_636),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1102),
.B(n_600),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1125),
.A2(n_1065),
.B1(n_600),
.B2(n_633),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_SL g1396 ( 
.A1(n_1099),
.A2(n_933),
.B(n_936),
.C(n_915),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_933),
.B(n_936),
.C(n_943),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1125),
.A2(n_1065),
.B1(n_600),
.B2(n_633),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1170),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1125),
.B(n_943),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1153),
.A2(n_1131),
.B(n_1182),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1175),
.A2(n_1096),
.A3(n_1058),
.B(n_1246),
.Y(n_1403)
);

NOR4xp25_ASAP7_75t_L g1404 ( 
.A(n_1238),
.B(n_1219),
.C(n_1216),
.D(n_1130),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1197),
.B(n_1102),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1175),
.A2(n_1096),
.A3(n_1058),
.B(n_1246),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1161),
.A2(n_936),
.B(n_933),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1102),
.B(n_1121),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1102),
.A2(n_936),
.B(n_933),
.C(n_607),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1170),
.Y(n_1413)
);

AOI21xp33_ASAP7_75t_L g1414 ( 
.A1(n_1201),
.A2(n_936),
.B(n_933),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1109),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1264),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1281),
.Y(n_1417)
);

INVx4_ASAP7_75t_L g1418 ( 
.A(n_1345),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1385),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1415),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1299),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1363),
.A2(n_1394),
.B1(n_1259),
.B2(n_1399),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1387),
.B(n_1391),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1275),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1373),
.A2(n_1402),
.B(n_1323),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1338),
.A2(n_1322),
.B(n_1340),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1383),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1295),
.B(n_1285),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1375),
.A2(n_1377),
.B(n_1368),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1322),
.A2(n_1253),
.B(n_1269),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1375),
.A2(n_1377),
.B1(n_1395),
.B2(n_1388),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1318),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1289),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1327),
.A2(n_1255),
.B(n_1331),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1372),
.A2(n_1389),
.B(n_1380),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1366),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1329),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1255),
.A2(n_1328),
.B(n_1309),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1398),
.B(n_1407),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1370),
.B(n_1374),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1412),
.A2(n_1411),
.B1(n_1410),
.B2(n_1408),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1386),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1405),
.B(n_1279),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1401),
.B(n_1271),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1288),
.A2(n_1409),
.B(n_1367),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1276),
.A2(n_1277),
.B(n_1308),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_SL g1448 ( 
.A1(n_1414),
.A2(n_1348),
.B(n_1364),
.C(n_1382),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1304),
.A2(n_1290),
.B(n_1288),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1397),
.A2(n_1324),
.B(n_1367),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1320),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1364),
.A2(n_1382),
.B(n_1404),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1283),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1333),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1339),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1287),
.A2(n_1312),
.B1(n_1256),
.B2(n_1343),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1329),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1256),
.A2(n_1381),
.B1(n_1271),
.B2(n_1321),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1318),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1393),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1404),
.A2(n_1278),
.B(n_1396),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1267),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1339),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1267),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1291),
.A2(n_1257),
.B1(n_1252),
.B2(n_1326),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1379),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1314),
.B(n_1315),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1319),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1337),
.B(n_1282),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1300),
.A2(n_1371),
.B(n_1262),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1362),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1335),
.B(n_1345),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1302),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1294),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1272),
.A2(n_1350),
.B(n_1307),
.C(n_1306),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1332),
.A2(n_1344),
.B1(n_1390),
.B2(n_1280),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1263),
.B(n_1358),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1300),
.A2(n_1371),
.B(n_1268),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1268),
.A2(n_1270),
.B(n_1347),
.Y(n_1479)
);

AOI21xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1384),
.A2(n_1392),
.B(n_1400),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1356),
.A2(n_1357),
.B(n_1362),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1265),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1254),
.B(n_1266),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1350),
.A2(n_1298),
.B(n_1352),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1273),
.A2(n_1305),
.A3(n_1378),
.B(n_1406),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1370),
.B(n_1374),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1360),
.A2(n_1301),
.B(n_1351),
.Y(n_1488)
);

AOI21xp33_ASAP7_75t_L g1489 ( 
.A1(n_1334),
.A2(n_1349),
.B(n_1286),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1310),
.A2(n_1359),
.B(n_1354),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1303),
.B(n_1317),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1316),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1361),
.A2(n_1297),
.B(n_1341),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1311),
.A2(n_1335),
.B1(n_1341),
.B2(n_1413),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1376),
.A2(n_1406),
.B(n_1403),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1286),
.B(n_1336),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1325),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1313),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1305),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1342),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_SL g1501 ( 
.A1(n_1390),
.A2(n_1305),
.B(n_1325),
.C(n_1293),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1349),
.A2(n_1390),
.B(n_1346),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1292),
.B(n_1353),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1376),
.A2(n_1378),
.B(n_1403),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1353),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1376),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1378),
.A2(n_1403),
.B(n_1406),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1274),
.A2(n_1296),
.B(n_1330),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1274),
.A2(n_1296),
.B(n_1330),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1274),
.A2(n_1296),
.B(n_1330),
.Y(n_1510)
);

INVxp33_ASAP7_75t_SL g1511 ( 
.A(n_1275),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1281),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1405),
.B(n_1197),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1287),
.B(n_1258),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1296),
.A2(n_1373),
.B(n_1365),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1295),
.B(n_1241),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1281),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1375),
.A2(n_1377),
.B1(n_915),
.B2(n_936),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_L g1520 ( 
.A(n_1265),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1258),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1296),
.A2(n_1373),
.B(n_1365),
.Y(n_1522)
);

OAI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1375),
.A2(n_634),
.B1(n_936),
.B2(n_933),
.C(n_915),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1258),
.Y(n_1525)
);

BUFx4f_ASAP7_75t_SL g1526 ( 
.A(n_1264),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1368),
.A2(n_801),
.B1(n_630),
.B2(n_513),
.C(n_1388),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1375),
.A2(n_936),
.B(n_933),
.Y(n_1528)
);

AO31x2_ASAP7_75t_L g1529 ( 
.A1(n_1355),
.A2(n_1284),
.A3(n_1296),
.B(n_1253),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1335),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1299),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1296),
.A2(n_1373),
.B(n_1365),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_SL g1533 ( 
.A1(n_1368),
.A2(n_933),
.B(n_936),
.C(n_1388),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1368),
.A2(n_801),
.B1(n_630),
.B2(n_513),
.C(n_1388),
.Y(n_1534)
);

AO222x2_ASAP7_75t_L g1535 ( 
.A1(n_1405),
.A2(n_1197),
.B1(n_634),
.B2(n_801),
.C1(n_513),
.C2(n_630),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1405),
.B(n_1197),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1296),
.A2(n_1373),
.B(n_1365),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1281),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1375),
.A2(n_1201),
.B1(n_1377),
.B2(n_1287),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1372),
.A2(n_1389),
.B(n_1380),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1331),
.A2(n_1328),
.B(n_1355),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1375),
.A2(n_936),
.B(n_933),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1375),
.A2(n_1201),
.B1(n_1377),
.B2(n_1287),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1339),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1368),
.A2(n_801),
.B1(n_630),
.B2(n_513),
.C(n_1388),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1299),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1265),
.B(n_1151),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1372),
.A2(n_1389),
.B(n_1380),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1339),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1299),
.Y(n_1552)
);

AO31x2_ASAP7_75t_L g1553 ( 
.A1(n_1355),
.A2(n_1284),
.A3(n_1296),
.B(n_1253),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_L g1554 ( 
.A(n_1265),
.B(n_1151),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1375),
.A2(n_1377),
.B1(n_915),
.B2(n_936),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1365),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1295),
.B(n_1241),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1372),
.A2(n_1389),
.B(n_1380),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1331),
.A2(n_1328),
.B(n_1355),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1383),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1527),
.A2(n_1547),
.B(n_1534),
.C(n_1523),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1442),
.B(n_1419),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1521),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1427),
.A2(n_1504),
.B(n_1495),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1526),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1519),
.A2(n_1555),
.B(n_1432),
.C(n_1533),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1477),
.B(n_1444),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1423),
.B(n_1440),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1539),
.A2(n_1544),
.B1(n_1445),
.B2(n_1422),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1428),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1539),
.A2(n_1544),
.B1(n_1445),
.B2(n_1430),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1465),
.B(n_1474),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1533),
.A2(n_1543),
.B(n_1528),
.C(n_1475),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1475),
.A2(n_1483),
.B(n_1448),
.C(n_1450),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1483),
.A2(n_1448),
.B(n_1452),
.C(n_1501),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1476),
.A2(n_1501),
.B1(n_1458),
.B2(n_1499),
.C(n_1461),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1484),
.B(n_1515),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1456),
.A2(n_1437),
.B1(n_1525),
.B2(n_1550),
.Y(n_1581)
);

O2A1O1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1494),
.A2(n_1561),
.B(n_1540),
.C(n_1535),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1451),
.B(n_1502),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1507),
.A2(n_1509),
.B(n_1508),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1462),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1507),
.A2(n_1508),
.B(n_1509),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1464),
.B(n_1563),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1456),
.A2(n_1446),
.B1(n_1471),
.B2(n_1460),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1493),
.A2(n_1517),
.B(n_1560),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1467),
.B(n_1513),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1454),
.Y(n_1591)
);

OAI31xp33_ASAP7_75t_L g1592 ( 
.A1(n_1535),
.A2(n_1536),
.A3(n_1560),
.B(n_1517),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1425),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1446),
.A2(n_1471),
.B1(n_1517),
.B2(n_1560),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1480),
.A2(n_1545),
.B(n_1551),
.C(n_1455),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1466),
.A2(n_1463),
.B(n_1471),
.C(n_1485),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1417),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1491),
.B(n_1429),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1491),
.B(n_1503),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1485),
.A2(n_1500),
.B1(n_1469),
.B2(n_1436),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1463),
.A2(n_1485),
.B(n_1497),
.C(n_1472),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1512),
.B(n_1518),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1497),
.A2(n_1472),
.B(n_1453),
.C(n_1489),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1496),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1538),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1441),
.B(n_1487),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1510),
.A2(n_1524),
.B(n_1559),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1520),
.A2(n_1526),
.B1(n_1492),
.B2(n_1420),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1497),
.A2(n_1506),
.B(n_1505),
.C(n_1459),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1541),
.B(n_1562),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1425),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1549),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1470),
.A2(n_1554),
.B(n_1479),
.C(n_1520),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1510),
.A2(n_1556),
.B(n_1559),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1492),
.A2(n_1416),
.B1(n_1420),
.B2(n_1530),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1511),
.A2(n_1531),
.B(n_1552),
.C(n_1421),
.Y(n_1616)
);

O2A1O1Ixp5_ASAP7_75t_L g1617 ( 
.A1(n_1418),
.A2(n_1548),
.B(n_1421),
.C(n_1531),
.Y(n_1617)
);

BUFx4_ASAP7_75t_R g1618 ( 
.A(n_1498),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1482),
.A2(n_1433),
.B1(n_1511),
.B2(n_1443),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1488),
.B(n_1481),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1433),
.B(n_1470),
.Y(n_1621)
);

OAI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1548),
.A2(n_1552),
.A3(n_1486),
.B(n_1457),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1498),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1443),
.A2(n_1468),
.B1(n_1537),
.B2(n_1522),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1468),
.A2(n_1532),
.B(n_1522),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1435),
.B(n_1486),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1490),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1516),
.A2(n_1522),
.B1(n_1532),
.B2(n_1537),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1490),
.B(n_1478),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1486),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1529),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1516),
.A2(n_1532),
.B1(n_1537),
.B2(n_1438),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1516),
.A2(n_1457),
.B(n_1479),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1424),
.A2(n_1558),
.B(n_1557),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1529),
.A2(n_1553),
.B1(n_1439),
.B2(n_1431),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1449),
.B(n_1553),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1449),
.B(n_1447),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1514),
.A2(n_1542),
.B1(n_1546),
.B2(n_1556),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1426),
.B(n_1477),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1477),
.B(n_1444),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1475),
.A2(n_1388),
.B(n_1368),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1515),
.B(n_1473),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1527),
.A2(n_943),
.B(n_1547),
.C(n_1534),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1465),
.B(n_1474),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1523),
.A2(n_1412),
.B(n_1555),
.C(n_1519),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1527),
.A2(n_1201),
.B1(n_1547),
.B2(n_1534),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1521),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1527),
.A2(n_1201),
.B1(n_1547),
.B2(n_1534),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1475),
.A2(n_1388),
.B(n_1368),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1475),
.A2(n_1388),
.B(n_1368),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1527),
.A2(n_943),
.B(n_1547),
.C(n_1534),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1533),
.A2(n_1388),
.B(n_1368),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1442),
.B(n_1419),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1442),
.B(n_1419),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1533),
.A2(n_1388),
.B(n_1368),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1527),
.A2(n_943),
.B(n_1547),
.C(n_1534),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1434),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1521),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1515),
.B(n_1473),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1442),
.B(n_1419),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1527),
.A2(n_1201),
.B1(n_1547),
.B2(n_1534),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1434),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1425),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1526),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1434),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1477),
.B(n_1444),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1566),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1583),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1583),
.B(n_1626),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1639),
.B(n_1636),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1659),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1591),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1629),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1646),
.A2(n_1661),
.B1(n_1648),
.B2(n_1572),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1641),
.B(n_1649),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1620),
.B(n_1627),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1631),
.B(n_1567),
.Y(n_1677)
);

BUFx12f_ASAP7_75t_L g1678 ( 
.A(n_1593),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1647),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1650),
.B(n_1601),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1658),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1567),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1565),
.B(n_1653),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1596),
.B(n_1620),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1632),
.A2(n_1628),
.B(n_1633),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1584),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1657),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1621),
.Y(n_1689)
);

AO21x2_ASAP7_75t_L g1690 ( 
.A1(n_1624),
.A2(n_1637),
.B(n_1574),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1662),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1594),
.B(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1665),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1594),
.B(n_1622),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1597),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1652),
.A2(n_1655),
.B(n_1569),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1588),
.B(n_1599),
.Y(n_1697)
);

BUFx2_ASAP7_75t_SL g1698 ( 
.A(n_1600),
.Y(n_1698)
);

OR2x6_ASAP7_75t_L g1699 ( 
.A(n_1625),
.B(n_1603),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1605),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1624),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1637),
.A2(n_1574),
.B(n_1572),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1584),
.B(n_1586),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1570),
.B(n_1640),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1654),
.B(n_1660),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1599),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1575),
.B(n_1644),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1581),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1602),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1575),
.B(n_1644),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1617),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1600),
.B(n_1607),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1607),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1609),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1581),
.B(n_1580),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1614),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1616),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1634),
.B(n_1606),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1578),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1672),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_SL g1721 ( 
.A(n_1681),
.B(n_1619),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1683),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1580),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1672),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1689),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1675),
.A2(n_1648),
.B1(n_1661),
.B2(n_1646),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1684),
.B(n_1585),
.Y(n_1727)
);

OAI33xp33_ASAP7_75t_L g1728 ( 
.A1(n_1707),
.A2(n_1710),
.A3(n_1715),
.B1(n_1719),
.B2(n_1697),
.B3(n_1645),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1675),
.A2(n_1577),
.B(n_1582),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1718),
.B(n_1587),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1718),
.B(n_1638),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1718),
.B(n_1670),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1670),
.B(n_1638),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1712),
.B(n_1573),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1671),
.B(n_1590),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1579),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1673),
.B(n_1613),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1689),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_SL g1739 ( 
.A(n_1681),
.B(n_1619),
.Y(n_1739)
);

BUFx4f_ASAP7_75t_L g1740 ( 
.A(n_1675),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1689),
.Y(n_1741)
);

OAI211xp5_ASAP7_75t_L g1742 ( 
.A1(n_1674),
.A2(n_1564),
.B(n_1576),
.C(n_1643),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1712),
.B(n_1598),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1715),
.B(n_1571),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1668),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1708),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1705),
.B(n_1635),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1674),
.A2(n_1656),
.B1(n_1651),
.B2(n_1589),
.Y(n_1748)
);

NOR4xp25_ASAP7_75t_SL g1749 ( 
.A(n_1717),
.B(n_1611),
.C(n_1663),
.D(n_1618),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1669),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1604),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1676),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1741),
.Y(n_1753)
);

AO21x2_ASAP7_75t_L g1754 ( 
.A1(n_1722),
.A2(n_1686),
.B(n_1711),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1736),
.A2(n_1702),
.B1(n_1694),
.B2(n_1681),
.Y(n_1755)
);

OAI31xp33_ASAP7_75t_L g1756 ( 
.A1(n_1742),
.A2(n_1701),
.A3(n_1719),
.B(n_1694),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1720),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1728),
.A2(n_1701),
.B1(n_1707),
.B2(n_1710),
.C(n_1694),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1736),
.A2(n_1702),
.B1(n_1681),
.B2(n_1697),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1726),
.A2(n_1681),
.B1(n_1696),
.B2(n_1697),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1726),
.A2(n_1681),
.B1(n_1696),
.B2(n_1699),
.Y(n_1762)
);

AOI31xp33_ASAP7_75t_L g1763 ( 
.A1(n_1728),
.A2(n_1615),
.A3(n_1608),
.B(n_1623),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1724),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1738),
.Y(n_1766)
);

AOI33xp33_ASAP7_75t_L g1767 ( 
.A1(n_1736),
.A2(n_1692),
.A3(n_1704),
.B1(n_1706),
.B2(n_1691),
.B3(n_1693),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_L g1768 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1768)
);

OAI321xp33_ASAP7_75t_L g1769 ( 
.A1(n_1748),
.A2(n_1685),
.A3(n_1680),
.B1(n_1699),
.B2(n_1692),
.C(n_1714),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1745),
.B(n_1667),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1747),
.A2(n_1702),
.B1(n_1690),
.B2(n_1692),
.C(n_1680),
.Y(n_1771)
);

OAI31xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1742),
.A2(n_1746),
.A3(n_1748),
.B(n_1731),
.Y(n_1772)
);

OAI31xp33_ASAP7_75t_L g1773 ( 
.A1(n_1747),
.A2(n_1592),
.A3(n_1680),
.B(n_1714),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1738),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1725),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1732),
.B(n_1706),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

CKINVDCx11_ASAP7_75t_R g1778 ( 
.A(n_1752),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1729),
.A2(n_1698),
.B1(n_1699),
.B2(n_1685),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1746),
.A2(n_1740),
.B1(n_1745),
.B2(n_1744),
.Y(n_1780)
);

OAI33xp33_ASAP7_75t_L g1781 ( 
.A1(n_1727),
.A2(n_1709),
.A3(n_1669),
.B1(n_1693),
.B2(n_1688),
.B3(n_1691),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1732),
.B(n_1706),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1679),
.C(n_1682),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1734),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1749),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1731),
.A2(n_1702),
.B1(n_1690),
.B2(n_1723),
.C(n_1727),
.Y(n_1786)
);

AND2x6_ASAP7_75t_SL g1787 ( 
.A(n_1723),
.B(n_1568),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1731),
.A2(n_1690),
.B1(n_1677),
.B2(n_1695),
.C(n_1700),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1735),
.B(n_1678),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1776),
.B(n_1732),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1778),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1754),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1776),
.B(n_1733),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1757),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1758),
.Y(n_1796)
);

CKINVDCx8_ASAP7_75t_R g1797 ( 
.A(n_1787),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1768),
.A2(n_1687),
.B(n_1703),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1754),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1772),
.B(n_1756),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1782),
.B(n_1733),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1765),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1783),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1771),
.A2(n_1713),
.B(n_1716),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1753),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1775),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1772),
.A2(n_1769),
.B(n_1756),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1733),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1734),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1775),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1784),
.B(n_1743),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1764),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1783),
.B(n_1690),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1768),
.A2(n_1687),
.B(n_1703),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1788),
.B(n_1769),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1750),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1794),
.B(n_1767),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1791),
.B(n_1797),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1815),
.B(n_1721),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1798),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1794),
.B(n_1775),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1794),
.B(n_1730),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1803),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1798),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1807),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1802),
.B(n_1730),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1806),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1804),
.B(n_1770),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1804),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1791),
.B(n_1789),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1803),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1815),
.B(n_1721),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1802),
.B(n_1809),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1803),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1801),
.B(n_1750),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1808),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1808),
.B(n_1759),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1809),
.B(n_1763),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1792),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_SL g1843 ( 
.A(n_1818),
.B(n_1785),
.C(n_1615),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1809),
.B(n_1730),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1792),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1790),
.B(n_1739),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1818),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1807),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1797),
.B(n_1678),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1805),
.B(n_1760),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1795),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1806),
.Y(n_1852)
);

OAI21xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1797),
.A2(n_1773),
.B(n_1761),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1817),
.A2(n_1773),
.B(n_1755),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1814),
.B(n_1735),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1805),
.B(n_1766),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1814),
.B(n_1774),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1795),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1807),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_SL g1860 ( 
.A(n_1811),
.B(n_1785),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1805),
.B(n_1743),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1798),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1817),
.A2(n_1779),
.B(n_1780),
.C(n_1737),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1831),
.B(n_1805),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1838),
.B(n_1811),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1820),
.B(n_1678),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1842),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1831),
.B(n_1805),
.Y(n_1869)
);

NAND2x2_ASAP7_75t_L g1870 ( 
.A(n_1837),
.B(n_1664),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1835),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1822),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1823),
.B(n_1790),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1823),
.B(n_1811),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1838),
.B(n_1805),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1855),
.B(n_1796),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1825),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1842),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1854),
.A2(n_1812),
.B1(n_1762),
.B2(n_1690),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1845),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1845),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1839),
.B(n_1813),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1851),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1837),
.B(n_1813),
.Y(n_1884)
);

A2O1A1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1853),
.A2(n_1812),
.B(n_1816),
.C(n_1698),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1853),
.A2(n_1781),
.B(n_1799),
.C(n_1800),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1851),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1821),
.B(n_1834),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1819),
.B(n_1824),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1819),
.B(n_1813),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1829),
.B(n_1810),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1858),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1824),
.B(n_1810),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1832),
.Y(n_1894)
);

NAND2xp33_ASAP7_75t_L g1895 ( 
.A(n_1843),
.B(n_1608),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1859),
.B(n_1739),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1858),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1828),
.B(n_1810),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1850),
.A2(n_1847),
.B1(n_1861),
.B2(n_1821),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1822),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1852),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1825),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1873),
.B(n_1859),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1894),
.B(n_1840),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1864),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1864),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1875),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1865),
.Y(n_1909)
);

INVx3_ASAP7_75t_SL g1910 ( 
.A(n_1865),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1866),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1873),
.B(n_1828),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1869),
.Y(n_1913)
);

CKINVDCx16_ASAP7_75t_R g1914 ( 
.A(n_1874),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1874),
.B(n_1844),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1877),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1902),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1882),
.B(n_1830),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1868),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1895),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1895),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1885),
.B(n_1849),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1876),
.B(n_1830),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1876),
.B(n_1855),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1889),
.B(n_1844),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1889),
.B(n_1846),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1901),
.B(n_1841),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1878),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_1884),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1871),
.B(n_1848),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1903),
.B(n_1871),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1910),
.A2(n_1885),
.B(n_1856),
.C(n_1886),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1904),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1920),
.A2(n_1899),
.B1(n_1879),
.B2(n_1872),
.C(n_1900),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1904),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1916),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1916),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1914),
.B(n_1867),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1921),
.A2(n_1860),
.B1(n_1821),
.B2(n_1834),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1923),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1910),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1914),
.B(n_1867),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1923),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1905),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1903),
.B(n_1890),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1906),
.Y(n_1946)
);

OAI21xp33_ASAP7_75t_L g1947 ( 
.A1(n_1922),
.A2(n_1891),
.B(n_1890),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1924),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1910),
.B(n_1827),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1908),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1924),
.Y(n_1951)
);

OAI21xp33_ASAP7_75t_SL g1952 ( 
.A1(n_1922),
.A2(n_1898),
.B(n_1893),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1909),
.A2(n_1863),
.B(n_1834),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1945),
.B(n_1931),
.Y(n_1954)
);

OAI21xp33_ASAP7_75t_SL g1955 ( 
.A1(n_1949),
.A2(n_1925),
.B(n_1926),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1946),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

NAND2x1_ASAP7_75t_L g1958 ( 
.A(n_1931),
.B(n_1827),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1938),
.B(n_1929),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1948),
.B(n_1918),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1941),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1941),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1944),
.B(n_1918),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1951),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1944),
.B(n_1925),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1942),
.B(n_1915),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1940),
.B(n_1915),
.Y(n_1967)
);

OAI21xp33_ASAP7_75t_L g1968 ( 
.A1(n_1952),
.A2(n_1927),
.B(n_1930),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1959),
.B(n_1911),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1966),
.B(n_1943),
.Y(n_1970)
);

NAND3xp33_ASAP7_75t_L g1971 ( 
.A(n_1961),
.B(n_1932),
.C(n_1949),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1962),
.B(n_1947),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1963),
.A2(n_1953),
.B1(n_1939),
.B2(n_1870),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1968),
.A2(n_1950),
.B(n_1908),
.C(n_1936),
.Y(n_1974)
);

OAI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1956),
.A2(n_1934),
.B1(n_1950),
.B2(n_1908),
.C(n_1907),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1955),
.B(n_1954),
.Y(n_1976)
);

OAI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1957),
.A2(n_1907),
.B1(n_1906),
.B2(n_1913),
.C(n_1962),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1960),
.B(n_1926),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1964),
.B(n_1965),
.C(n_1967),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1958),
.Y(n_1980)
);

O2A1O1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1975),
.A2(n_1972),
.B(n_1974),
.C(n_1977),
.Y(n_1981)
);

OAI211xp5_ASAP7_75t_L g1982 ( 
.A1(n_1971),
.A2(n_1937),
.B(n_1935),
.C(n_1933),
.Y(n_1982)
);

AOI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1979),
.A2(n_1906),
.B1(n_1907),
.B2(n_1913),
.C(n_1928),
.Y(n_1983)
);

OAI31xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1973),
.A2(n_1913),
.A3(n_1919),
.B(n_1928),
.Y(n_1984)
);

OAI322xp33_ASAP7_75t_L g1985 ( 
.A1(n_1969),
.A2(n_1976),
.A3(n_1973),
.B1(n_1980),
.B2(n_1978),
.C1(n_1919),
.C2(n_1970),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1975),
.A2(n_1917),
.B1(n_1872),
.B2(n_1900),
.C(n_1826),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1978),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1987),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1982),
.Y(n_1989)
);

NOR2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1985),
.B(n_1917),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1981),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1983),
.B(n_1827),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1986),
.Y(n_1993)
);

INVx1_ASAP7_75t_SL g1994 ( 
.A(n_1984),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1987),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1994),
.A2(n_1912),
.B(n_1896),
.Y(n_1996)
);

OAI211xp5_ASAP7_75t_L g1997 ( 
.A1(n_1989),
.A2(n_1827),
.B(n_1912),
.C(n_1897),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1991),
.A2(n_1988),
.B(n_1992),
.Y(n_1998)
);

AOI211xp5_ASAP7_75t_L g1999 ( 
.A1(n_1995),
.A2(n_1883),
.B(n_1880),
.C(n_1881),
.Y(n_1999)
);

NAND4xp75_ASAP7_75t_L g2000 ( 
.A(n_1990),
.B(n_1892),
.C(n_1887),
.D(n_1893),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1993),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1998),
.B(n_1896),
.Y(n_2002)
);

NAND3xp33_ASAP7_75t_SL g2003 ( 
.A(n_1996),
.B(n_2001),
.C(n_1993),
.Y(n_2003)
);

AND3x4_ASAP7_75t_L g2004 ( 
.A(n_2000),
.B(n_1997),
.C(n_1999),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1996),
.B(n_1888),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2003),
.Y(n_2006)
);

NOR2x1p5_ASAP7_75t_L g2007 ( 
.A(n_2002),
.B(n_1857),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_2006),
.A2(n_2005),
.B1(n_2007),
.B2(n_2004),
.Y(n_2008)
);

AOI322xp5_ASAP7_75t_L g2009 ( 
.A1(n_2006),
.A2(n_1834),
.A3(n_1821),
.B1(n_1826),
.B2(n_1862),
.C1(n_1793),
.C2(n_1800),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_2008),
.A2(n_1870),
.B1(n_1888),
.B2(n_1862),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_2009),
.A2(n_1888),
.B1(n_1896),
.B2(n_1898),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_2010),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_2011),
.A2(n_1888),
.B1(n_1800),
.B2(n_1793),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_2013),
.A2(n_1857),
.B1(n_1836),
.B2(n_1833),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2012),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_SL g2016 ( 
.A1(n_2015),
.A2(n_1612),
.B1(n_1836),
.B2(n_1833),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_2016),
.B(n_2014),
.C(n_1799),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2017),
.B(n_1793),
.Y(n_2018)
);

XNOR2xp5_ASAP7_75t_L g2019 ( 
.A(n_2018),
.B(n_1749),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2019),
.A2(n_1846),
.B1(n_1793),
.B2(n_1799),
.Y(n_2020)
);

AOI211xp5_ASAP7_75t_L g2021 ( 
.A1(n_2020),
.A2(n_1595),
.B(n_1800),
.C(n_1799),
.Y(n_2021)
);


endmodule