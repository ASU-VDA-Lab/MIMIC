module fake_netlist_1_10288_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_3), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g13 ( .A1(n_9), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_10), .B(n_4), .Y(n_14) );
NOR2x1_ASAP7_75t_L g15 ( .A(n_12), .B(n_7), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_11), .B(n_9), .Y(n_16) );
AOI22xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_13), .B1(n_15), .B2(n_5), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_6), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_17), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NOR3xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .C(n_19), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_22), .Y(n_25) );
INVx3_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
endmodule