module fake_jpeg_31939_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_53),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_45),
.B1(n_71),
.B2(n_69),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_51),
.B1(n_46),
.B2(n_45),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_46),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_57),
.B1(n_64),
.B2(n_62),
.Y(n_89)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_91),
.Y(n_125)
);

OAI22x1_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_58),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_103),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_61),
.B1(n_59),
.B2(n_58),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_3),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_35),
.B(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_16),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_29),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_34),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_38),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_126),
.B1(n_123),
.B2(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_132),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_153),
.A2(n_130),
.B1(n_133),
.B2(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_129),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.C(n_135),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_146),
.C(n_135),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_150),
.B(n_151),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_149),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_148),
.Y(n_163)
);

XNOR2x2_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_143),
.Y(n_164)
);


endmodule