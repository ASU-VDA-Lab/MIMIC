module real_jpeg_29307_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_0),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_36),
.B1(n_92),
.B2(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_22),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_42),
.B(n_90),
.C(n_92),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_1),
.B(n_29),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_1),
.A2(n_29),
.B(n_59),
.C(n_68),
.D(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_26),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_51),
.B(n_134),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_1),
.A2(n_22),
.B(n_32),
.C(n_74),
.D(n_164),
.Y(n_163)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_3),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_66),
.Y(n_133)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_10),
.B(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_47),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_116),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_114),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_80),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_18),
.B(n_80),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_57),
.C(n_71),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_19),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_38),
.C(n_44),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_31),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_22),
.A2(n_41),
.B(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_29),
.A3(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_25),
.B(n_35),
.Y(n_164)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_32),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_28),
.B(n_30),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_28),
.A2(n_46),
.A3(n_61),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_29),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_40),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_40),
.B(n_103),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_41),
.A2(n_42),
.B1(n_92),
.B2(n_93),
.Y(n_99)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_46),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_51),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_52),
.A2(n_140),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_56),
.B(n_135),
.Y(n_134)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_57),
.B(n_71),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_67),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_59),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_70),
.A2(n_112),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_70),
.B(n_91),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_72),
.B(n_76),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_79),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_96),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_154),
.Y(n_153)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_169),
.B(n_173),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_159),
.B(n_168),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_136),
.B(n_158),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_124),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_130),
.C(n_132),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_145),
.B(n_157),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_156),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_161),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);


endmodule