module fake_jpeg_7369_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_32),
.B1(n_18),
.B2(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_19),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_18),
.B1(n_33),
.B2(n_22),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_23),
.B1(n_17),
.B2(n_27),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_63),
.B1(n_67),
.B2(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_63)
);

NAND2xp67_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_16),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_27),
.B1(n_17),
.B2(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_28),
.B1(n_16),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_16),
.B1(n_31),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_31),
.B1(n_34),
.B2(n_21),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_77),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_80),
.B(n_83),
.Y(n_142)
);

BUFx12f_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_92),
.B1(n_100),
.B2(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_11),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_102),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_11),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_15),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_59),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_48),
.A2(n_21),
.B(n_25),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_112),
.B(n_21),
.Y(n_130)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_0),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_131),
.B(n_106),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_53),
.B1(n_70),
.B2(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_122),
.B1(n_100),
.B2(n_92),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_50),
.B1(n_51),
.B2(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_125),
.B1(n_127),
.B2(n_98),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_70),
.B1(n_54),
.B2(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_54),
.B1(n_49),
.B2(n_45),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_45),
.C(n_54),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_132),
.C(n_108),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_49),
.B1(n_34),
.B2(n_31),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_141),
.B(n_118),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_0),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_65),
.C(n_25),
.Y(n_132)
);

OAI22x1_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_95),
.B1(n_104),
.B2(n_110),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_151),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_153),
.B(n_166),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_86),
.B1(n_88),
.B2(n_111),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_173),
.B1(n_175),
.B2(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_105),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_99),
.B(n_82),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_160),
.B(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_87),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_164),
.C(n_113),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_82),
.C(n_93),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_78),
.B(n_77),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_171),
.B(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_75),
.B1(n_109),
.B2(n_80),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_96),
.B1(n_89),
.B2(n_98),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_94),
.B1(n_101),
.B2(n_14),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_101),
.B(n_1),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_138),
.B1(n_137),
.B2(n_3),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_14),
.B1(n_12),
.B2(n_3),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_117),
.C(n_115),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_115),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_115),
.B1(n_131),
.B2(n_113),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_153),
.B1(n_174),
.B2(n_145),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_131),
.B(n_113),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_189),
.B(n_198),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_131),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_209),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_117),
.B(n_139),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_140),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_168),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_208),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_139),
.B(n_138),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_137),
.B(n_140),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_0),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_1),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_224),
.B(n_234),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_146),
.B(n_159),
.C(n_171),
.D(n_174),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_228),
.Y(n_250)
);

AO32x1_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_174),
.A3(n_156),
.B1(n_143),
.B2(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_156),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_169),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_179),
.C(n_185),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_163),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_178),
.B(n_6),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_172),
.B1(n_175),
.B2(n_173),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_231),
.Y(n_252)
);

XNOR2x2_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_4),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_236),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_236),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_4),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_4),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_5),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_251),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_203),
.B1(n_177),
.B2(n_197),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_230),
.B1(n_232),
.B2(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_194),
.C(n_182),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_247),
.C(n_253),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_206),
.B1(n_203),
.B2(n_195),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_249),
.B1(n_256),
.B2(n_224),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_200),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_180),
.B1(n_178),
.B2(n_183),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_186),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_208),
.C(n_188),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_234),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_220),
.C(n_222),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_221),
.A2(n_178),
.B1(n_209),
.B2(n_7),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_226),
.B(n_210),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_275),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_257),
.B1(n_249),
.B2(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_274),
.Y(n_292)
);

AO21x2_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_230),
.B(n_219),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_257),
.B(n_248),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_233),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_276),
.C(n_279),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_256),
.B1(n_259),
.B2(n_9),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_226),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_222),
.C(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_226),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_5),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_6),
.C(n_7),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_7),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_280),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_252),
.B1(n_238),
.B2(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_271),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_265),
.C(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_290),
.C(n_263),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_291),
.B(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_253),
.C(n_255),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_238),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_268),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_267),
.B1(n_8),
.B2(n_9),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_305),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_279),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_266),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_275),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_306),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_292),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_270),
.B(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_7),
.C(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_8),
.C(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_295),
.C(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_316),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

INVx11_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_297),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_314),
.C(n_317),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_283),
.B(n_308),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_315),
.B(n_319),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_299),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_320),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_330),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_325),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_325),
.Y(n_336)
);


endmodule