module fake_netlist_6_330_n_756 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_756);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_756;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_703;
wire n_578;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_611;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_0),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_45),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_53),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_30),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_82),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_59),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_91),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_47),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_84),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_50),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_35),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_124),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_32),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_61),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_95),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_73),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g193 ( 
.A(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_36),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_31),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_123),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_131),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_29),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_62),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_40),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_2),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_19),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_4),
.B(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_6),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_7),
.B(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_7),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_9),
.B(n_10),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

CKINVDCx8_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_9),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_20),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_10),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_11),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_167),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_206),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_R g255 ( 
.A(n_158),
.B(n_12),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_13),
.Y(n_256)
);

BUFx6f_ASAP7_75t_SL g257 ( 
.A(n_219),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_167),
.B1(n_179),
.B2(n_186),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_159),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_186),
.B1(n_179),
.B2(n_171),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g271 ( 
.A1(n_228),
.A2(n_213),
.B(n_171),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_162),
.Y(n_273)
);

AO21x2_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_208),
.B(n_207),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_168),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_169),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_170),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_174),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_205),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_242),
.B(n_238),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_215),
.B(n_176),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_220),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_178),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_242),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_185),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_218),
.B(n_204),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_214),
.B1(n_216),
.B2(n_226),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_190),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_222),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_224),
.B(n_202),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_238),
.A2(n_201),
.B1(n_200),
.B2(n_197),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_233),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_282),
.B(n_242),
.Y(n_307)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_239),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_220),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_277),
.B(n_231),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_245),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_230),
.B1(n_225),
.B2(n_247),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_265),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_263),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_253),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_273),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_271),
.B(n_248),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_274),
.A2(n_230),
.B1(n_225),
.B2(n_256),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_254),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_288),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_274),
.A2(n_230),
.B1(n_225),
.B2(n_251),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_243),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_243),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_243),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_243),
.Y(n_332)
);

OAI221xp5_ASAP7_75t_L g333 ( 
.A1(n_271),
.A2(n_252),
.B1(n_251),
.B2(n_246),
.C(n_241),
.Y(n_333)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_276),
.B(n_299),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_267),
.B(n_241),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_258),
.B(n_246),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_260),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_261),
.B(n_231),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_298),
.B(n_191),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_252),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_258),
.B(n_21),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_258),
.B(n_22),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_14),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_L g355 ( 
.A(n_258),
.B(n_255),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_276),
.B(n_24),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_261),
.B(n_255),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_284),
.B(n_15),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_279),
.B(n_15),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_25),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_26),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_280),
.B(n_16),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_290),
.B(n_16),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_284),
.B(n_289),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_319),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_270),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_291),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_293),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_291),
.B(n_296),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_330),
.A2(n_296),
.B(n_305),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_270),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_296),
.B(n_305),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_270),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_297),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_270),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_297),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_305),
.B(n_297),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_297),
.B(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_302),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_281),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_361),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_351),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_310),
.A2(n_257),
.B1(n_262),
.B2(n_302),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

OR2x6_ASAP7_75t_SL g395 ( 
.A(n_358),
.B(n_289),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_334),
.B(n_275),
.Y(n_396)
);

O2A1O1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_355),
.A2(n_268),
.B(n_266),
.C(n_285),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_343),
.A2(n_257),
.B1(n_262),
.B2(n_268),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_285),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_317),
.A2(n_292),
.B(n_266),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_323),
.B(n_344),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_311),
.B(n_27),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_338),
.A2(n_292),
.B(n_28),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_354),
.A2(n_292),
.B(n_17),
.C(n_34),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_337),
.A2(n_292),
.B(n_33),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_37),
.Y(n_407)
);

O2A1O1Ixp5_ASAP7_75t_L g408 ( 
.A1(n_321),
.A2(n_94),
.B(n_38),
.C(n_39),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_368),
.B(n_17),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_333),
.A2(n_155),
.B1(n_42),
.B2(n_43),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_41),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_307),
.B(n_44),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_321),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_51),
.B(n_52),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_363),
.A2(n_55),
.B(n_56),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_341),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_364),
.A2(n_348),
.B(n_352),
.Y(n_417)
);

O2A1O1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_354),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_362),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_312),
.B(n_66),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_67),
.C(n_68),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_69),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_340),
.A2(n_70),
.B(n_74),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_366),
.B(n_75),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_366),
.B(n_76),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_320),
.B(n_77),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_309),
.B(n_78),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_329),
.B(n_342),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_79),
.Y(n_433)
);

AOI221xp5_ASAP7_75t_L g434 ( 
.A1(n_314),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.C(n_88),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_314),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_370),
.A2(n_93),
.B(n_96),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_336),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_345),
.A2(n_97),
.B(n_100),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_438),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

AO21x1_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_322),
.B(n_346),
.Y(n_443)
);

AO31x2_ASAP7_75t_L g444 ( 
.A1(n_393),
.A2(n_322),
.A3(n_346),
.B(n_345),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_376),
.B(n_325),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_416),
.Y(n_447)
);

OAI22x1_ASAP7_75t_L g448 ( 
.A1(n_372),
.A2(n_325),
.B1(n_308),
.B2(n_356),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_381),
.A2(n_356),
.B(n_308),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g450 ( 
.A1(n_390),
.A2(n_373),
.B(n_433),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_378),
.A2(n_101),
.B(n_102),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_377),
.A2(n_154),
.B(n_105),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_387),
.A2(n_103),
.B(n_106),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

AOI221x1_ASAP7_75t_L g455 ( 
.A1(n_393),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.C(n_112),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_391),
.B(n_113),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_374),
.B(n_114),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_388),
.A2(n_152),
.B(n_118),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_399),
.A2(n_383),
.B(n_386),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_374),
.A2(n_117),
.B(n_121),
.Y(n_460)
);

NOR4xp25_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_404),
.C(n_422),
.D(n_418),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_401),
.A2(n_122),
.B(n_125),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_392),
.B(n_126),
.Y(n_464)
);

AOI221x1_ASAP7_75t_L g465 ( 
.A1(n_410),
.A2(n_417),
.B1(n_398),
.B2(n_424),
.C(n_400),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_411),
.A2(n_127),
.B(n_128),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_130),
.C(n_132),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_389),
.A2(n_134),
.B(n_135),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_434),
.A2(n_136),
.B(n_137),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

AOI221xp5_ASAP7_75t_L g474 ( 
.A1(n_410),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.C(n_142),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_382),
.B(n_145),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_397),
.A2(n_148),
.B(n_149),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_396),
.A2(n_151),
.B(n_432),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_436),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_405),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_420),
.A2(n_439),
.B(n_423),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

A2O1A1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_379),
.A2(n_435),
.B(n_413),
.C(n_408),
.Y(n_483)
);

NOR2x1_ASAP7_75t_R g484 ( 
.A(n_412),
.B(n_375),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

NAND2x1p5_ASAP7_75t_L g486 ( 
.A(n_402),
.B(n_429),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_398),
.A2(n_415),
.B(n_414),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_426),
.A2(n_431),
.B(n_403),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_395),
.B(n_419),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_406),
.A2(n_427),
.B(n_440),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_437),
.A2(n_381),
.B(n_377),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_391),
.Y(n_492)
);

AO31x2_ASAP7_75t_L g493 ( 
.A1(n_393),
.A2(n_354),
.A3(n_404),
.B(n_410),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_374),
.A2(n_258),
.B(n_399),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_449),
.A2(n_481),
.B(n_491),
.Y(n_495)
);

OAI21x1_ASAP7_75t_SL g496 ( 
.A1(n_462),
.A2(n_478),
.B(n_456),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_492),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_443),
.B(n_459),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_447),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_494),
.A2(n_452),
.B(n_477),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_470),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_446),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_445),
.A2(n_457),
.B(n_483),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_487),
.A2(n_455),
.B(n_458),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_464),
.A2(n_490),
.B(n_466),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_488),
.A2(n_482),
.B(n_485),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_460),
.A2(n_486),
.B(n_451),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_450),
.A2(n_472),
.B1(n_474),
.B2(n_485),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_482),
.A2(n_473),
.B(n_475),
.Y(n_512)
);

AO21x2_ASAP7_75t_L g513 ( 
.A1(n_461),
.A2(n_476),
.B(n_467),
.Y(n_513)
);

BUFx8_ASAP7_75t_SL g514 ( 
.A(n_469),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_442),
.B(n_446),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_442),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_471),
.A2(n_451),
.B(n_453),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_448),
.A2(n_453),
.B(n_489),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_446),
.B(n_479),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_454),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

NOR2x1_ASAP7_75t_SL g523 ( 
.A(n_454),
.B(n_484),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_493),
.Y(n_524)
);

BUFx2_ASAP7_75t_SL g525 ( 
.A(n_454),
.Y(n_525)
);

INVx4_ASAP7_75t_SL g526 ( 
.A(n_493),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_493),
.A2(n_450),
.B(n_445),
.C(n_483),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_480),
.B(n_372),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_446),
.Y(n_529)
);

AO31x2_ASAP7_75t_L g530 ( 
.A1(n_443),
.A2(n_465),
.A3(n_448),
.B(n_483),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_445),
.A2(n_263),
.B1(n_259),
.B2(n_483),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_449),
.A2(n_481),
.B(n_381),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_445),
.B(n_376),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_454),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_450),
.A2(n_487),
.B(n_483),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_502),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_531),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_504),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_515),
.Y(n_543)
);

AO21x2_ASAP7_75t_L g544 ( 
.A1(n_527),
.A2(n_505),
.B(n_500),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_537),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_524),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_531),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

INVx3_ASAP7_75t_SL g549 ( 
.A(n_499),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_503),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_515),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_527),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_529),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_529),
.Y(n_559)
);

AO21x2_ASAP7_75t_L g560 ( 
.A1(n_505),
.A2(n_517),
.B(n_535),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_496),
.A2(n_510),
.B(n_508),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_523),
.B(n_534),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_526),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_535),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_497),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_532),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_530),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_519),
.B(n_525),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_516),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_516),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_530),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_530),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_540),
.B(n_498),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_557),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_498),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_566),
.Y(n_579)
);

AOI221xp5_ASAP7_75t_L g580 ( 
.A1(n_551),
.A2(n_510),
.B1(n_513),
.B2(n_499),
.C(n_536),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_546),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_538),
.B(n_547),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_541),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_557),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_513),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_558),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_550),
.Y(n_588)
);

AOI221xp5_ASAP7_75t_L g589 ( 
.A1(n_547),
.A2(n_536),
.B1(n_520),
.B2(n_506),
.C(n_514),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_550),
.Y(n_591)
);

NOR2x1_ASAP7_75t_SL g592 ( 
.A(n_565),
.B(n_563),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_506),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_552),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_556),
.Y(n_596)
);

BUFx2_ASAP7_75t_SL g597 ( 
.A(n_562),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_554),
.B(n_520),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_562),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_565),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_539),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_562),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_559),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_568),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_545),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_545),
.B(n_509),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_564),
.B(n_509),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_564),
.B(n_495),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_568),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

AO31x2_ASAP7_75t_L g612 ( 
.A1(n_561),
.A2(n_507),
.A3(n_574),
.B(n_573),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_542),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_570),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_549),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_542),
.B(n_571),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_574),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_569),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_605),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_575),
.B(n_560),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_544),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_605),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_602),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_583),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_593),
.B(n_544),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_575),
.B(n_560),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_544),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_610),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_600),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_582),
.B(n_549),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_604),
.B(n_580),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_581),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_594),
.B(n_548),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_611),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_606),
.B(n_549),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_594),
.B(n_567),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_594),
.B(n_567),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_615),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_581),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_594),
.B(n_595),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_598),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_606),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_622),
.B(n_608),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_608),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_641),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_620),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_601),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_620),
.Y(n_655)
);

AND2x4_ASAP7_75t_SL g656 ( 
.A(n_627),
.B(n_586),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_601),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_623),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_628),
.B(n_609),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_624),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_635),
.B(n_596),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_623),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_637),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_609),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_631),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_612),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_630),
.B(n_607),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_637),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_621),
.B(n_612),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_637),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_633),
.B(n_647),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_644),
.A2(n_589),
.B1(n_590),
.B2(n_603),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_629),
.B(n_640),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_646),
.B(n_640),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_638),
.B(n_592),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_631),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_676),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_676),
.Y(n_679)
);

AOI221xp5_ASAP7_75t_L g680 ( 
.A1(n_660),
.A2(n_661),
.B1(n_657),
.B2(n_654),
.C(n_652),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_629),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_663),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_672),
.B(n_647),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_650),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_677),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_677),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_653),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_671),
.B(n_618),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_655),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_658),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_659),
.B(n_642),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_656),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_673),
.B(n_639),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_664),
.B(n_643),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_662),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_664),
.B(n_625),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_683),
.A2(n_675),
.B1(n_619),
.B2(n_618),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_680),
.B(n_665),
.C(n_669),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_684),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_681),
.B(n_650),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_686),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_696),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_686),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_683),
.A2(n_675),
.B(n_599),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_682),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_688),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_688),
.B(n_644),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_700),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_698),
.A2(n_695),
.B1(n_687),
.B2(n_689),
.C(n_690),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_681),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_704),
.A2(n_707),
.B(n_702),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_699),
.B(n_691),
.Y(n_712)
);

OAI21xp33_ASAP7_75t_L g713 ( 
.A1(n_697),
.A2(n_666),
.B(n_669),
.Y(n_713)
);

AOI21xp33_ASAP7_75t_SL g714 ( 
.A1(n_703),
.A2(n_693),
.B(n_682),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_711),
.B(n_692),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_709),
.A2(n_666),
.B1(n_700),
.B2(n_675),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_SL g717 ( 
.A1(n_708),
.A2(n_656),
.B1(n_597),
.B2(n_705),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_710),
.B(n_712),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_674),
.B1(n_619),
.B2(n_649),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_SL g720 ( 
.A(n_715),
.B(n_714),
.C(n_703),
.Y(n_720)
);

OAI211xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_685),
.B(n_679),
.C(n_678),
.Y(n_721)
);

AND4x1_ASAP7_75t_L g722 ( 
.A(n_718),
.B(n_590),
.C(n_616),
.D(n_598),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_716),
.B(n_701),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_719),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_720),
.B(n_585),
.C(n_603),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_694),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_723),
.B(n_599),
.C(n_613),
.Y(n_727)
);

XNOR2x1_ASAP7_75t_L g728 ( 
.A(n_726),
.B(n_722),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_727),
.Y(n_729)
);

NAND3x1_ASAP7_75t_L g730 ( 
.A(n_725),
.B(n_721),
.C(n_552),
.Y(n_730)
);

NOR2x1_ASAP7_75t_L g731 ( 
.A(n_727),
.B(n_569),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_730),
.A2(n_701),
.B(n_585),
.Y(n_732)
);

NAND2x1_ASAP7_75t_L g733 ( 
.A(n_731),
.B(n_569),
.Y(n_733)
);

OA22x2_ASAP7_75t_L g734 ( 
.A1(n_729),
.A2(n_597),
.B1(n_674),
.B2(n_663),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_576),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_728),
.B(n_651),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_R g738 ( 
.A(n_737),
.B(n_572),
.Y(n_738)
);

OAI211xp5_ASAP7_75t_L g739 ( 
.A1(n_736),
.A2(n_576),
.B(n_572),
.C(n_619),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_735),
.B(n_651),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_734),
.A2(n_674),
.B1(n_576),
.B2(n_667),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_SL g742 ( 
.A1(n_733),
.A2(n_596),
.B1(n_634),
.B2(n_648),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_732),
.A2(n_639),
.B1(n_648),
.B2(n_668),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_743),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_740),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_SL g746 ( 
.A1(n_742),
.A2(n_738),
.B1(n_741),
.B2(n_739),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

AOI21xp33_ASAP7_75t_L g748 ( 
.A1(n_744),
.A2(n_668),
.B(n_670),
.Y(n_748)
);

OAI22x1_ASAP7_75t_L g749 ( 
.A1(n_745),
.A2(n_747),
.B1(n_746),
.B2(n_670),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_636),
.B(n_645),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_SL g751 ( 
.A(n_749),
.B(n_587),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_748),
.A2(n_591),
.B(n_578),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_750),
.B(n_578),
.Y(n_753)
);

OAI222xp33_ASAP7_75t_L g754 ( 
.A1(n_752),
.A2(n_591),
.B1(n_587),
.B2(n_636),
.C1(n_645),
.C2(n_588),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_753),
.A2(n_617),
.B(n_614),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_754),
.B1(n_638),
.B2(n_588),
.Y(n_756)
);


endmodule