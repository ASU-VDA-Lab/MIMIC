module fake_jpeg_29015_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_66),
.Y(n_115)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_23),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g154 ( 
.A(n_68),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_21),
.B(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_9),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_87),
.Y(n_129)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_8),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_96),
.Y(n_127)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_43),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_33),
.Y(n_135)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_44),
.B1(n_19),
.B2(n_26),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_123),
.A2(n_138),
.B1(n_146),
.B2(n_150),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_48),
.B1(n_30),
.B2(n_35),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_130),
.A2(n_36),
.B1(n_26),
.B2(n_32),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_20),
.B(n_42),
.C(n_47),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_131),
.B(n_157),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_147),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_60),
.B1(n_71),
.B2(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_56),
.B(n_19),
.C(n_33),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_28),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_75),
.A2(n_19),
.B1(n_42),
.B2(n_47),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_54),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_20),
.B1(n_47),
.B2(n_42),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_62),
.B(n_48),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_27),
.B1(n_20),
.B2(n_34),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_162),
.A2(n_18),
.B1(n_28),
.B2(n_32),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_166),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx6_ASAP7_75t_SL g249 ( 
.A(n_167),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_169),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_70),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_171),
.A2(n_216),
.B1(n_219),
.B2(n_18),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_176),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_45),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_118),
.B(n_35),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_180),
.B(n_207),
.Y(n_257)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_181),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_128),
.A2(n_98),
.B1(n_90),
.B2(n_82),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_214),
.B1(n_216),
.B2(n_125),
.Y(n_227)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_129),
.A2(n_26),
.B(n_34),
.C(n_32),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_45),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_208),
.Y(n_253)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_91),
.B1(n_88),
.B2(n_67),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_133),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_198),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_200),
.A2(n_211),
.B1(n_220),
.B2(n_40),
.Y(n_256)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_202),
.Y(n_264)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_140),
.B(n_159),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_111),
.B(n_70),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_206),
.B1(n_218),
.B2(n_120),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_36),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_50),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_212),
.B(n_215),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_128),
.A2(n_105),
.B1(n_34),
.B2(n_28),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_18),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_140),
.B(n_50),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_156),
.B(n_27),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_227),
.A2(n_234),
.B1(n_243),
.B2(n_248),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_229),
.A2(n_245),
.B(n_255),
.C(n_236),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_125),
.B1(n_142),
.B2(n_108),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_167),
.A2(n_123),
.B(n_138),
.C(n_27),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_142),
.B1(n_108),
.B2(n_121),
.Y(n_243)
);

AOI22x1_ASAP7_75t_L g244 ( 
.A1(n_168),
.A2(n_161),
.B1(n_121),
.B2(n_149),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_244),
.A2(n_43),
.B(n_2),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_247),
.A2(n_166),
.B1(n_50),
.B2(n_43),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_168),
.A2(n_161),
.B1(n_149),
.B2(n_112),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_192),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_252),
.B(n_204),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_258),
.B1(n_261),
.B2(n_204),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_179),
.A2(n_40),
.B1(n_69),
.B2(n_50),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_193),
.A2(n_69),
.B1(n_140),
.B2(n_50),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_217),
.CI(n_169),
.CON(n_268),
.SN(n_268)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_174),
.A2(n_173),
.B1(n_215),
.B2(n_196),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_211),
.B1(n_178),
.B2(n_186),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_265),
.A2(n_276),
.B1(n_295),
.B2(n_234),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_172),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_217),
.B(n_182),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_267),
.A2(n_271),
.B(n_288),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_268),
.A2(n_277),
.B(n_246),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_223),
.B(n_169),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_275),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_231),
.B(n_245),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_190),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_189),
.B1(n_170),
.B2(n_199),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_SL g277 ( 
.A(n_230),
.B(n_203),
.C(n_208),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_191),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_290),
.Y(n_329)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_249),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_205),
.B1(n_218),
.B2(n_206),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_282),
.A2(n_285),
.B1(n_292),
.B2(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_213),
.B1(n_183),
.B2(n_181),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_231),
.B(n_244),
.C(n_248),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_231),
.A2(n_185),
.B(n_188),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_228),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_222),
.B(n_219),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_194),
.C(n_187),
.Y(n_291)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

NOR4xp25_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_11),
.C(n_2),
.D(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_296),
.B(n_300),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_229),
.B(n_251),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_43),
.C(n_0),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_299),
.C(n_229),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_2),
.C(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_222),
.B(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_242),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_259),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_326),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_247),
.B1(n_243),
.B2(n_239),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g357 ( 
.A1(n_305),
.A2(n_313),
.B1(n_332),
.B2(n_336),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_283),
.A2(n_261),
.B1(n_221),
.B2(n_246),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_297),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_287),
.A2(n_237),
.B(n_229),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_321),
.B(n_324),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_264),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_328),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_250),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_318),
.C(n_268),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_251),
.C(n_242),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_229),
.B(n_236),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_297),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_267),
.A2(n_254),
.B(n_232),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_254),
.B1(n_224),
.B2(n_241),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_270),
.A2(n_240),
.A3(n_232),
.B1(n_241),
.B2(n_225),
.Y(n_327)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_278),
.B(n_240),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_265),
.A2(n_224),
.B1(n_259),
.B2(n_238),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_335),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_295),
.B(n_296),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_7),
.B(n_11),
.C(n_12),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_358),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_282),
.B1(n_269),
.B2(n_285),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_338),
.A2(n_332),
.B1(n_314),
.B2(n_328),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_277),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_363),
.C(n_367),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_300),
.Y(n_344)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_268),
.B(n_288),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_345),
.Y(n_377)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_311),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_361),
.Y(n_387)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_349),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_350),
.B(n_360),
.Y(n_393)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_313),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_352),
.Y(n_396)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_276),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_356),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_313),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_314),
.B1(n_324),
.B2(n_306),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_290),
.B(n_294),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_368),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_286),
.C(n_284),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_280),
.Y(n_364)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_309),
.A2(n_269),
.B1(n_273),
.B2(n_301),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_366),
.B1(n_303),
.B2(n_304),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_332),
.A2(n_273),
.B1(n_279),
.B2(n_293),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_7),
.C(n_11),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_319),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_369),
.A2(n_371),
.B1(n_346),
.B2(n_357),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_370),
.A2(n_373),
.B1(n_374),
.B2(n_383),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_366),
.A2(n_326),
.B1(n_330),
.B2(n_307),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_312),
.B1(n_316),
.B2(n_320),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_343),
.B1(n_342),
.B2(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_357),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_306),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_348),
.C(n_350),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_365),
.A2(n_316),
.B1(n_320),
.B2(n_315),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_315),
.B1(n_323),
.B2(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_392),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_357),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_347),
.A2(n_302),
.B1(n_322),
.B2(n_336),
.Y(n_389)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_354),
.A2(n_323),
.B1(n_322),
.B2(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_362),
.B(n_302),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_398),
.B(n_394),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_384),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_411),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_341),
.B1(n_360),
.B2(n_352),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_402),
.A2(n_425),
.B1(n_385),
.B2(n_392),
.Y(n_428)
);

FAx1_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_358),
.CI(n_341),
.CON(n_403),
.SN(n_403)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_419),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_364),
.Y(n_406)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_399),
.Y(n_407)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_410),
.A2(n_378),
.B1(n_361),
.B2(n_318),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_344),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_357),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_418),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_348),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_393),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_363),
.C(n_340),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_421),
.Y(n_445)
);

OAI21xp33_ASAP7_75t_L g419 ( 
.A1(n_377),
.A2(n_340),
.B(n_342),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_381),
.B(n_359),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_422),
.A2(n_423),
.B1(n_386),
.B2(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_381),
.B(n_368),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_390),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_428),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_388),
.B1(n_391),
.B2(n_387),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_431),
.A2(n_433),
.B1(n_410),
.B2(n_412),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_409),
.A2(n_370),
.B1(n_374),
.B2(n_373),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_432),
.A2(n_414),
.B1(n_420),
.B2(n_422),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_404),
.A2(n_388),
.B1(n_391),
.B2(n_380),
.Y(n_433)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_437),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_379),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_405),
.B(n_393),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_440),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_403),
.B(n_372),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_395),
.B(n_390),
.Y(n_441)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_367),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_402),
.C(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_454),
.B1(n_460),
.B2(n_431),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_448),
.B(n_462),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_426),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_458),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_433),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_428),
.A2(n_432),
.B1(n_414),
.B2(n_446),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_401),
.C(n_420),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_461),
.C(n_463),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_406),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_434),
.B1(n_401),
.B2(n_417),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_411),
.C(n_395),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_407),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_417),
.C(n_423),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_472),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_429),
.C(n_439),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_334),
.C(n_331),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_445),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_470),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_386),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_476),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_463),
.A2(n_430),
.B(n_434),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_479),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_408),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_474),
.B(n_475),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_448),
.A2(n_429),
.B(n_427),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_351),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_355),
.B(n_353),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_478),
.B(n_470),
.Y(n_490)
);

AO21x2_ASAP7_75t_SL g478 ( 
.A1(n_447),
.A2(n_454),
.B(n_458),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_456),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_408),
.B1(n_376),
.B2(n_336),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_471),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_484),
.Y(n_502)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_482),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_16),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_467),
.A2(n_325),
.B1(n_11),
.B2(n_13),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g486 ( 
.A(n_472),
.B(n_325),
.Y(n_486)
);

NOR2x1_ASAP7_75t_SL g497 ( 
.A(n_486),
.B(n_7),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_465),
.A2(n_325),
.B1(n_14),
.B2(n_16),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_473),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_469),
.C(n_468),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_466),
.C(n_478),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_498),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_491),
.A2(n_464),
.B(n_477),
.Y(n_494)
);

AO21x1_ASAP7_75t_L g504 ( 
.A1(n_494),
.A2(n_497),
.B(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_495),
.B(n_496),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_478),
.C(n_14),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_16),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_16),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_489),
.B(n_481),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_503),
.A2(n_507),
.B(n_499),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_504),
.A2(n_505),
.B(n_482),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_485),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_509),
.A2(n_510),
.B(n_511),
.Y(n_512)
);

A2O1A1O1Ixp25_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_490),
.B(n_501),
.C(n_486),
.D(n_496),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_510),
.A2(n_508),
.B(n_501),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_506),
.Y(n_514)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_512),
.B(n_483),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_17),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_17),
.Y(n_517)
);


endmodule