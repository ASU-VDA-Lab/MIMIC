module fake_jpeg_4665_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_23),
.B1(n_30),
.B2(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_50),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_38),
.B1(n_28),
.B2(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_30),
.B1(n_23),
.B2(n_17),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_15),
.B1(n_31),
.B2(n_21),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_26),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_70),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_80),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_84),
.B(n_82),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_101),
.Y(n_123)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_53),
.B1(n_66),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_49),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_43),
.B1(n_48),
.B2(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_108),
.B1(n_54),
.B2(n_39),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_62),
.B1(n_66),
.B2(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_84),
.B1(n_72),
.B2(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_64),
.B1(n_87),
.B2(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_124),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_125),
.B(n_74),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_63),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_101),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_63),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_44),
.C(n_73),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_110),
.C(n_104),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_116),
.B(n_126),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_147),
.B(n_16),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_152),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_140),
.C(n_153),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_146),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_90),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_96),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_159),
.Y(n_164)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_64),
.B1(n_65),
.B2(n_81),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_150),
.B1(n_121),
.B2(n_70),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_156),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_26),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_37),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_132),
.C(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_125),
.A3(n_115),
.B1(n_113),
.B2(n_128),
.C1(n_74),
.C2(n_134),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_173),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_99),
.B1(n_100),
.B2(n_97),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_179),
.B1(n_155),
.B2(n_153),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_135),
.C(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_99),
.B1(n_100),
.B2(n_118),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_21),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_181),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_95),
.B(n_114),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_31),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_159),
.C(n_138),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_196),
.C(n_203),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_135),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_143),
.Y(n_216)
);

NAND2x1_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_138),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_21),
.B(n_31),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_156),
.B1(n_136),
.B2(n_154),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_170),
.B1(n_169),
.B2(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_146),
.B1(n_143),
.B2(n_114),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_102),
.B1(n_37),
.B2(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_146),
.C(n_143),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_164),
.B(n_173),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_219),
.B(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_190),
.C(n_204),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_181),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_216),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_195),
.B(n_161),
.CI(n_169),
.CON(n_215),
.SN(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_177),
.B1(n_114),
.B2(n_102),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_187),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_193),
.B1(n_189),
.B2(n_195),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_222),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_221),
.C(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_230),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_203),
.C(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_199),
.C(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_102),
.B1(n_141),
.B2(n_10),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_31),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_31),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_21),
.Y(n_236)
);

OAI322xp33_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_212),
.A3(n_219),
.B1(n_215),
.B2(n_208),
.C1(n_207),
.C2(n_220),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_248),
.B(n_7),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_208),
.B(n_215),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_7),
.B(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_207),
.C(n_21),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_246),
.C(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_8),
.C(n_14),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_8),
.C(n_14),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_7),
.C(n_12),
.Y(n_247)
);

OAI322xp33_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_26),
.A3(n_6),
.B1(n_11),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_250),
.A2(n_3),
.B(n_9),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_252),
.B(n_257),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_258),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_37),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_240),
.C(n_9),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_4),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_249),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_244),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_263),
.B(n_267),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_266),
.C(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_0),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_254),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_1),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_261),
.A2(n_259),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_3),
.C(n_10),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_1),
.B(n_2),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_1),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_2),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_277),
.B(n_2),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_275),
.B(n_274),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_2),
.Y(n_280)
);


endmodule