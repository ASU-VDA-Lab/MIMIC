module real_aes_8570_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_1078;
wire n_495;
wire n_892;
wire n_994;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_973;
wire n_504;
wire n_725;
wire n_671;
wire n_1081;
wire n_960;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_756;
wire n_404;
wire n_728;
wire n_598;
wire n_713;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_1136;
wire n_579;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1033;
wire n_1028;
wire n_1014;
wire n_1083;
wire n_727;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_1090;
wire n_456;
wire n_717;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_719;
wire n_566;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_1102;
wire n_1076;
wire n_463;
wire n_601;
wire n_804;
wire n_396;
wire n_661;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g662 ( .A(n_0), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g730 ( .A(n_1), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_2), .A2(n_240), .B1(n_479), .B2(n_485), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g885 ( .A1(n_3), .A2(n_182), .B1(n_334), .B2(n_428), .C1(n_535), .C2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_4), .A2(n_255), .B1(n_488), .B2(n_626), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_5), .A2(n_119), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_6), .A2(n_166), .B1(n_605), .B2(n_657), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_7), .A2(n_109), .B1(n_741), .B2(n_969), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_8), .A2(n_95), .B1(n_535), .B2(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_9), .A2(n_236), .B1(n_468), .B2(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g899 ( .A(n_10), .B(n_900), .Y(n_899) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_11), .A2(n_226), .B1(n_411), .B2(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g1074 ( .A(n_11), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_12), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_13), .A2(n_176), .B1(n_491), .B2(n_824), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_14), .A2(n_360), .B1(n_435), .B2(n_643), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_15), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_16), .A2(n_164), .B1(n_505), .B2(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g679 ( .A(n_17), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_18), .A2(n_196), .B1(n_521), .B2(n_573), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_19), .A2(n_250), .B1(n_505), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_20), .A2(n_321), .B1(n_511), .B2(n_512), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_21), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g836 ( .A1(n_22), .A2(n_76), .B1(n_285), .B2(n_435), .C1(n_593), .C2(n_669), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_23), .A2(n_232), .B1(n_813), .B2(n_964), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_24), .A2(n_308), .B1(n_545), .B2(n_787), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_25), .Y(n_930) );
AOI22xp5_ASAP7_75t_SL g628 ( .A1(n_26), .A2(n_247), .B1(n_602), .B2(n_629), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_27), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_28), .A2(n_306), .B1(n_503), .B2(n_554), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_29), .A2(n_252), .B1(n_488), .B2(n_491), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_30), .A2(n_364), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_31), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_32), .A2(n_246), .B1(n_741), .B2(n_824), .Y(n_1023) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_33), .A2(n_133), .B1(n_411), .B2(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g1082 ( .A(n_34), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_35), .A2(n_179), .B1(n_474), .B2(n_486), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_36), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_37), .A2(n_64), .B1(n_741), .B2(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_38), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_39), .A2(n_67), .B1(n_491), .B2(n_790), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_40), .A2(n_73), .B1(n_657), .B2(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g707 ( .A(n_41), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_42), .A2(n_295), .B1(n_535), .B2(n_667), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_43), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_44), .A2(n_69), .B1(n_493), .B2(n_607), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_45), .A2(n_170), .B1(n_611), .B2(n_824), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_46), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_47), .A2(n_139), .B1(n_508), .B2(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_48), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g986 ( .A(n_49), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_50), .A2(n_366), .B1(n_577), .B2(n_665), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_51), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_52), .A2(n_214), .B1(n_442), .B2(n_530), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g1126 ( .A(n_53), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_54), .A2(n_324), .B1(n_533), .B2(n_570), .Y(n_917) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_55), .A2(n_301), .B1(n_320), .B2(n_532), .C1(n_533), .C2(n_534), .Y(n_531) );
AOI22xp5_ASAP7_75t_SL g625 ( .A1(n_56), .A2(n_315), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_57), .A2(n_300), .B1(n_883), .B2(n_982), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_58), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_59), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_60), .A2(n_134), .B1(n_779), .B2(n_847), .Y(n_846) );
AOI22xp5_ASAP7_75t_SL g736 ( .A1(n_61), .A2(n_223), .B1(n_505), .B2(n_627), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_62), .A2(n_88), .B1(n_441), .B2(n_568), .Y(n_801) );
INVx1_ASAP7_75t_L g686 ( .A(n_63), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_65), .A2(n_331), .B1(n_830), .B2(n_831), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_66), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_68), .A2(n_219), .B1(n_632), .B2(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_70), .B(n_534), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_71), .A2(n_205), .B1(n_511), .B2(n_1117), .Y(n_1116) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_72), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_74), .A2(n_362), .B1(n_547), .B2(n_558), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_75), .A2(n_272), .B1(n_441), .B2(n_577), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_77), .A2(n_107), .B1(n_535), .B2(n_831), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_78), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_79), .Y(n_928) );
INVx1_ASAP7_75t_L g1086 ( .A(n_80), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_81), .A2(n_142), .B1(n_609), .B2(n_834), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_82), .A2(n_354), .B1(n_491), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g728 ( .A(n_83), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_84), .A2(n_159), .B1(n_785), .B2(n_787), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_85), .A2(n_283), .B1(n_491), .B2(n_512), .Y(n_1115) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_86), .B(n_633), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_87), .A2(n_208), .B1(n_468), .B2(n_473), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_89), .A2(n_108), .B1(n_458), .B2(n_463), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_90), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_91), .A2(n_221), .B1(n_521), .B2(n_525), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_92), .A2(n_230), .B1(n_847), .B2(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g433 ( .A(n_93), .Y(n_433) );
INVx1_ASAP7_75t_L g683 ( .A(n_94), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_96), .A2(n_113), .B1(n_488), .B2(n_782), .Y(n_781) );
AOI22xp5_ASAP7_75t_SL g739 ( .A1(n_97), .A2(n_114), .B1(n_740), .B2(n_741), .Y(n_739) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_98), .A2(n_262), .B1(n_411), .B2(n_412), .Y(n_418) );
INVx1_ASAP7_75t_L g1071 ( .A(n_98), .Y(n_1071) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_99), .A2(n_100), .B1(n_458), .B2(n_463), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_101), .A2(n_271), .B1(n_474), .B2(n_604), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_102), .A2(n_357), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_103), .A2(n_355), .B1(n_611), .B2(n_612), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_104), .A2(n_372), .B1(n_658), .B2(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_105), .A2(n_377), .B1(n_969), .B2(n_1003), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_106), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_110), .A2(n_291), .B1(n_813), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_111), .A2(n_310), .B1(n_607), .B2(n_609), .Y(n_606) );
OA22x2_ASAP7_75t_L g497 ( .A1(n_112), .A2(n_498), .B1(n_499), .B2(n_536), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_112), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_115), .A2(n_209), .B1(n_485), .B2(n_633), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_116), .A2(n_129), .B1(n_741), .B2(n_834), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_117), .A2(n_121), .B1(n_533), .B2(n_643), .Y(n_1019) );
INVx1_ASAP7_75t_L g733 ( .A(n_118), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_120), .A2(n_350), .B1(n_527), .B2(n_577), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_122), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_123), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_124), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_125), .B(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_126), .A2(n_154), .B1(n_511), .B2(n_1099), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_127), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_128), .A2(n_244), .B1(n_604), .B2(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_130), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_131), .A2(n_282), .B1(n_463), .B2(n_485), .Y(n_653) );
INVx1_ASAP7_75t_L g1110 ( .A(n_132), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_132), .A2(n_1110), .B1(n_1112), .B2(n_1136), .Y(n_1111) );
INVx1_ASAP7_75t_L g1075 ( .A(n_133), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_135), .B(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_136), .A2(n_157), .B1(n_507), .B2(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_137), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_138), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_140), .A2(n_145), .B1(n_485), .B2(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_141), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_141), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_143), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_144), .A2(n_263), .B1(n_665), .B2(n_808), .Y(n_860) );
XNOR2x2_ASAP7_75t_L g647 ( .A(n_146), .B(n_648), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_147), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_148), .A2(n_197), .B1(n_629), .B2(n_696), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_149), .Y(n_845) );
INVx1_ASAP7_75t_L g996 ( .A(n_150), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_151), .A2(n_193), .B1(n_468), .B2(n_473), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_152), .A2(n_338), .B1(n_515), .B2(n_517), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_153), .A2(n_178), .B1(n_481), .B2(n_834), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_155), .A2(n_261), .B1(n_441), .B2(n_577), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g1094 ( .A1(n_156), .A2(n_242), .B1(n_545), .B2(n_779), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_158), .A2(n_361), .B1(n_435), .B2(n_643), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_160), .A2(n_266), .B1(n_512), .B2(n_967), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_161), .A2(n_187), .B1(n_474), .B2(n_790), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_162), .A2(n_276), .B1(n_527), .B2(n_530), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_163), .Y(n_913) );
AND2x6_ASAP7_75t_L g385 ( .A(n_165), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_165), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_167), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_168), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_169), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_171), .A2(n_358), .B1(n_554), .B2(n_790), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_172), .A2(n_239), .B1(n_530), .B2(n_535), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_173), .A2(n_373), .B1(n_741), .B2(n_824), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_174), .Y(n_908) );
AOI222xp33_ASAP7_75t_L g1011 ( .A1(n_175), .A2(n_189), .B1(n_211), .B2(n_441), .C1(n_669), .C2(n_886), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_177), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_180), .Y(n_931) );
INVx1_ASAP7_75t_L g448 ( .A(n_181), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_183), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_184), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_185), .A2(n_268), .B1(n_511), .B2(n_815), .Y(n_814) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_186), .A2(n_248), .B1(n_411), .B2(n_415), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_186), .B(n_1073), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_188), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_190), .A2(n_267), .B1(n_602), .B2(n_626), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_191), .A2(n_251), .B1(n_481), .B2(n_607), .Y(n_875) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_192), .A2(n_224), .B1(n_293), .B2(n_435), .C1(n_441), .C2(n_669), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_194), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g1128 ( .A(n_195), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_198), .A2(n_381), .B1(n_435), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g404 ( .A(n_199), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_200), .A2(n_337), .B1(n_458), .B2(n_481), .Y(n_692) );
INVx1_ASAP7_75t_L g445 ( .A(n_201), .Y(n_445) );
AOI22xp5_ASAP7_75t_SL g631 ( .A1(n_202), .A2(n_278), .B1(n_632), .B2(n_633), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_203), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_204), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_206), .A2(n_238), .B1(n_612), .B2(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_207), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_210), .A2(n_344), .B1(n_474), .B2(n_515), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_212), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_213), .B(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_215), .Y(n_858) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_216), .A2(n_249), .B1(n_527), .B2(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_217), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g1057 ( .A1(n_218), .A2(n_374), .B1(n_502), .B2(n_627), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_220), .Y(n_589) );
INVx1_ASAP7_75t_L g1085 ( .A(n_222), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_225), .A2(n_347), .B1(n_813), .B2(n_964), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_227), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_228), .A2(n_944), .B1(n_972), .B2(n_973), .Y(n_943) );
INVx1_ASAP7_75t_L g972 ( .A(n_228), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_229), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_231), .A2(n_370), .B1(n_612), .B2(n_787), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_233), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_234), .A2(n_298), .B1(n_515), .B2(n_547), .Y(n_923) );
XNOR2xp5_ASAP7_75t_L g795 ( .A(n_235), .B(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_237), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_241), .A2(n_378), .B1(n_468), .B2(n_508), .Y(n_924) );
INVx2_ASAP7_75t_L g390 ( .A(n_243), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_245), .A2(n_329), .B1(n_435), .B2(n_442), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_253), .A2(n_265), .B1(n_626), .B2(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1081 ( .A(n_254), .Y(n_1081) );
OA22x2_ASAP7_75t_L g673 ( .A1(n_256), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_256), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_257), .A2(n_290), .B1(n_609), .B2(n_658), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_258), .A2(n_839), .B1(n_868), .B2(n_869), .Y(n_838) );
INVx1_ASAP7_75t_L g868 ( .A(n_258), .Y(n_868) );
INVx1_ASAP7_75t_L g1091 ( .A(n_259), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_260), .A2(n_313), .B1(n_635), .B2(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g704 ( .A(n_264), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_269), .A2(n_380), .B1(n_507), .B2(n_508), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_270), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_273), .A2(n_311), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_274), .A2(n_319), .B1(n_520), .B2(n_524), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_275), .A2(n_294), .B1(n_547), .B2(n_609), .Y(n_1004) );
NAND2xp5_ASAP7_75t_SL g898 ( .A(n_277), .B(n_573), .Y(n_898) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_279), .A2(n_383), .B(n_391), .C(n_1076), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_280), .A2(n_318), .B1(n_544), .B2(n_545), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_281), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_284), .A2(n_367), .B1(n_573), .B2(n_663), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_286), .Y(n_747) );
INVx1_ASAP7_75t_L g411 ( .A(n_287), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_287), .Y(n_413) );
INVx1_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
INVx1_ASAP7_75t_L g1044 ( .A(n_289), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_292), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_296), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_297), .Y(n_723) );
INVx1_ASAP7_75t_L g1042 ( .A(n_299), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_302), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_303), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_304), .A2(n_353), .B1(n_528), .B2(n_831), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_305), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_307), .B(n_1088), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_309), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_312), .A2(n_341), .B1(n_577), .B2(n_643), .Y(n_884) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_314), .B(n_521), .Y(n_806) );
AO22x2_ASAP7_75t_L g579 ( .A1(n_316), .A2(n_580), .B1(n_613), .B2(n_614), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_316), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_317), .A2(n_345), .B1(n_568), .B2(n_570), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_322), .Y(n_1134) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_323), .A2(n_1078), .B1(n_1101), .B2(n_1102), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_323), .Y(n_1101) );
AND2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_326), .A2(n_335), .B1(n_458), .B2(n_489), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_327), .Y(n_551) );
INVx1_ASAP7_75t_L g386 ( .A(n_328), .Y(n_386) );
XOR2x2_ASAP7_75t_L g999 ( .A(n_330), .B(n_1000), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_332), .B(n_883), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_333), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g731 ( .A(n_336), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_339), .Y(n_951) );
AOI22xp5_ASAP7_75t_SL g909 ( .A1(n_340), .A2(n_910), .B1(n_932), .B2(n_933), .Y(n_909) );
INVx1_ASAP7_75t_L g933 ( .A(n_340), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_342), .A2(n_359), .B1(n_665), .B2(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g689 ( .A(n_343), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_346), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_348), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_349), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_351), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_352), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_356), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_363), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_365), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_368), .A2(n_539), .B1(n_540), .B2(n_578), .Y(n_538) );
INVx1_ASAP7_75t_L g578 ( .A(n_368), .Y(n_578) );
INVx1_ASAP7_75t_L g681 ( .A(n_369), .Y(n_681) );
INVx1_ASAP7_75t_L g1090 ( .A(n_371), .Y(n_1090) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_375), .Y(n_1046) );
OA22x2_ASAP7_75t_L g757 ( .A1(n_376), .A2(n_758), .B1(n_759), .B2(n_791), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_376), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_379), .Y(n_1016) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_386), .Y(n_1067) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_387), .A2(n_1066), .B(n_1109), .Y(n_1108) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_793), .B1(n_1061), .B2(n_1062), .C(n_1063), .Y(n_391) );
INVxp67_ASAP7_75t_L g1061 ( .A(n_392), .Y(n_1061) );
AOI22xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B1(n_757), .B2(n_792), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI22xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_617), .B1(n_618), .B2(n_756), .Y(n_394) );
INVx1_ASAP7_75t_L g756 ( .A(n_395), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_494), .B1(n_495), .B2(n_616), .Y(n_395) );
INVx1_ASAP7_75t_L g616 ( .A(n_396), .Y(n_616) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_455), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_426), .C(n_444), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_421), .B2(n_422), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_405), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
OAI221xp5_ASAP7_75t_SL g857 ( .A1(n_405), .A2(n_422), .B1(n_858), .B2(n_859), .C(n_860), .Y(n_857) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g584 ( .A(n_406), .Y(n_584) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_406), .Y(n_1043) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_407), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_407), .A2(n_704), .B(n_705), .Y(n_703) );
OAI22xp5_ASAP7_75t_SL g912 ( .A1(n_407), .A2(n_423), .B1(n_913), .B2(n_914), .Y(n_912) );
BUFx3_ASAP7_75t_L g1125 ( .A(n_407), .Y(n_1125) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_416), .Y(n_407) );
INVx2_ASAP7_75t_L g484 ( .A(n_408), .Y(n_484) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_414), .Y(n_408) );
AND2x2_ASAP7_75t_L g425 ( .A(n_409), .B(n_414), .Y(n_425) );
AND2x2_ASAP7_75t_L g462 ( .A(n_409), .B(n_439), .Y(n_462) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g430 ( .A(n_410), .B(n_414), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_410), .B(n_420), .Y(n_440) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_413), .Y(n_415) );
INVx2_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_417), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g486 ( .A(n_417), .B(n_462), .Y(n_486) );
AND2x4_ASAP7_75t_L g523 ( .A(n_417), .B(n_484), .Y(n_523) );
AND2x6_ASAP7_75t_L g525 ( .A(n_417), .B(n_425), .Y(n_525) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g432 ( .A(n_418), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
INVx1_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_418), .B(n_420), .Y(n_466) );
AND2x2_ASAP7_75t_L g431 ( .A(n_419), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g461 ( .A(n_420), .B(n_454), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_422), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_678) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_423), .A2(n_446), .B1(n_707), .B2(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g765 ( .A(n_423), .Y(n_765) );
OA211x2_ASAP7_75t_L g880 ( .A1(n_423), .A2(n_881), .B(n_882), .C(n_884), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_423), .A2(n_584), .B1(n_947), .B2(n_948), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_423), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g587 ( .A(n_424), .Y(n_587) );
AND2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_461), .Y(n_472) );
AND2x4_ASAP7_75t_L g493 ( .A(n_425), .B(n_431), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_425), .B(n_461), .Y(n_726) );
OAI21xp33_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_433), .B(n_434), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_427), .A2(n_683), .B(n_684), .Y(n_682) );
OAI222xp33_ASAP7_75t_L g949 ( .A1(n_427), .A2(n_569), .B1(n_865), .B2(n_950), .C1(n_951), .C2(n_952), .Y(n_949) );
OAI21xp33_ASAP7_75t_L g1045 ( .A1(n_427), .A2(n_1046), .B(n_1047), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_427), .A2(n_769), .B1(n_1085), .B2(n_1086), .C(n_1087), .Y(n_1084) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g799 ( .A(n_428), .Y(n_799) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g532 ( .A(n_429), .Y(n_532) );
INVx4_ASAP7_75t_L g565 ( .A(n_429), .Y(n_565) );
INVx2_ASAP7_75t_L g639 ( .A(n_429), .Y(n_639) );
INVx2_ASAP7_75t_SL g711 ( .A(n_429), .Y(n_711) );
INVx2_ASAP7_75t_L g894 ( .A(n_429), .Y(n_894) );
AND2x6_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g451 ( .A(n_430), .Y(n_451) );
AND2x4_ASAP7_75t_L g530 ( .A(n_430), .B(n_453), .Y(n_530) );
AND2x6_ASAP7_75t_L g483 ( .A(n_431), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g490 ( .A(n_431), .B(n_462), .Y(n_490) );
INVx4_ASAP7_75t_L g569 ( .A(n_435), .Y(n_569) );
INVx2_ASAP7_75t_L g753 ( .A(n_435), .Y(n_753) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx4f_ASAP7_75t_SL g533 ( .A(n_436), .Y(n_533) );
BUFx2_ASAP7_75t_L g592 ( .A(n_436), .Y(n_592) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_436), .Y(n_688) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_436), .Y(n_886) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_438), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_439), .Y(n_447) );
AND2x4_ASAP7_75t_L g442 ( .A(n_440), .B(n_443), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_440), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g528 ( .A(n_440), .B(n_529), .Y(n_528) );
BUFx4f_ASAP7_75t_L g570 ( .A(n_441), .Y(n_570) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx12f_ASAP7_75t_L g535 ( .A(n_442), .Y(n_535) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_442), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_448), .B2(n_449), .Y(n_444) );
INVx4_ASAP7_75t_L g598 ( .A(n_446), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_446), .A2(n_686), .B1(n_687), .B2(n_689), .Y(n_685) );
BUFx3_ASAP7_75t_L g774 ( .A(n_446), .Y(n_774) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_446), .Y(n_955) );
AND2x2_ASAP7_75t_L g633 ( .A(n_447), .B(n_465), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_449), .A2(n_773), .B1(n_774), .B2(n_775), .Y(n_772) );
OAI22xp5_ASAP7_75t_SL g918 ( .A1(n_449), .A2(n_746), .B1(n_919), .B2(n_920), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_449), .A2(n_746), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_450), .A2(n_596), .B1(n_597), .B2(n_599), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g958 ( .A(n_450), .Y(n_958) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_477), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
BUFx4f_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g780 ( .A(n_459), .Y(n_780) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx3_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
BUFx3_ASAP7_75t_L g824 ( .A(n_460), .Y(n_824) );
BUFx3_ASAP7_75t_L g971 ( .A(n_460), .Y(n_971) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_461), .B(n_462), .Y(n_562) );
AND2x4_ASAP7_75t_L g464 ( .A(n_462), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g852 ( .A(n_463), .Y(n_852) );
BUFx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g517 ( .A(n_464), .Y(n_517) );
BUFx3_ASAP7_75t_L g547 ( .A(n_464), .Y(n_547) );
BUFx3_ASAP7_75t_L g612 ( .A(n_464), .Y(n_612) );
BUFx3_ASAP7_75t_L g632 ( .A(n_464), .Y(n_632) );
INVx1_ASAP7_75t_L g724 ( .A(n_464), .Y(n_724) );
BUFx3_ASAP7_75t_L g741 ( .A(n_464), .Y(n_741) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x6_ASAP7_75t_L g475 ( .A(n_466), .B(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g507 ( .A(n_470), .Y(n_507) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_470), .Y(n_549) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g604 ( .A(n_471), .Y(n_604) );
INVx3_ASAP7_75t_L g627 ( .A(n_471), .Y(n_627) );
INVx1_ASAP7_75t_L g657 ( .A(n_471), .Y(n_657) );
INVx5_ASAP7_75t_L g790 ( .A(n_471), .Y(n_790) );
INVx8_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g508 ( .A(n_474), .Y(n_508) );
BUFx2_ASAP7_75t_L g605 ( .A(n_474), .Y(n_605) );
BUFx4f_ASAP7_75t_SL g813 ( .A(n_474), .Y(n_813) );
INVx6_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g658 ( .A(n_475), .Y(n_658) );
INVx1_ASAP7_75t_SL g855 ( .A(n_475), .Y(n_855) );
INVx1_ASAP7_75t_SL g995 ( .A(n_475), .Y(n_995) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_480), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx5_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g611 ( .A(n_482), .Y(n_611) );
INVx1_ASAP7_75t_L g651 ( .A(n_482), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_482), .B(n_730), .Y(n_729) );
INVx4_ASAP7_75t_L g815 ( .A(n_482), .Y(n_815) );
INVx2_ASAP7_75t_L g1096 ( .A(n_482), .Y(n_1096) );
INVx11_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx11_ASAP7_75t_L g513 ( .A(n_483), .Y(n_513) );
INVx4_ASAP7_75t_L g516 ( .A(n_485), .Y(n_516) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g609 ( .A(n_486), .Y(n_609) );
BUFx3_ASAP7_75t_L g635 ( .A(n_486), .Y(n_635) );
INVx2_ASAP7_75t_L g715 ( .A(n_486), .Y(n_715) );
BUFx3_ASAP7_75t_L g787 ( .A(n_486), .Y(n_787) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g511 ( .A(n_489), .Y(n_511) );
BUFx3_ASAP7_75t_L g847 ( .A(n_489), .Y(n_847) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_490), .Y(n_558) );
INVx2_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
BUFx2_ASAP7_75t_SL g629 ( .A(n_490), .Y(n_629) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g502 ( .A(n_492), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_492), .A2(n_608), .B1(n_719), .B2(n_720), .Y(n_718) );
INVx2_ASAP7_75t_L g826 ( .A(n_492), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_492), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
INVx2_ASAP7_75t_L g967 ( .A(n_492), .Y(n_967) );
INVx6_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx3_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
BUFx3_ASAP7_75t_L g602 ( .A(n_493), .Y(n_602) );
BUFx3_ASAP7_75t_L g652 ( .A(n_493), .Y(n_652) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AO22x1_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_537), .B2(n_615), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g536 ( .A(n_499), .Y(n_536) );
NAND4xp75_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .C(n_518), .D(n_531), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g626 ( .A(n_513), .Y(n_626) );
INVx4_ASAP7_75t_L g740 ( .A(n_513), .Y(n_740) );
INVx4_ASAP7_75t_L g1003 ( .A(n_513), .Y(n_1003) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g544 ( .A(n_516), .Y(n_544) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_519), .B(n_526), .Y(n_518) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
INVx5_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g663 ( .A(n_522), .Y(n_663) );
INVx2_ASAP7_75t_L g883 ( .A(n_522), .Y(n_883) );
INVx2_ASAP7_75t_L g900 ( .A(n_522), .Y(n_900) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_525), .Y(n_573) );
BUFx2_ASAP7_75t_L g982 ( .A(n_525), .Y(n_982) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g643 ( .A(n_528), .Y(n_643) );
INVx1_ASAP7_75t_L g666 ( .A(n_528), .Y(n_666) );
BUFx2_ASAP7_75t_L g830 ( .A(n_528), .Y(n_830) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_530), .Y(n_577) );
BUFx2_ASAP7_75t_SL g667 ( .A(n_530), .Y(n_667) );
BUFx3_ASAP7_75t_L g831 ( .A(n_530), .Y(n_831) );
BUFx2_ASAP7_75t_SL g1048 ( .A(n_530), .Y(n_1048) );
INVx3_ASAP7_75t_L g590 ( .A(n_532), .Y(n_590) );
INVx1_ASAP7_75t_L g862 ( .A(n_533), .Y(n_862) );
BUFx4f_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g594 ( .A(n_535), .Y(n_594) );
INVx1_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_579), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_541), .B(n_563), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_550), .C(n_555), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g782 ( .A(n_553), .Y(n_782) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_559), .B2(n_560), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_557), .A2(n_560), .B1(n_930), .B2(n_931), .Y(n_929) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_562), .B(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B(n_567), .Y(n_564) );
INVx4_ASAP7_75t_L g669 ( .A(n_565), .Y(n_669) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_565), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
BUFx2_ASAP7_75t_L g767 ( .A(n_565), .Y(n_767) );
OAI21xp5_ASAP7_75t_SL g915 ( .A1(n_565), .A2(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g769 ( .A(n_568), .Y(n_769) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_569), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .C(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g805 ( .A(n_573), .Y(n_805) );
INVx1_ASAP7_75t_SL g809 ( .A(n_577), .Y(n_809) );
INVx1_ASAP7_75t_SL g613 ( .A(n_580), .Y(n_613) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_581), .B(n_600), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_588), .C(n_595), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_586), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g661 ( .A(n_587), .Y(n_661) );
INVx1_ASAP7_75t_SL g1083 ( .A(n_587), .Y(n_1083) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_591), .Y(n_588) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_SL g746 ( .A(n_598), .Y(n_746) );
AND4x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .C(n_606), .D(n_610), .Y(n_600) );
INVx1_ASAP7_75t_L g844 ( .A(n_602), .Y(n_844) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx3_ASAP7_75t_L g834 ( .A(n_608), .Y(n_834) );
BUFx2_ASAP7_75t_L g850 ( .A(n_609), .Y(n_850) );
INVx1_ASAP7_75t_L g786 ( .A(n_611), .Y(n_786) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
XOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_670), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_646), .B2(n_647), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
XOR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_645), .Y(n_623) );
NAND4xp75_ASAP7_75t_SL g624 ( .A(n_625), .B(n_628), .C(n_630), .D(n_636), .Y(n_624) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND4xp75_ASAP7_75t_L g648 ( .A(n_649), .B(n_654), .C(n_659), .D(n_668), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
INVx2_ASAP7_75t_L g842 ( .A(n_651), .Y(n_842) );
INVx3_ASAP7_75t_L g697 ( .A(n_652), .Y(n_697) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
OA211x2_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B(n_662), .C(n_664), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_661), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AO22x2_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_699), .B2(n_755), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_690), .Y(n_676) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_682), .C(n_685), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g748 ( .A1(n_680), .A2(n_749), .B(n_750), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_680), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1080) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g755 ( .A(n_699), .Y(n_755) );
XOR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_732), .Y(n_699) );
XNOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_731), .Y(n_700) );
AND3x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_713), .C(n_721), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .C(n_709), .Y(n_702) );
OAI222xp33_ASAP7_75t_L g861 ( .A1(n_711), .A2(n_862), .B1(n_863), .B2(n_864), .C1(n_865), .C2(n_867), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g962 ( .A(n_715), .Y(n_962) );
INVx2_ASAP7_75t_L g1120 ( .A(n_715), .Y(n_1120) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_727), .C(n_729), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_722) );
XNOR2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND3x1_ASAP7_75t_SL g734 ( .A(n_735), .B(n_738), .C(n_743), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .C(n_751), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_746), .A2(n_957), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
INVx1_ASAP7_75t_L g792 ( .A(n_757), .Y(n_792) );
INVx1_ASAP7_75t_L g791 ( .A(n_759), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_776), .Y(n_759) );
NOR3xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_766), .C(n_772), .Y(n_760) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_770), .C(n_771), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_767), .A2(n_1128), .B1(n_1129), .B2(n_1130), .C(n_1131), .Y(n_1127) );
NOR2xp67_ASAP7_75t_L g776 ( .A(n_777), .B(n_783), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_788), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_787), .Y(n_1099) );
BUFx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_790), .Y(n_964) );
INVx1_ASAP7_75t_L g1062 ( .A(n_793), .Y(n_1062) );
XOR2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_939), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_817), .B1(n_937), .B2(n_938), .Y(n_794) );
INVx1_ASAP7_75t_L g937 ( .A(n_795), .Y(n_937) );
NAND4xp75_ASAP7_75t_SL g796 ( .A(n_797), .B(n_810), .C(n_814), .D(n_816), .Y(n_796) );
NOR2xp67_ASAP7_75t_L g797 ( .A(n_798), .B(n_802), .Y(n_797) );
OAI21xp5_ASAP7_75t_SL g798 ( .A1(n_799), .A2(n_800), .B(n_801), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .C(n_807), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_SL g927 ( .A(n_815), .Y(n_927) );
INVx1_ASAP7_75t_L g938 ( .A(n_817), .Y(n_938) );
XOR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_871), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_838), .B2(n_870), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
XOR2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_837), .Y(n_820) );
NAND4xp75_ASAP7_75t_L g821 ( .A(n_822), .B(n_827), .C(n_832), .D(n_836), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
BUFx3_ASAP7_75t_L g1117 ( .A(n_824), .Y(n_1117) );
AND2x2_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .Y(n_827) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g870 ( .A(n_838), .Y(n_870) );
INVx1_ASAP7_75t_L g869 ( .A(n_839), .Y(n_869) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_856), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_848), .Y(n_840) );
OAI221xp5_ASAP7_75t_SL g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_845), .C(n_846), .Y(n_841) );
OAI221xp5_ASAP7_75t_SL g848 ( .A1(n_849), .A2(n_851), .B1(n_852), .B2(n_853), .C(n_854), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2xp33_ASAP7_75t_SL g856 ( .A(n_857), .B(n_861), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_862), .A2(n_955), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_866), .Y(n_1088) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_866), .Y(n_1132) );
AO22x1_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_888), .B1(n_889), .B2(n_936), .Y(n_871) );
INVx2_ASAP7_75t_SL g936 ( .A(n_872), .Y(n_936) );
XOR2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_887), .Y(n_872) );
NAND4xp75_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .C(n_880), .D(n_885), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1129 ( .A(n_886), .Y(n_1129) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AO22x2_ASAP7_75t_SL g889 ( .A1(n_890), .A2(n_909), .B1(n_934), .B2(n_935), .Y(n_889) );
INVx4_ASAP7_75t_SL g934 ( .A(n_890), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_890), .A2(n_934), .B1(n_943), .B2(n_974), .Y(n_942) );
XOR2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_908), .Y(n_890) );
NAND3x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_902), .C(n_905), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_897), .Y(n_892) );
OAI21xp5_ASAP7_75t_SL g893 ( .A1(n_894), .A2(n_895), .B(n_896), .Y(n_893) );
OAI21xp5_ASAP7_75t_SL g985 ( .A1(n_894), .A2(n_986), .B(n_987), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_894), .A2(n_1016), .B(n_1017), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .C(n_901), .Y(n_897) );
AND2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
AND2x2_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g935 ( .A(n_909), .Y(n_935) );
INVx1_ASAP7_75t_L g932 ( .A(n_910), .Y(n_932) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_921), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .C(n_918), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_929), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
AOI22xp5_ASAP7_75t_SL g939 ( .A1(n_940), .A2(n_1033), .B1(n_1034), .B2(n_1060), .Y(n_939) );
INVx1_ASAP7_75t_L g1060 ( .A(n_940), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B1(n_975), .B2(n_1032), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g974 ( .A(n_943), .Y(n_974) );
INVx1_ASAP7_75t_L g973 ( .A(n_944), .Y(n_973) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_959), .Y(n_944) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_949), .C(n_953), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_953) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_965), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_963), .Y(n_960) );
NAND2xp5_ASAP7_75t_SL g965 ( .A(n_966), .B(n_968), .Y(n_965) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1032 ( .A(n_975), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_997), .B1(n_998), .B2(n_1031), .Y(n_975) );
INVx1_ASAP7_75t_SL g1031 ( .A(n_976), .Y(n_1031) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
XOR2x2_ASAP7_75t_SL g977 ( .A(n_978), .B(n_996), .Y(n_977) );
NAND2x1p5_ASAP7_75t_L g978 ( .A(n_979), .B(n_988), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_985), .Y(n_979) );
NAND3xp33_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .C(n_984), .Y(n_980) );
NOR2x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
AO22x1_ASAP7_75t_SL g998 ( .A1(n_999), .A2(n_1012), .B1(n_1029), .B2(n_1030), .Y(n_998) );
INVx1_ASAP7_75t_L g1029 ( .A(n_999), .Y(n_1029) );
NAND4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1005), .C(n_1008), .D(n_1011), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1004), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1007), .Y(n_1005) );
AND2x2_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
INVx3_ASAP7_75t_SL g1030 ( .A(n_1012), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_1012), .A2(n_1030), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
XOR2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1028), .Y(n_1012) );
NAND2xp5_ASAP7_75t_SL g1013 ( .A(n_1014), .B(n_1021), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1018), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_SL g1037 ( .A(n_1038), .Y(n_1037) );
XNOR2x1_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1059), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1052), .Y(n_1039) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1045), .C(n_1049), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1056), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
INVx1_ASAP7_75t_SL g1063 ( .A(n_1064), .Y(n_1063) );
NOR2x1_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1069), .Y(n_1064) );
OR2x2_ASAP7_75t_SL g1139 ( .A(n_1065), .B(n_1070), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1068), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
OAI322xp33_ASAP7_75t_L g1076 ( .A1(n_1067), .A2(n_1077), .A3(n_1103), .B1(n_1107), .B2(n_1110), .C1(n_1111), .C2(n_1137), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1067), .B(n_1106), .Y(n_1109) );
CKINVDCx16_ASAP7_75t_R g1106 ( .A(n_1068), .Y(n_1106) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_1070), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1075), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_1078), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1092), .Y(n_1078) );
NOR3xp33_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1084), .C(n_1089), .Y(n_1079) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1097), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1100), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_SL g1136 ( .A(n_1112), .Y(n_1136) );
AND2x2_ASAP7_75t_SL g1112 ( .A(n_1113), .B(n_1122), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1118), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1121), .Y(n_1118) );
NOR3xp33_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1127), .C(n_1133), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g1137 ( .A(n_1138), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g1138 ( .A(n_1139), .Y(n_1138) );
endmodule