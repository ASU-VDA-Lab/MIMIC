module fake_ariane_3074_n_197 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_197);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_197;

wire n_83;
wire n_56;
wire n_60;
wire n_190;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVxp33_ASAP7_75t_SL g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_37),
.Y(n_62)
);

AO21x2_ASAP7_75t_L g63 ( 
.A1(n_33),
.A2(n_59),
.B(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_0),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_5),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_35),
.A2(n_6),
.B1(n_12),
.B2(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_R g85 ( 
.A(n_76),
.B(n_44),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_54),
.B(n_38),
.C(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_69),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_44),
.B(n_57),
.C(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

HB1xp67_ASAP7_75t_SL g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_76),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

AOI221x1_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_82),
.B1(n_73),
.B2(n_75),
.C(n_74),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_69),
.Y(n_109)
);

NAND3x1_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_81),
.C(n_75),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_63),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_63),
.Y(n_114)
);

AO31x2_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_74),
.A3(n_63),
.B(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_71),
.B(n_62),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_103),
.B(n_100),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx9p33_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_68),
.B(n_60),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_99),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_67),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_67),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_90),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_86),
.B(n_95),
.C(n_97),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_93),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_99),
.B1(n_92),
.B2(n_105),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_92),
.B(n_123),
.C(n_113),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_124),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_124),
.B1(n_110),
.B2(n_120),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_108),
.B(n_112),
.C(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_111),
.B1(n_120),
.B2(n_117),
.Y(n_135)
);

O2A1O1Ixp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_101),
.B(n_118),
.C(n_109),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_109),
.B(n_114),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_103),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_103),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_61),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_114),
.B(n_123),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_93),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_84),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_103),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_100),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_136),
.B(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_127),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_144),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_141),
.Y(n_158)
);

AOI211xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_128),
.B(n_141),
.C(n_135),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_126),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_154),
.B(n_152),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_155),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_160),
.B(n_163),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_156),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_150),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_151),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_158),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_155),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_171),
.B1(n_159),
.B2(n_160),
.C(n_165),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_180),
.B1(n_162),
.B2(n_176),
.C(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_166),
.B(n_162),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

AOI211x1_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_180),
.B(n_164),
.C(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_183),
.C(n_184),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_191),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_192),
.B(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_194),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_162),
.B(n_168),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_182),
.B1(n_185),
.B2(n_169),
.C(n_170),
.Y(n_197)
);


endmodule