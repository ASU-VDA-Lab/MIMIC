module fake_jpeg_3871_n_283 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_283);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_46),
.CON(n_74),
.SN(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_30),
.B1(n_19),
.B2(n_15),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_59),
.B(n_27),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_62),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_31),
.B1(n_16),
.B2(n_30),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_80),
.B1(n_84),
.B2(n_97),
.Y(n_123)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_13),
.C(n_22),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_8),
.B(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_24),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_23),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_26),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_91),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_36),
.A2(n_28),
.B1(n_14),
.B2(n_27),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_40),
.Y(n_91)
);

BUFx2_ASAP7_75t_R g94 ( 
.A(n_33),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_26),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_14),
.B1(n_27),
.B2(n_2),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_25),
.B1(n_18),
.B2(n_28),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_109),
.B1(n_96),
.B2(n_74),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_14),
.B1(n_7),
.B2(n_3),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_74),
.B(n_47),
.C(n_48),
.Y(n_129)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_136),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_90),
.B1(n_50),
.B2(n_59),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_81),
.B1(n_87),
.B2(n_64),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_141),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_94),
.B(n_65),
.C(n_47),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_156),
.B(n_122),
.Y(n_170)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_79),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_60),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_67),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_75),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_75),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_83),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_70),
.B(n_83),
.C(n_6),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_98),
.B1(n_120),
.B2(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_73),
.B1(n_63),
.B2(n_66),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_116),
.B1(n_114),
.B2(n_100),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_155),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_63),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_111),
.B(n_1),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_98),
.B(n_112),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_118),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_175),
.Y(n_209)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_107),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_141),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_167),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_184),
.B(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_101),
.B1(n_122),
.B2(n_116),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_180),
.B1(n_137),
.B2(n_142),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_70),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_100),
.A3(n_114),
.B1(n_113),
.B2(n_125),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_125),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_145),
.B(n_155),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_102),
.B(n_93),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_153),
.B(n_136),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_132),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_193),
.C(n_198),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_147),
.C(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_200),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_210),
.B1(n_173),
.B2(n_169),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_128),
.C(n_158),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_127),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_173),
.B(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_156),
.Y(n_206)
);

OAI322xp33_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_192),
.A3(n_191),
.B1(n_203),
.B2(n_205),
.C1(n_207),
.C2(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_183),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_130),
.B1(n_139),
.B2(n_129),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_167),
.B1(n_187),
.B2(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_156),
.B1(n_148),
.B2(n_140),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_212),
.B(n_186),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_127),
.B(n_1),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_66),
.Y(n_214)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_179),
.B(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_231),
.C(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_226),
.B(n_230),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_235),
.A2(n_248),
.B(n_249),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_213),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_247),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_202),
.C(n_201),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_231),
.C(n_242),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_227),
.B(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_259),
.B1(n_163),
.B2(n_241),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_216),
.B1(n_219),
.B2(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_162),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_260),
.B(n_240),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_235),
.Y(n_263)
);

OA21x2_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_242),
.B(n_237),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_223),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_241),
.B1(n_233),
.B2(n_161),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_249),
.C(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_267),
.B1(n_196),
.B2(n_268),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_174),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_176),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_276),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_240),
.C(n_214),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_278),
.B(n_188),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_279),
.Y(n_283)
);


endmodule