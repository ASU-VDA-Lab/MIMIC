module fake_jpeg_1439_n_312 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_66),
.Y(n_109)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_0),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_77),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_18),
.B1(n_66),
.B2(n_64),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_21),
.B1(n_32),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_34),
.B1(n_24),
.B2(n_38),
.Y(n_77)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_40),
.B1(n_29),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_83),
.B1(n_95),
.B2(n_99),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_40),
.B1(n_29),
.B2(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_25),
.B1(n_33),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_87),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_102),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_28),
.B1(n_26),
.B2(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_52),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_20),
.B1(n_19),
.B2(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_20),
.B1(n_19),
.B2(n_6),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_102),
.B(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_111),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_46),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_15),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_114),
.A2(n_147),
.B1(n_128),
.B2(n_141),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_122),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_131),
.Y(n_152)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_14),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_123),
.B(n_127),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_124),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_9),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_10),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_80),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_11),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_125),
.B(n_124),
.Y(n_165)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_97),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_103),
.B(n_105),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_160),
.B(n_165),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_82),
.B1(n_78),
.B2(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_139),
.B1(n_145),
.B2(n_117),
.Y(n_193)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_69),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_169),
.C(n_175),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_110),
.B(n_69),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_82),
.B1(n_94),
.B2(n_103),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_162),
.B1(n_156),
.B2(n_154),
.Y(n_196)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_105),
.B1(n_94),
.B2(n_76),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_76),
.C(n_112),
.Y(n_169)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_132),
.C(n_136),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_183),
.Y(n_189)
);

AO22x2_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_135),
.B1(n_129),
.B2(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_149),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_129),
.A2(n_120),
.B1(n_146),
.B2(n_133),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_160),
.B(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_203),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_140),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_212),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_200),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_201),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_205),
.B1(n_171),
.B2(n_196),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_117),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_195),
.C(n_171),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_139),
.C(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_197),
.B1(n_207),
.B2(n_213),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_150),
.B1(n_162),
.B2(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_151),
.B(n_164),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_170),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_169),
.B(n_172),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_208),
.B(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_163),
.B1(n_183),
.B2(n_172),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_157),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_159),
.B1(n_166),
.B2(n_161),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_161),
.B(n_166),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_171),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_171),
.B1(n_191),
.B2(n_205),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_237),
.B(n_216),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_200),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_209),
.C(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_234),
.B1(n_226),
.B2(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_198),
.A2(n_188),
.B1(n_187),
.B2(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_229),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_187),
.B1(n_189),
.B2(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_186),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_213),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_216),
.B(n_237),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_209),
.B(n_185),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_250),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_255),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_214),
.B1(n_224),
.B2(n_215),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_248),
.B1(n_229),
.B2(n_228),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

NOR4xp25_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_230),
.C(n_236),
.D(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_251),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_266),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_250),
.B1(n_246),
.B2(n_245),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_244),
.B1(n_240),
.B2(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_231),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_268),
.Y(n_279)
);

XNOR2x2_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_240),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_220),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_218),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_239),
.C(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_259),
.C(n_265),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_276),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_249),
.B1(n_245),
.B2(n_254),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_267),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_256),
.B(n_241),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_254),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_253),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_270),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_259),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_291),
.C(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_280),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_282),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_SL g293 ( 
.A1(n_287),
.A2(n_273),
.B(n_271),
.C(n_277),
.Y(n_293)
);

AOI31xp33_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_296),
.A3(n_276),
.B(n_221),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_291),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_274),
.B(n_284),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_282),
.C(n_241),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_219),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_293),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_276),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_302),
.A2(n_303),
.B1(n_295),
.B2(n_296),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_306),
.B(n_302),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_227),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_308),
.Y(n_312)
);


endmodule