module real_jpeg_22394_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_0),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_0),
.A2(n_52),
.B1(n_53),
.B2(n_104),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_104),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_0),
.A2(n_28),
.B1(n_32),
.B2(n_104),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_92),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_2),
.A2(n_28),
.B1(n_32),
.B2(n_92),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_98),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_98),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_109),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_109),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_28),
.B1(n_32),
.B2(n_102),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_102),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_182)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_7),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_269)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_71),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_71),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_11),
.B(n_22),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_49),
.B(n_52),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_86),
.B1(n_87),
.B2(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_63),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_11),
.A2(n_25),
.B(n_197),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_13),
.A2(n_31),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_13),
.A2(n_31),
.B1(n_52),
.B2(n_53),
.Y(n_234)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_59),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_14),
.A2(n_25),
.A3(n_48),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_30),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B(n_28),
.C(n_29),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_22),
.A2(n_27),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_22),
.A2(n_27),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_25),
.Y(n_121)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_24),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_24),
.A2(n_29),
.B1(n_106),
.B2(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_24),
.B(n_107),
.Y(n_193)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g106 ( 
.A(n_28),
.B(n_107),
.CON(n_106),
.SN(n_106)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_34),
.B(n_41),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_76),
.B(n_332),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_72),
.C(n_74),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_42),
.A2(n_43),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_55),
.C(n_64),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_44),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_44),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_44),
.A2(n_55),
.B1(n_302),
.B2(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B(n_54),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_51),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_51),
.B1(n_91),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_45),
.A2(n_51),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_45),
.A2(n_51),
.B1(n_161),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_45),
.A2(n_51),
.B1(n_182),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_45),
.A2(n_51),
.B1(n_97),
.B2(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_45),
.A2(n_51),
.B1(n_93),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_45),
.A2(n_51),
.B1(n_236),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_45),
.A2(n_51),
.B1(n_54),
.B2(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_47),
.B(n_59),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_48),
.A2(n_50),
.B(n_107),
.C(n_157),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_51),
.B(n_107),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_53),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_55),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_62),
.B(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_57),
.A2(n_63),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_57),
.A2(n_63),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_61),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_61),
.B1(n_103),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_58),
.A2(n_61),
.B1(n_134),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_58),
.A2(n_61),
.B1(n_117),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_58),
.A2(n_61),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_64),
.A2(n_65),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_69),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_66),
.A2(n_69),
.B1(n_115),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_66),
.A2(n_69),
.B1(n_243),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_74),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_325),
.B(n_331),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_294),
.A3(n_317),
.B1(n_323),
.B2(n_324),
.C(n_334),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_273),
.B(n_293),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_249),
.B(n_272),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_140),
.B(n_225),
.C(n_248),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_125),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_82),
.B(n_125),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_110),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_84),
.B(n_94),
.C(n_110),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_85),
.B(n_90),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_88),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_123),
.B1(n_124),
.B2(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_86),
.A2(n_150),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_86),
.A2(n_124),
.B1(n_153),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_86),
.A2(n_124),
.B1(n_139),
.B2(n_184),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_86),
.A2(n_89),
.B1(n_166),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_86),
.A2(n_166),
.B(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_87),
.B(n_107),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_105),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_112),
.B(n_118),
.C(n_119),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_132),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_224),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_219),
.B(n_223),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_205),
.B(n_218),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_186),
.B(n_204),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_174),
.B(n_185),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_162),
.B(n_173),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_168),
.B(n_172),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_194),
.B1(n_202),
.B2(n_203),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_215),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_227),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_247),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_238),
.C(n_247),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_241),
.C(n_246),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_246),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_271),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_264),
.B2(n_265),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_265),
.C(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_257),
.C(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_267),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_268),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_267),
.A2(n_285),
.B(n_288),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_275),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_291),
.B2(n_292),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_284),
.C(n_292),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B(n_283),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_296),
.C(n_307),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_296),
.B1(n_297),
.B2(n_322),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_283),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_309),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_309),
.Y(n_324)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_303),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_306),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_311),
.C(n_316),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_308),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_328),
.Y(n_330)
);


endmodule