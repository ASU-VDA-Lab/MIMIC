module fake_jpeg_29597_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_70),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_55),
.B1(n_51),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_53),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_52),
.B1(n_51),
.B2(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_67),
.B1(n_58),
.B2(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_65),
.B1(n_48),
.B2(n_49),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_85),
.B1(n_88),
.B2(n_84),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_47),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_61),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_50),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_9),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_60),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_60),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_56),
.B1(n_60),
.B2(n_2),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_124),
.B1(n_128),
.B2(n_12),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_3),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_133),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_4),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_25),
.A3(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_30),
.B(n_39),
.C(n_17),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_21),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.C(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_24),
.C(n_42),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_11),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_154),
.B1(n_156),
.B2(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_12),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_29),
.C(n_38),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_33),
.C(n_18),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_128),
.B1(n_131),
.B2(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

OAI322xp33_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_155),
.A3(n_139),
.B1(n_141),
.B2(n_147),
.C1(n_145),
.C2(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_163),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B1(n_168),
.B2(n_160),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_169),
.B(n_158),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_159),
.B(n_20),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);


endmodule