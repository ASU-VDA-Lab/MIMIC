module fake_jpeg_19365_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_27),
.B1(n_14),
.B2(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_34),
.B1(n_27),
.B2(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_19),
.B1(n_13),
.B2(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_12),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_17),
.C(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_27),
.B1(n_19),
.B2(n_12),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B(n_36),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_26),
.B(n_23),
.C(n_22),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_29),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_43),
.C(n_44),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_8),
.C(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_36),
.B1(n_22),
.B2(n_20),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_28),
.B(n_36),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_36),
.B(n_32),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_40),
.B(n_37),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_48),
.B1(n_40),
.B2(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_3),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_18),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_18),
.B1(n_11),
.B2(n_10),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_2),
.B(n_3),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_59),
.B(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_53),
.B(n_60),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_72),
.B(n_75),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_68),
.B(n_52),
.C(n_18),
.D(n_11),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_76),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_5),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_84),
.C(n_89),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_20),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_86),
.B1(n_83),
.B2(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_6),
.A3(n_7),
.B1(n_11),
.B2(n_18),
.C1(n_32),
.C2(n_93),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_11),
.Y(n_105)
);


endmodule