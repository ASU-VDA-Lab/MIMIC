module fake_jpeg_15218_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_82),
.Y(n_98)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_46),
.B1(n_50),
.B2(n_54),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_77),
.B1(n_60),
.B2(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_61),
.B1(n_46),
.B2(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_54),
.B1(n_58),
.B2(n_55),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_89),
.B1(n_91),
.B2(n_10),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_61),
.B(n_53),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_6),
.B(n_7),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_57),
.B1(n_52),
.B2(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_49),
.B1(n_48),
.B2(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_94),
.B1(n_103),
.B2(n_83),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_49),
.B1(n_1),
.B2(n_3),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_102),
.B1(n_8),
.B2(n_9),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_26),
.B1(n_42),
.B2(n_41),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_111),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_10),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_113),
.B(n_114),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_81),
.B1(n_12),
.B2(n_13),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_95),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_104),
.B(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_119),
.C(n_118),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_114),
.B1(n_103),
.B2(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_115),
.B1(n_101),
.B2(n_90),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_11),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_115),
.B(n_18),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_124),
.C(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_134),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_129),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_127),
.B(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_20),
.B(n_21),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_141)
);

AOI21x1_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_28),
.B(n_29),
.Y(n_142)
);

OAI21x1_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_32),
.B(n_33),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_34),
.B(n_36),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_38),
.B(n_40),
.Y(n_146)
);


endmodule