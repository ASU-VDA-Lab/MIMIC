module fake_aes_10931_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NOR2xp67_ASAP7_75t_L g4 ( .A(n_2), .B(n_1), .Y(n_4) );
AOI21xp5_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
INVx4_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AND2x4_ASAP7_75t_SL g8 ( .A(n_7), .B(n_3), .Y(n_8) );
OAI221xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_7), .B1(n_5), .B2(n_4), .C(n_2), .Y(n_9) );
OAI21xp5_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_4), .B(n_0), .Y(n_10) );
XNOR2x1_ASAP7_75t_L g11 ( .A(n_10), .B(n_0), .Y(n_11) );
OAI21xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_1), .B(n_10), .Y(n_12) );
endmodule