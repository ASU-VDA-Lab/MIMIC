module fake_netlist_6_229_n_181 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_40, n_181);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;
input n_40;

output n_181;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_130;
wire n_84;
wire n_78;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_18),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

NOR2xp67_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_56),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_52),
.B(n_64),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_42),
.C(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_48),
.B1(n_54),
.B2(n_47),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_53),
.B(n_46),
.Y(n_89)
);

AOI21x1_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_45),
.B(n_43),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_65),
.B(n_49),
.C(n_5),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_25),
.B(n_37),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_8),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_9),
.B(n_12),
.C(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_81),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OR2x6_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_75),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_82),
.B(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_99),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2x1_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_82),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_75),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_82),
.B(n_70),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_81),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND4xp25_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_107),
.C(n_72),
.D(n_74),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_101),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_106),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_127),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_111),
.C(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_106),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_93),
.C(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_118),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_118),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_128),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_129),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_143),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_123),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

NAND2x1_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_149),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_138),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_109),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_154),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_109),
.C(n_39),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_82),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_36),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_78),
.B1(n_157),
.B2(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_78),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_173),
.B1(n_158),
.B2(n_175),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_157),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_177),
.B1(n_159),
.B2(n_160),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_168),
.B(n_172),
.Y(n_180)
);

OAI221xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_170),
.B1(n_159),
.B2(n_165),
.C(n_78),
.Y(n_181)
);


endmodule