module fake_netlist_1_7054_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
BUFx10_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_3), .Y(n_8) );
OAI22xp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_5), .B1(n_2), .B2(n_1), .Y(n_9) );
A2O1A1Ixp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B(n_7), .C(n_1), .Y(n_10) );
AOI32xp33_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_8), .A3(n_7), .B1(n_1), .B2(n_0), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_2), .Y(n_12) );
AOI22xp33_ASAP7_75t_SL g13 ( .A1(n_12), .A2(n_11), .B1(n_0), .B2(n_1), .Y(n_13) );
endmodule