module fake_jpeg_25849_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_65),
.A2(n_96),
.B1(n_103),
.B2(n_45),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_37),
.B1(n_23),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_75),
.B(n_83),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_37),
.B1(n_42),
.B2(n_35),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_35),
.B1(n_33),
.B2(n_26),
.Y(n_77)
);

OR2x4_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_17),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_65),
.C(n_95),
.Y(n_120)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_26),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_33),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_22),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_18),
.B1(n_64),
.B2(n_24),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_18),
.B1(n_36),
.B2(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_18),
.B1(n_31),
.B2(n_28),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_30),
.B1(n_25),
.B2(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_22),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_21),
.B1(n_36),
.B2(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_27),
.B1(n_36),
.B2(n_25),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_22),
.A3(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_32),
.B1(n_29),
.B2(n_17),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_120),
.B1(n_129),
.B2(n_69),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_98),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_47),
.B(n_46),
.C(n_43),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_135),
.B(n_103),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_85),
.A2(n_25),
.B1(n_27),
.B2(n_15),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_97),
.B1(n_105),
.B2(n_67),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_47),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_133),
.C(n_70),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_94),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_47),
.B1(n_46),
.B2(n_20),
.Y(n_129)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_16),
.C(n_34),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_153),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_141),
.B(n_148),
.Y(n_181)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_149),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_130),
.B1(n_109),
.B2(n_118),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_102),
.B1(n_93),
.B2(n_67),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_106),
.B1(n_128),
.B2(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_147),
.B(n_157),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_15),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_96),
.B1(n_102),
.B2(n_69),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_156),
.B1(n_161),
.B2(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_34),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_66),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_66),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_114),
.B(n_20),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_160),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_109),
.C(n_123),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_20),
.B1(n_34),
.B2(n_32),
.Y(n_161)
);

CKINVDCx11_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_70),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_34),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_153),
.B1(n_131),
.B2(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_178),
.B1(n_184),
.B2(n_191),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_107),
.C(n_135),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_4),
.C(n_5),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_123),
.B1(n_126),
.B2(n_137),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_116),
.B(n_125),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_170),
.B(n_177),
.C(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_113),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_121),
.B1(n_113),
.B2(n_116),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_116),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_117),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_188),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_126),
.B1(n_137),
.B2(n_44),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_110),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_133),
.B1(n_116),
.B2(n_118),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_148),
.B1(n_164),
.B2(n_161),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_117),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_160),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_32),
.C(n_29),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_140),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_204),
.C(n_210),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_143),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_145),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_217),
.B(n_221),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_174),
.B1(n_186),
.B2(n_187),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_173),
.B(n_143),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_216),
.B1(n_227),
.B2(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_14),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_0),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_2),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_4),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_5),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_212),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_166),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_233),
.A2(n_171),
.B(n_227),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_184),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_237),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_175),
.A3(n_168),
.B1(n_196),
.B2(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_191),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_187),
.B1(n_181),
.B2(n_167),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_181),
.B1(n_193),
.B2(n_183),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_179),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_168),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_204),
.C(n_200),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_264),
.C(n_256),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_256),
.B(n_252),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_214),
.B1(n_176),
.B2(n_210),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_233),
.B1(n_237),
.B2(n_236),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_220),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_265),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_268),
.B1(n_240),
.B2(n_235),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_218),
.C(n_245),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_178),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_202),
.B1(n_208),
.B2(n_216),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_275),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_171),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_235),
.B(n_233),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_243),
.B1(n_233),
.B2(n_236),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_251),
.B1(n_246),
.B2(n_259),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_283),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

OAI22x1_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_238),
.B1(n_273),
.B2(n_268),
.Y(n_282)
);

AOI22x1_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_267),
.B1(n_274),
.B2(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_234),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_248),
.B1(n_241),
.B2(n_230),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_246),
.C(n_250),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_230),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_6),
.C(n_8),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_294),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_257),
.B(n_232),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_305),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_276),
.Y(n_315)
);

OAI322xp33_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_259),
.A3(n_232),
.B1(n_169),
.B2(n_263),
.C1(n_272),
.C2(n_5),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_10),
.B(n_11),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_295),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_309),
.B(n_310),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_286),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_290),
.C(n_283),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_313),
.C(n_293),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_299),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.Y(n_323)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_308),
.C(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_321),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_296),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_301),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_326),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_310),
.C(n_292),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_297),
.B(n_298),
.Y(n_326)
);

INVx11_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_277),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_316),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_328),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.C(n_329),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_330),
.B(n_331),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_327),
.B1(n_281),
.B2(n_304),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_304),
.B(n_305),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_300),
.Y(n_341)
);


endmodule