module fake_jpeg_26036_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_22),
.B1(n_36),
.B2(n_38),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_59),
.Y(n_83)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_86),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

AOI22x1_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_81),
.B1(n_89),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_22),
.B1(n_23),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_92),
.B1(n_30),
.B2(n_35),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_45),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_32),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_28),
.B(n_45),
.Y(n_128)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_84),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_18),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_48),
.B1(n_44),
.B2(n_23),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_30),
.B1(n_24),
.B2(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_24),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_23),
.B1(n_30),
.B2(n_36),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_93),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_29),
.B1(n_20),
.B2(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_97),
.B1(n_73),
.B2(n_69),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_127),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_83),
.B1(n_89),
.B2(n_81),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_21),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_13),
.B(n_14),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_31),
.B(n_27),
.C(n_28),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_21),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_135),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_67),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_110),
.B1(n_100),
.B2(n_107),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_138),
.B1(n_100),
.B2(n_107),
.Y(n_174)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_143),
.Y(n_165)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_109),
.B1(n_101),
.B2(n_124),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_90),
.B1(n_82),
.B2(n_95),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_91),
.B1(n_120),
.B2(n_34),
.Y(n_188)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_75),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_145),
.C(n_112),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_147),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_17),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_154),
.B(n_80),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_21),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_34),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_104),
.B(n_112),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_160),
.B(n_180),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_145),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_127),
.B(n_117),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_121),
.A3(n_103),
.B1(n_99),
.B2(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_179),
.B1(n_149),
.B2(n_130),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_34),
.Y(n_212)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_176),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_129),
.C(n_113),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_150),
.C(n_139),
.Y(n_196)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_172),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_188),
.B1(n_135),
.B2(n_137),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_113),
.B1(n_122),
.B2(n_100),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_177),
.B1(n_136),
.B2(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_122),
.B1(n_118),
.B2(n_91),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_184),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_17),
.B1(n_26),
.B2(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_108),
.B(n_115),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_21),
.B(n_115),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_154),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_189),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_203),
.B(n_209),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_154),
.B(n_143),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_193),
.A2(n_200),
.B(n_208),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_196),
.C(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_206),
.B1(n_214),
.B2(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_198),
.B(n_204),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_152),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_152),
.B(n_151),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_211),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_163),
.A2(n_120),
.B(n_21),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_26),
.B(n_17),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_217),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_26),
.B(n_17),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_219),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_34),
.B1(n_26),
.B2(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_170),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_2),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_0),
.B(n_2),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_8),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_167),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_229),
.B1(n_235),
.B2(n_236),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_239),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_243),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_184),
.B1(n_176),
.B2(n_169),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_171),
.C(n_168),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_185),
.B1(n_164),
.B2(n_167),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_162),
.B1(n_177),
.B2(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_240),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_200),
.B1(n_198),
.B2(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_202),
.B1(n_214),
.B2(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_209),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_220),
.C(n_212),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_190),
.C(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_193),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_265),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_203),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_253),
.A2(n_224),
.B1(n_227),
.B2(n_219),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_267),
.Y(n_286)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.Y(n_280)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_238),
.B(n_162),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_222),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_190),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_231),
.B(n_217),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_269),
.Y(n_284)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_230),
.C(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_274),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_245),
.C(n_234),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_240),
.C(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_277),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_237),
.C(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_225),
.B1(n_242),
.B2(n_226),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_283),
.B1(n_253),
.B2(n_254),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_247),
.C(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_281),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_222),
.B1(n_246),
.B2(n_172),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_288),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_250),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_249),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_266),
.B1(n_263),
.B2(n_218),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_263),
.B1(n_266),
.B2(n_222),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_272),
.B1(n_277),
.B2(n_287),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_9),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_9),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_8),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_6),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_8),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_6),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_280),
.C(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_308),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_10),
.CI(n_15),
.CON(n_307),
.SN(n_307)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_315),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_7),
.B(n_15),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_303),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_323),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_301),
.C(n_299),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_311),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_290),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_304),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_311),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_307),
.B1(n_315),
.B2(n_313),
.Y(n_329)
);

AOI21x1_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_330),
.B(n_324),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_327),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_317),
.B(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_331),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_328),
.B(n_323),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_300),
.B1(n_293),
.B2(n_14),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_12),
.B(n_16),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_3),
.B(n_4),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_5),
.C(n_3),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_4),
.C(n_5),
.Y(n_341)
);


endmodule