module fake_jpeg_27473_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_47),
.B1(n_30),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_34),
.B1(n_17),
.B2(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_34),
.B1(n_17),
.B2(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_70),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_0),
.B(n_2),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_42),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_16),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_29),
.B1(n_33),
.B2(n_25),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_45),
.B1(n_66),
.B2(n_33),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_33),
.B1(n_25),
.B2(n_19),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_19),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_98),
.C(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_69),
.C(n_71),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_25),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_91),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_16),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_108),
.Y(n_141)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_56),
.C(n_54),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_80),
.B1(n_79),
.B2(n_86),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_62),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_121),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_76),
.B(n_74),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_127),
.B(n_73),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_77),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_91),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_135),
.B(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_82),
.B1(n_51),
.B2(n_52),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_98),
.B1(n_93),
.B2(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_90),
.B1(n_52),
.B2(n_45),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_126),
.B1(n_139),
.B2(n_73),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_51),
.B1(n_49),
.B2(n_80),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_84),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_100),
.Y(n_154)
);

NAND2x1_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_92),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_144),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_156),
.B1(n_122),
.B2(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_147),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_163),
.B(n_117),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_167),
.B1(n_125),
.B2(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_157),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_103),
.B1(n_112),
.B2(n_49),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_105),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_135),
.B(n_131),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_178),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_119),
.B(n_130),
.C(n_138),
.D(n_121),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_180),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_149),
.C(n_159),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_124),
.B1(n_80),
.B2(n_85),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_124),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_132),
.B(n_134),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_4),
.B(n_5),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_62),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_167),
.B1(n_147),
.B2(n_146),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_198),
.B1(n_201),
.B2(n_179),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_144),
.B1(n_155),
.B2(n_153),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_134),
.A3(n_161),
.B1(n_165),
.B2(n_156),
.C1(n_143),
.C2(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_151),
.B1(n_166),
.B2(n_99),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_207),
.B(n_177),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_192),
.B1(n_196),
.B2(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_209),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_169),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_6),
.C(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_173),
.C(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_213),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_194),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_217),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_175),
.B(n_189),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_219),
.B(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_192),
.B1(n_195),
.B2(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_178),
.C(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_219),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_193),
.C(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_176),
.Y(n_240)
);

AOI31xp67_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_232),
.A3(n_209),
.B(n_199),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_246),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_224),
.C(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_227),
.B1(n_229),
.B2(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_252),
.B1(n_8),
.B2(n_9),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_234),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_9),
.B(n_10),
.Y(n_260)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_6),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_260),
.B(n_11),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_7),
.C(n_8),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_265),
.C(n_263),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_256),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_258),
.C(n_265),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_266),
.B1(n_14),
.B2(n_15),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_12),
.Y(n_270)
);


endmodule