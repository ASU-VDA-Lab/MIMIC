module real_aes_12262_n_5 (n_4, n_0, n_3, n_2, n_1, n_5);
input n_4;
input n_0;
input n_3;
input n_2;
input n_1;
output n_5;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_6;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
NAND3xp33_ASAP7_75t_SL g6 ( .A(n_0), .B(n_7), .C(n_9), .Y(n_6) );
BUFx3_ASAP7_75t_L g23 ( .A(n_1), .Y(n_23) );
BUFx2_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
AOI31xp33_ASAP7_75t_L g5 ( .A1(n_6), .A2(n_16), .A3(n_18), .B(n_24), .Y(n_5) );
INVx1_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
INVx1_ASAP7_75t_SL g9 ( .A(n_10), .Y(n_9) );
INVx1_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
INVx5_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
BUFx8_ASAP7_75t_SL g12 ( .A(n_13), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_16), .B(n_18), .Y(n_24) );
INVx1_ASAP7_75t_SL g16 ( .A(n_17), .Y(n_16) );
INVxp67_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
endmodule