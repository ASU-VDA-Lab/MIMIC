module real_aes_4827_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_287;
wire n_905;
wire n_503;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_0), .A2(n_22), .B1(n_321), .B2(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_1), .A2(n_69), .B1(n_341), .B2(n_346), .Y(n_340) );
INVx1_ASAP7_75t_SL g402 ( .A(n_2), .Y(n_402) );
INVx1_ASAP7_75t_L g464 ( .A(n_3), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_3), .A2(n_111), .B1(n_709), .B2(n_730), .Y(n_742) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_4), .Y(n_687) );
AND2x4_ASAP7_75t_L g697 ( .A(n_4), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g706 ( .A(n_4), .B(n_242), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_5), .A2(n_72), .B1(n_594), .B2(n_597), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_6), .A2(n_144), .B1(n_385), .B2(n_388), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_7), .A2(n_83), .B1(n_672), .B2(n_945), .Y(n_944) );
AOI21xp33_ASAP7_75t_SL g470 ( .A1(n_8), .A2(n_310), .B(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_9), .A2(n_232), .B1(n_376), .B2(n_377), .Y(n_634) );
INVx1_ASAP7_75t_L g419 ( .A(n_10), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_11), .A2(n_27), .B1(n_338), .B2(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_12), .A2(n_195), .B1(n_351), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_13), .A2(n_215), .B1(n_379), .B2(n_380), .Y(n_633) );
INVx1_ASAP7_75t_L g534 ( .A(n_14), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_15), .A2(n_29), .B1(n_504), .B2(n_583), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_16), .Y(n_707) );
INVxp33_ASAP7_75t_SL g723 ( .A(n_17), .Y(n_723) );
AO22x1_ASAP7_75t_L g644 ( .A1(n_18), .A2(n_131), .B1(n_393), .B2(n_394), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_19), .A2(n_127), .B1(n_600), .B2(n_667), .Y(n_666) );
AO22x2_ASAP7_75t_L g762 ( .A1(n_20), .A2(n_64), .B1(n_709), .B2(n_730), .Y(n_762) );
AO22x1_ASAP7_75t_L g763 ( .A1(n_21), .A2(n_248), .B1(n_735), .B2(n_741), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_23), .A2(n_46), .B1(n_321), .B2(n_454), .Y(n_940) );
INVx1_ASAP7_75t_L g674 ( .A(n_24), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_25), .A2(n_123), .B1(n_376), .B2(n_377), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_26), .A2(n_58), .B1(n_376), .B2(n_380), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_28), .A2(n_91), .B1(n_373), .B2(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g523 ( .A(n_30), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_31), .A2(n_108), .B1(n_705), .B2(n_728), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_32), .A2(n_373), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g280 ( .A(n_33), .Y(n_280) );
INVxp67_ASAP7_75t_L g293 ( .A(n_33), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_33), .B(n_181), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_34), .A2(n_191), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_35), .A2(n_202), .B1(n_699), .B2(n_709), .Y(n_768) );
AOI21xp33_ASAP7_75t_SL g566 ( .A1(n_36), .A2(n_567), .B(n_569), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_37), .A2(n_110), .B1(n_735), .B2(n_737), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_38), .B(n_475), .Y(n_474) );
AO22x1_ASAP7_75t_L g642 ( .A1(n_39), .A2(n_122), .B1(n_387), .B2(n_391), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_40), .A2(n_67), .B1(n_384), .B2(n_385), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_41), .B(n_265), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_42), .A2(n_241), .B1(n_330), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_43), .A2(n_228), .B1(n_661), .B2(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g911 ( .A(n_44), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_45), .A2(n_105), .B1(n_357), .B2(n_360), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_47), .A2(n_78), .B1(n_376), .B2(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_48), .A2(n_182), .B1(n_454), .B2(n_477), .Y(n_476) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_49), .B(n_538), .Y(n_537) );
OAI22x1_ASAP7_75t_L g587 ( .A1(n_50), .A2(n_588), .B1(n_621), .B2(n_622), .Y(n_587) );
INVx1_ASAP7_75t_L g622 ( .A(n_50), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_51), .A2(n_219), .B1(n_730), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_52), .A2(n_231), .B1(n_320), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_53), .A2(n_136), .B1(n_337), .B2(n_346), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_54), .B(n_374), .Y(n_632) );
INVx1_ASAP7_75t_L g520 ( .A(n_55), .Y(n_520) );
INVx2_ASAP7_75t_L g685 ( .A(n_56), .Y(n_685) );
INVxp33_ASAP7_75t_SL g710 ( .A(n_57), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_59), .A2(n_155), .B1(n_347), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_60), .A2(n_193), .B1(n_325), .B2(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_61), .A2(n_210), .B1(n_610), .B2(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g424 ( .A(n_62), .Y(n_424) );
INVx1_ASAP7_75t_L g696 ( .A(n_63), .Y(n_696) );
AND2x4_ASAP7_75t_L g702 ( .A(n_63), .B(n_685), .Y(n_702) );
INVx1_ASAP7_75t_SL g736 ( .A(n_63), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_65), .A2(n_165), .B1(n_442), .B2(n_483), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_66), .A2(n_188), .B1(n_393), .B2(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_68), .B(n_258), .Y(n_512) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_70), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_71), .A2(n_133), .B1(n_379), .B2(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g550 ( .A(n_73), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_74), .A2(n_171), .B1(n_379), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_75), .A2(n_84), .B1(n_613), .B2(n_615), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_76), .A2(n_82), .B1(n_315), .B2(n_522), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_77), .A2(n_178), .B1(n_449), .B2(n_671), .C(n_673), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_79), .A2(n_218), .B1(n_442), .B2(n_443), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_80), .B(n_380), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_81), .A2(n_209), .B1(n_358), .B2(n_480), .Y(n_935) );
AO22x1_ASAP7_75t_L g283 ( .A1(n_85), .A2(n_170), .B1(n_284), .B2(n_295), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_86), .A2(n_197), .B1(n_480), .B2(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g266 ( .A(n_87), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_87), .B(n_180), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_88), .A2(n_204), .B1(n_338), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_89), .A2(n_94), .B1(n_342), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_90), .A2(n_217), .B1(n_309), .B2(n_314), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_92), .A2(n_128), .B1(n_709), .B2(n_730), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_93), .A2(n_138), .B1(n_486), .B2(n_487), .Y(n_485) );
AO221x2_ASAP7_75t_L g691 ( .A1(n_95), .A2(n_97), .B1(n_692), .B2(n_699), .C(n_703), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_96), .A2(n_233), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_98), .A2(n_247), .B1(n_694), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g637 ( .A(n_99), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_100), .B(n_450), .Y(n_528) );
XOR2x2_ASAP7_75t_L g252 ( .A(n_101), .B(n_253), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_102), .A2(n_160), .B1(n_384), .B2(n_390), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_103), .A2(n_157), .B1(n_351), .B2(n_507), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_104), .A2(n_239), .B1(n_387), .B2(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g472 ( .A(n_106), .Y(n_472) );
INVx1_ASAP7_75t_L g460 ( .A(n_107), .Y(n_460) );
XNOR2x1_ASAP7_75t_L g434 ( .A(n_108), .B(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_109), .A2(n_158), .B1(n_351), .B2(n_446), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_112), .A2(n_220), .B1(n_651), .B2(n_653), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_113), .A2(n_120), .B1(n_354), .B2(n_506), .Y(n_578) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_114), .A2(n_238), .B1(n_384), .B2(n_390), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_115), .A2(n_216), .B1(n_390), .B2(n_391), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_116), .A2(n_190), .B1(n_384), .B2(n_385), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_117), .A2(n_187), .B1(n_387), .B2(n_391), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_118), .A2(n_194), .B1(n_735), .B2(n_737), .Y(n_734) );
XOR2x2_ASAP7_75t_L g904 ( .A(n_118), .B(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_118), .A2(n_927), .B1(n_929), .B2(n_946), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_119), .A2(n_208), .B1(n_330), .B2(n_358), .Y(n_437) );
INVx1_ASAP7_75t_L g421 ( .A(n_121), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_124), .A2(n_130), .B1(n_315), .B2(n_522), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_125), .A2(n_256), .B(n_283), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_126), .A2(n_149), .B1(n_351), .B2(n_353), .Y(n_350) );
XOR2xp5_ASAP7_75t_L g929 ( .A(n_129), .B(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_132), .A2(n_141), .B1(n_347), .B2(n_481), .Y(n_934) );
AOI22x1_ASAP7_75t_L g646 ( .A1(n_134), .A2(n_647), .B1(n_648), .B2(n_675), .Y(n_646) );
INVx1_ASAP7_75t_L g675 ( .A(n_134), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_135), .A2(n_150), .B1(n_385), .B2(n_388), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_137), .B(n_565), .Y(n_564) );
CKINVDCx14_ASAP7_75t_R g368 ( .A(n_139), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_140), .A2(n_148), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_142), .A2(n_185), .B1(n_342), .B2(n_509), .Y(n_508) );
XNOR2x2_ASAP7_75t_L g629 ( .A(n_143), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_145), .B(n_295), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_146), .A2(n_173), .B1(n_694), .B2(n_705), .Y(n_769) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_147), .A2(n_169), .B1(n_320), .B2(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g417 ( .A(n_151), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_152), .A2(n_222), .B1(n_342), .B2(n_439), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_153), .A2(n_196), .B1(n_456), .B2(n_458), .C(n_459), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_154), .A2(n_226), .B1(n_387), .B2(n_391), .Y(n_410) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_156), .A2(n_181), .B1(n_265), .B2(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g307 ( .A(n_156), .Y(n_307) );
AOI21xp5_ASAP7_75t_SL g415 ( .A1(n_159), .A2(n_373), .B(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_161), .A2(n_183), .B1(n_393), .B2(n_394), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_162), .A2(n_179), .B1(n_450), .B2(n_477), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_163), .A2(n_235), .B1(n_483), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_164), .A2(n_166), .B1(n_393), .B2(n_394), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_167), .A2(n_221), .B1(n_329), .B2(n_337), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_168), .A2(n_234), .B1(n_390), .B2(n_391), .Y(n_913) );
INVx1_ASAP7_75t_L g719 ( .A(n_172), .Y(n_719) );
INVx1_ASAP7_75t_L g570 ( .A(n_174), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_175), .A2(n_211), .B1(n_379), .B2(n_919), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_176), .A2(n_212), .B1(n_338), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_177), .A2(n_200), .B1(n_694), .B2(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g282 ( .A(n_180), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_180), .B(n_304), .Y(n_303) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_181), .A2(n_206), .B(n_294), .Y(n_318) );
INVx1_ASAP7_75t_L g413 ( .A(n_184), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_186), .A2(n_227), .B1(n_385), .B2(n_388), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_189), .A2(n_201), .B1(n_393), .B2(n_394), .Y(n_546) );
INVx1_ASAP7_75t_L g526 ( .A(n_192), .Y(n_526) );
INVx1_ASAP7_75t_L g516 ( .A(n_198), .Y(n_516) );
INVx1_ASAP7_75t_L g561 ( .A(n_199), .Y(n_561) );
INVx1_ASAP7_75t_SL g529 ( .A(n_203), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_205), .A2(n_245), .B1(n_384), .B2(n_390), .Y(n_547) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_206), .B(n_236), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_207), .A2(n_244), .B1(n_907), .B2(n_909), .C(n_910), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_213), .A2(n_223), .B1(n_452), .B2(n_454), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_214), .A2(n_243), .B1(n_600), .B2(n_601), .C(n_602), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_224), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_225), .A2(n_237), .B1(n_342), .B2(n_662), .Y(n_937) );
AOI21xp33_ASAP7_75t_SL g548 ( .A1(n_229), .A2(n_373), .B(n_549), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_230), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_236), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_240), .B(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g698 ( .A(n_242), .Y(n_698) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_242), .Y(n_949) );
INVx1_ASAP7_75t_L g603 ( .A(n_246), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_429), .B(n_679), .C(n_688), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_250), .A2(n_429), .B(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_364), .B1(n_427), .B2(n_428), .Y(n_250) );
BUFx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g427 ( .A(n_252), .Y(n_427) );
NOR2x1_ASAP7_75t_L g253 ( .A(n_254), .B(n_327), .Y(n_253) );
NAND3xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_308), .C(n_319), .Y(n_254) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g475 ( .A(n_259), .Y(n_475) );
INVx2_ASAP7_75t_L g565 ( .A(n_259), .Y(n_565) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g672 ( .A(n_261), .Y(n_672) );
INVx3_ASAP7_75t_L g908 ( .A(n_261), .Y(n_908) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
AND2x2_ASAP7_75t_L g326 ( .A(n_262), .B(n_323), .Y(n_326) );
AND2x2_ASAP7_75t_L g343 ( .A(n_262), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g348 ( .A(n_262), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g374 ( .A(n_262), .B(n_271), .Y(n_374) );
AND2x4_ASAP7_75t_L g379 ( .A(n_262), .B(n_323), .Y(n_379) );
AND2x4_ASAP7_75t_L g387 ( .A(n_262), .B(n_344), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_262), .B(n_334), .Y(n_388) );
AND2x2_ASAP7_75t_L g484 ( .A(n_262), .B(n_344), .Y(n_484) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g313 ( .A(n_263), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
INVx1_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_266), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_268), .A2(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g291 ( .A(n_270), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g333 ( .A(n_270), .Y(n_333) );
AND2x4_ASAP7_75t_L g311 ( .A(n_271), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g316 ( .A(n_271), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g355 ( .A(n_271), .B(n_332), .Y(n_355) );
AND2x2_ASAP7_75t_L g373 ( .A(n_271), .B(n_312), .Y(n_373) );
AND2x4_ASAP7_75t_L g377 ( .A(n_271), .B(n_317), .Y(n_377) );
AND2x4_ASAP7_75t_L g394 ( .A(n_271), .B(n_332), .Y(n_394) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_277), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_273), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g323 ( .A(n_273), .B(n_277), .Y(n_323) );
OR2x2_ASAP7_75t_L g335 ( .A(n_273), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g344 ( .A(n_273), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_276), .B(n_303), .C(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx4_ASAP7_75t_L g450 ( .A(n_285), .Y(n_450) );
INVx2_ASAP7_75t_L g575 ( .A(n_285), .Y(n_575) );
INVx3_ASAP7_75t_L g600 ( .A(n_285), .Y(n_600) );
INVx5_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g469 ( .A(n_286), .Y(n_469) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
AND2x4_ASAP7_75t_L g380 ( .A(n_287), .B(n_291), .Y(n_380) );
AND2x2_ASAP7_75t_L g919 ( .A(n_287), .B(n_291), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
INVx2_ASAP7_75t_SL g461 ( .A(n_295), .Y(n_461) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_296), .B(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_296), .Y(n_473) );
INVx1_ASAP7_75t_L g518 ( .A(n_296), .Y(n_518) );
INVx2_ASAP7_75t_L g572 ( .A(n_296), .Y(n_572) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx3_ASAP7_75t_L g605 ( .A(n_297), .Y(n_605) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .Y(n_297) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_299), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_304), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g317 ( .A(n_305), .B(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g457 ( .A(n_311), .Y(n_457) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_311), .Y(n_596) );
INVx2_ASAP7_75t_L g943 ( .A(n_311), .Y(n_943) );
AND2x4_ASAP7_75t_L g322 ( .A(n_312), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g376 ( .A(n_312), .B(n_323), .Y(n_376) );
AND2x4_ASAP7_75t_L g332 ( .A(n_313), .B(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx4_ASAP7_75t_L g524 ( .A(n_315), .Y(n_524) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_316), .Y(n_454) );
INVx3_ASAP7_75t_L g598 ( .A(n_316), .Y(n_598) );
AND2x4_ASAP7_75t_L g339 ( .A(n_317), .B(n_334), .Y(n_339) );
AND2x4_ASAP7_75t_L g363 ( .A(n_317), .B(n_344), .Y(n_363) );
AND2x4_ASAP7_75t_L g385 ( .A(n_317), .B(n_334), .Y(n_385) );
AND2x4_ASAP7_75t_L g391 ( .A(n_317), .B(n_344), .Y(n_391) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g449 ( .A(n_322), .Y(n_449) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_322), .Y(n_514) );
INVx1_ASAP7_75t_L g568 ( .A(n_322), .Y(n_568) );
AND2x4_ASAP7_75t_L g352 ( .A(n_323), .B(n_332), .Y(n_352) );
AND2x4_ASAP7_75t_L g393 ( .A(n_323), .B(n_332), .Y(n_393) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g453 ( .A(n_326), .Y(n_453) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_326), .Y(n_477) );
NAND4xp25_ASAP7_75t_SL g327 ( .A(n_328), .B(n_340), .C(n_350), .D(n_356), .Y(n_327) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_331), .Y(n_480) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_331), .Y(n_583) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x4_ASAP7_75t_L g359 ( .A(n_332), .B(n_344), .Y(n_359) );
AND2x4_ASAP7_75t_L g384 ( .A(n_332), .B(n_349), .Y(n_384) );
AND2x4_ASAP7_75t_L g390 ( .A(n_332), .B(n_344), .Y(n_390) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g349 ( .A(n_335), .Y(n_349) );
INVx1_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
BUFx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx6_ASAP7_75t_L g444 ( .A(n_339), .Y(n_444) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx8_ASAP7_75t_L g661 ( .A(n_343), .Y(n_661) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx12f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_348), .Y(n_502) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_348), .Y(n_585) );
BUFx3_ASAP7_75t_L g664 ( .A(n_348), .Y(n_664) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_352), .Y(n_506) );
INVx3_ASAP7_75t_L g614 ( .A(n_352), .Y(n_614) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx5_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g446 ( .A(n_355), .Y(n_446) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_355), .Y(n_507) );
INVx1_ASAP7_75t_L g656 ( .A(n_355), .Y(n_656) );
BUFx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_359), .Y(n_486) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_359), .Y(n_504) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx4_ASAP7_75t_L g439 ( .A(n_362), .Y(n_439) );
INVx1_ASAP7_75t_L g487 ( .A(n_362), .Y(n_487) );
INVx4_ASAP7_75t_L g509 ( .A(n_362), .Y(n_509) );
INVx2_ASAP7_75t_L g580 ( .A(n_362), .Y(n_580) );
INVx1_ASAP7_75t_L g619 ( .A(n_362), .Y(n_619) );
INVx4_ASAP7_75t_L g662 ( .A(n_362), .Y(n_662) );
INVx8_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g428 ( .A(n_364), .Y(n_428) );
OAI22xp33_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_366), .B1(n_398), .B2(n_399), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_395), .Y(n_367) );
NAND3xp33_ASAP7_75t_SL g395 ( .A(n_368), .B(n_396), .C(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_382), .Y(n_370) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g371 ( .A(n_372), .B(n_375), .C(n_378), .D(n_381), .Y(n_371) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_373), .Y(n_909) );
INVx2_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_374), .Y(n_538) );
INVx2_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
INVx2_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVxp67_ASAP7_75t_L g396 ( .A(n_382), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .C(n_389), .D(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_411), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_418), .C(n_423), .Y(n_411) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_415), .Y(n_412) );
INVx2_ASAP7_75t_L g458 ( .A(n_414), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_418) );
INVxp67_ASAP7_75t_L g540 ( .A(n_422), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .B(n_426), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_555), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_495), .B1(n_553), .B2(n_554), .Y(n_430) );
INVx2_ASAP7_75t_L g553 ( .A(n_431), .Y(n_553) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
XNOR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_462), .Y(n_433) );
NAND4xp75_ASAP7_75t_L g435 ( .A(n_436), .B(n_440), .C(n_447), .D(n_455), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g481 ( .A(n_444), .Y(n_481) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_453), .Y(n_668) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_SL g522 ( .A(n_457), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI21x1_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_489), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_463), .B(n_476), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_466), .B(n_478), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_474), .C(n_476), .Y(n_466) );
INVx1_ASAP7_75t_L g493 ( .A(n_467), .Y(n_493) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_473), .B(n_550), .Y(n_549) );
INVxp67_ASAP7_75t_L g491 ( .A(n_474), .Y(n_491) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_475), .Y(n_601) );
INVx3_ASAP7_75t_L g527 ( .A(n_477), .Y(n_527) );
BUFx3_ASAP7_75t_L g592 ( .A(n_477), .Y(n_592) );
INVx1_ASAP7_75t_L g494 ( .A(n_478), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .C(n_485), .D(n_488), .Y(n_478) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_486), .Y(n_609) );
BUFx12f_ASAP7_75t_L g658 ( .A(n_486), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_530), .B1(n_551), .B2(n_552), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
XOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_529), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
AND4x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_505), .D(n_508), .Y(n_500) );
BUFx2_ASAP7_75t_SL g615 ( .A(n_507), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .C(n_525), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_512), .B(n_513), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_523), .B2(n_524), .Y(n_519) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_529), .A2(n_704), .B1(n_708), .B2(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g552 ( .A(n_530), .Y(n_552) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
XNOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .C(n_541), .Y(n_536) );
NAND4xp25_ASAP7_75t_SL g542 ( .A(n_543), .B(n_544), .C(n_545), .D(n_548), .Y(n_542) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_626), .B1(n_677), .B2(n_678), .Y(n_555) );
INVx1_ASAP7_75t_L g677 ( .A(n_556), .Y(n_677) );
AO22x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_586), .B1(n_623), .B2(n_624), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g625 ( .A(n_560), .Y(n_625) );
XNOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NOR4xp75_ASAP7_75t_L g562 ( .A(n_563), .B(n_573), .C(n_577), .D(n_581), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g611 ( .A(n_583), .Y(n_611) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g623 ( .A(n_587), .Y(n_623) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_606), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_589), .B(n_606), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_599), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_604), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx4_ASAP7_75t_L g638 ( .A(n_605), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_607), .B(n_616), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g652 ( .A(n_614), .Y(n_652) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g678 ( .A(n_626), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_645), .B2(n_676), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_639), .Y(n_630) );
AND4x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .C(n_634), .D(n_635), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_638), .B(n_911), .Y(n_910) );
INVx4_ASAP7_75t_L g945 ( .A(n_638), .Y(n_945) );
NOR4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .C(n_643), .D(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g676 ( .A(n_645), .Y(n_676) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND4xp75_ASAP7_75t_L g648 ( .A(n_649), .B(n_659), .C(n_665), .D(n_670), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_657), .Y(n_649) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_686), .C(n_687), .Y(n_682) );
AND2x2_ASAP7_75t_L g923 ( .A(n_683), .B(n_924), .Y(n_923) );
AND2x2_ASAP7_75t_L g928 ( .A(n_683), .B(n_925), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_683), .A2(n_687), .B(n_736), .Y(n_950) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AO21x1_ASAP7_75t_L g947 ( .A1(n_684), .A2(n_948), .B(n_950), .Y(n_947) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g695 ( .A(n_685), .B(n_696), .Y(n_695) );
AND3x4_ASAP7_75t_L g735 ( .A(n_685), .B(n_697), .C(n_736), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_686), .B(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_687), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_898), .B1(n_900), .B2(n_921), .C(n_926), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_711), .B(n_817), .C(n_868), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_690), .A2(n_818), .B(n_850), .Y(n_817) );
INVx1_ASAP7_75t_L g886 ( .A(n_690), .Y(n_886) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI311xp33_ASAP7_75t_L g850 ( .A1(n_691), .A2(n_851), .A3(n_859), .B(n_861), .C(n_864), .Y(n_850) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_693), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_720) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
AND2x4_ASAP7_75t_L g705 ( .A(n_695), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g737 ( .A(n_695), .B(n_706), .Y(n_737) );
AND2x2_ASAP7_75t_L g741 ( .A(n_695), .B(n_706), .Y(n_741) );
AND2x4_ASAP7_75t_L g701 ( .A(n_697), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_697), .B(n_702), .Y(n_722) );
AND2x4_ASAP7_75t_L g730 ( .A(n_697), .B(n_702), .Y(n_730) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g709 ( .A(n_702), .B(n_706), .Y(n_709) );
AND2x2_ASAP7_75t_L g728 ( .A(n_702), .B(n_706), .Y(n_728) );
AND2x2_ASAP7_75t_L g746 ( .A(n_702), .B(n_706), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B1(n_708), .B2(n_710), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g899 ( .A(n_705), .Y(n_899) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND5xp2_ASAP7_75t_L g711 ( .A(n_712), .B(n_748), .C(n_757), .D(n_789), .E(n_810), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_743), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_724), .Y(n_715) );
AND2x2_ASAP7_75t_L g758 ( .A(n_716), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g776 ( .A(n_716), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_716), .B(n_726), .Y(n_793) );
AND2x2_ASAP7_75t_L g883 ( .A(n_716), .B(n_777), .Y(n_883) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_717), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g785 ( .A(n_717), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_717), .B(n_756), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_717), .B(n_744), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_717), .B(n_761), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_717), .B(n_788), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_717), .B(n_725), .Y(n_843) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_717), .Y(n_862) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_724), .A2(n_770), .B(n_785), .C(n_786), .Y(n_784) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_731), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_725), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_725), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g795 ( .A(n_725), .B(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g806 ( .A(n_725), .B(n_753), .Y(n_806) );
OR2x2_ASAP7_75t_L g830 ( .A(n_725), .B(n_732), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_725), .B(n_739), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_725), .B(n_753), .Y(n_875) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g782 ( .A(n_726), .B(n_739), .Y(n_782) );
INVx1_ASAP7_75t_L g800 ( .A(n_726), .Y(n_800) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_732), .B(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_739), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_733), .Y(n_753) );
AND2x2_ASAP7_75t_L g796 ( .A(n_733), .B(n_739), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_733), .A2(n_821), .B1(n_823), .B2(n_825), .Y(n_820) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
OR2x2_ASAP7_75t_L g752 ( .A(n_739), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g770 ( .A(n_739), .Y(n_770) );
AND2x2_ASAP7_75t_L g777 ( .A(n_739), .B(n_753), .Y(n_777) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_744), .Y(n_756) );
OR2x2_ASAP7_75t_L g760 ( .A(n_744), .B(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g780 ( .A(n_744), .Y(n_780) );
AND2x2_ASAP7_75t_L g788 ( .A(n_744), .B(n_761), .Y(n_788) );
AND2x4_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_750), .B(n_754), .Y(n_749) );
INVx1_ASAP7_75t_L g894 ( .A(n_750), .Y(n_894) );
INVx1_ASAP7_75t_L g773 ( .A(n_752), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_752), .B(n_843), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_753), .B(n_799), .Y(n_798) );
OAI222xp33_ASAP7_75t_L g790 ( .A1(n_754), .A2(n_786), .B1(n_791), .B2(n_794), .C1(n_797), .C2(n_801), .Y(n_790) );
OAI211xp5_ASAP7_75t_L g851 ( .A1(n_754), .A2(n_852), .B(n_854), .C(n_857), .Y(n_851) );
AND2x2_ASAP7_75t_L g890 ( .A(n_754), .B(n_766), .Y(n_890) );
AND3x1_ASAP7_75t_L g895 ( .A(n_754), .B(n_799), .C(n_883), .Y(n_895) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g840 ( .A(n_755), .Y(n_840) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g809 ( .A(n_756), .B(n_761), .Y(n_809) );
AOI311xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_764), .A3(n_770), .B(n_771), .C(n_781), .Y(n_757) );
AOI222xp33_ASAP7_75t_L g810 ( .A1(n_759), .A2(n_761), .B1(n_777), .B2(n_811), .C1(n_813), .C2(n_814), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_759), .A2(n_832), .B1(n_835), .B2(n_836), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_759), .A2(n_881), .B1(n_884), .B2(n_887), .C(n_891), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_759), .B(n_841), .Y(n_892) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g783 ( .A(n_760), .B(n_767), .Y(n_783) );
INVx1_ASAP7_75t_L g804 ( .A(n_761), .Y(n_804) );
CKINVDCx6p67_ASAP7_75t_R g827 ( .A(n_761), .Y(n_827) );
OR2x2_ASAP7_75t_L g860 ( .A(n_761), .B(n_766), .Y(n_860) );
OR2x6_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_764), .B(n_809), .Y(n_829) );
INVx3_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g789 ( .A1(n_765), .A2(n_790), .B1(n_799), .B2(n_802), .C1(n_805), .C2(n_807), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_765), .B(n_809), .Y(n_808) );
INVx5_ASAP7_75t_L g819 ( .A(n_765), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_765), .B(n_785), .Y(n_879) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g779 ( .A(n_766), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g845 ( .A(n_766), .B(n_803), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_766), .B(n_827), .Y(n_867) );
INVx3_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g802 ( .A(n_767), .B(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g863 ( .A(n_767), .B(n_787), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_770), .B(n_792), .Y(n_791) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g872 ( .A(n_772), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_773), .B(n_792), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_L g861 ( .A1(n_774), .A2(n_797), .B(n_862), .C(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_L g866 ( .A(n_775), .B(n_799), .Y(n_866) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_776), .B(n_805), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_776), .B(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g835 ( .A(n_777), .B(n_799), .Y(n_835) );
AND2x2_ASAP7_75t_L g841 ( .A(n_777), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g876 ( .A(n_777), .Y(n_876) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g826 ( .A(n_780), .B(n_827), .Y(n_826) );
OAI21xp5_ASAP7_75t_SL g781 ( .A1(n_782), .A2(n_783), .B(n_784), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_SL g864 ( .A1(n_782), .A2(n_855), .B(n_865), .C(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g873 ( .A(n_783), .Y(n_873) );
AND2x2_ASAP7_75t_L g813 ( .A(n_785), .B(n_796), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_785), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g855 ( .A(n_785), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_785), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_787), .B(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_795), .A2(n_836), .B(n_845), .Y(n_849) );
INVx1_ASAP7_75t_L g822 ( .A(n_796), .Y(n_822) );
AND2x2_ASAP7_75t_L g858 ( .A(n_796), .B(n_799), .Y(n_858) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_799), .B(n_883), .Y(n_882) );
INVx3_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g828 ( .A1(n_801), .A2(n_829), .B(n_830), .C(n_831), .Y(n_828) );
AOI211xp5_ASAP7_75t_L g869 ( .A1(n_802), .A2(n_811), .B(n_870), .C(n_874), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_803), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_806), .A2(n_808), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g897 ( .A1(n_809), .A2(n_846), .B(n_858), .Y(n_897) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI211xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B(n_828), .C(n_838), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_L g893 ( .A1(n_819), .A2(n_894), .B(n_895), .C(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g888 ( .A(n_826), .Y(n_888) );
INVx1_ASAP7_75t_L g856 ( .A(n_830), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND3xp33_ASAP7_75t_SL g838 ( .A(n_839), .B(n_844), .C(n_849), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_855), .B(n_858), .C(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_880), .C(n_893), .Y(n_868) );
INVxp67_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
AOI21xp33_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B(n_877), .Y(n_874) );
INVxp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
INVxp67_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_892), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_899), .Y(n_898) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
NAND3x1_ASAP7_75t_L g905 ( .A(n_906), .B(n_912), .C(n_915), .Y(n_905) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
AND2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
AND4x1_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .C(n_918), .D(n_920), .Y(n_915) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
BUFx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NOR2x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_938), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .C(n_936), .D(n_937), .Y(n_933) );
NAND4xp25_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .C(n_941), .D(n_944), .Y(n_938) );
INVx3_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
BUFx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_949), .Y(n_948) );
endmodule