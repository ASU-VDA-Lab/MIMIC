module fake_ariane_1315_n_38 (n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_4, n_38);

input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_4;

output n_38;

wire n_8;
wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_27;
wire n_29;
wire n_17;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_9;
wire n_11;
wire n_34;
wire n_26;
wire n_14;
wire n_36;
wire n_33;
wire n_19;
wire n_30;
wire n_31;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_35;
wire n_10;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_11),
.B1(n_8),
.B2(n_3),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

AOI33xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_16),
.A3(n_17),
.B1(n_4),
.B2(n_6),
.B3(n_0),
.Y(n_25)
);

OR2x6_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_17),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_15),
.B(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

AOI222xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_24),
.B1(n_14),
.B2(n_25),
.C1(n_31),
.C2(n_27),
.Y(n_33)
);

OAI221xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_26),
.B1(n_29),
.B2(n_14),
.C(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_29),
.B1(n_26),
.B2(n_6),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_36),
.C(n_26),
.Y(n_38)
);


endmodule