module fake_jpeg_12474_n_97 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_39),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_26),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_24),
.B(n_27),
.C(n_25),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_39),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_57),
.B1(n_46),
.B2(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_67),
.Y(n_76)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_1),
.B(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_44),
.B1(n_40),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_13),
.B1(n_21),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_67),
.B1(n_58),
.B2(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_4),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_73),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_12),
.C(n_18),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_72),
.C(n_78),
.Y(n_79)
);

INVxp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_4),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_74),
.B2(n_75),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_15),
.Y(n_90)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_81),
.B1(n_80),
.B2(n_85),
.C(n_5),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_87),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_8),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_14),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_16),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_17),
.C(n_22),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_6),
.Y(n_97)
);


endmodule