module fake_jpeg_14719_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_54),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_45),
.B1(n_42),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_59),
.B1(n_33),
.B2(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_53),
.B(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_35),
.B1(n_17),
.B2(n_25),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_68),
.B(n_31),
.C(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_32),
.B(n_30),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_70),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_91),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_42),
.B1(n_39),
.B2(n_25),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_77),
.B(n_78),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_22),
.C(n_39),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_76),
.B(n_82),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_42),
.B1(n_25),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_89),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_22),
.B1(n_20),
.B2(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_28),
.C(n_33),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_2),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_98),
.B(n_2),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_27),
.B(n_3),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_24),
.B1(n_21),
.B2(n_27),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_27),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_4),
.Y(n_157)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_16),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_16),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_4),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_86),
.B1(n_100),
.B2(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_135),
.B1(n_147),
.B2(n_155),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_83),
.B(n_97),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_134),
.A2(n_157),
.B(n_5),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_92),
.B1(n_77),
.B2(n_86),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_94),
.C(n_105),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_126),
.C(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_146),
.B1(n_109),
.B2(n_110),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_97),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_160),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_82),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_82),
.B1(n_79),
.B2(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_152),
.Y(n_173)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_72),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_130),
.B1(n_127),
.B2(n_111),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_5),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_15),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_177),
.B(n_185),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_180),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_113),
.A3(n_126),
.B1(n_118),
.B2(n_117),
.C1(n_15),
.C2(n_132),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_169),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_136),
.C(n_134),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_115),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_125),
.B1(n_114),
.B2(n_122),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_124),
.B1(n_72),
.B2(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_152),
.A3(n_138),
.B1(n_137),
.B2(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_121),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_116),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_137),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_195),
.C(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_138),
.B(n_147),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_202),
.B(n_163),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_133),
.B(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_202),
.B1(n_203),
.B2(n_186),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_129),
.C(n_124),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_218),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_171),
.B1(n_163),
.B2(n_175),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_219),
.B1(n_212),
.B2(n_204),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_200),
.B(n_188),
.Y(n_223)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_171),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_221),
.C(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_199),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_203),
.B1(n_198),
.B2(n_186),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_166),
.B1(n_178),
.B2(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_161),
.C(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_231),
.B(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_233),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_210),
.B1(n_220),
.B2(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_234),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_196),
.B(n_198),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_211),
.CI(n_207),
.CON(n_234),
.SN(n_234)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_238),
.B(n_228),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_221),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_190),
.B(n_180),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_240),
.A2(n_244),
.B(n_182),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_233),
.B(n_185),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_245),
.A2(n_251),
.B(n_235),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_229),
.C(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_250),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_209),
.B(n_234),
.C(n_224),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_167),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_224),
.B(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_12),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_254),
.B(n_255),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_218),
.B(n_167),
.Y(n_254)
);

OAI21x1_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_247),
.B(n_218),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_260),
.B(n_6),
.C(n_8),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_183),
.B1(n_129),
.B2(n_8),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_258),
.A2(n_6),
.B(n_7),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_9),
.Y(n_265)
);


endmodule