module fake_netlist_5_735_n_1274 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1274);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1274;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_252;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_94),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_128),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_41),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_61),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_25),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_54),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_35),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_95),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_91),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_117),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_85),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_71),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_100),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_27),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_59),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_12),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_53),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_73),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_29),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_90),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_171),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_83),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_24),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_106),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_55),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_21),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_74),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_69),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_77),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_5),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_167),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_44),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_152),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_177),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_148),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_64),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_88),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_38),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_175),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_136),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_140),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_25),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_176),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_143),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_103),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_46),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_62),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_108),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_52),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_96),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_124),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_43),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_112),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_170),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_133),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_149),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_42),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_155),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_19),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_35),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_6),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_245),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_217),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_224),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_193),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_241),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_231),
.B(n_0),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_233),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_200),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_191),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_219),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_220),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_301),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_248),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_254),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_264),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_211),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_225),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_301),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_195),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_225),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_195),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_227),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_196),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_213),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_186),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_196),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_R g347 ( 
.A(n_218),
.B(n_49),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_204),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_188),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_194),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_231),
.B(n_0),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_198),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_204),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_203),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_216),
.B(n_1),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_205),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_207),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_209),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_265),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_212),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_216),
.B(n_1),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_226),
.B(n_2),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_222),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_214),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_266),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_229),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_282),
.B(n_3),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_222),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_267),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_268),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_237),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_226),
.B(n_4),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_275),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_286),
.B(n_4),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_208),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_232),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_239),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_291),
.B(n_5),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_247),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_291),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_235),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_249),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_234),
.B(n_6),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_238),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_240),
.Y(n_395)
);

BUFx8_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_344),
.B(n_184),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

BUFx12f_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_253),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_315),
.A2(n_262),
.B(n_256),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_344),
.B(n_184),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_344),
.B(n_185),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_185),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_311),
.B(n_260),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_390),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_263),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_277),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_283),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_285),
.B(n_284),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_L g433 ( 
.A(n_309),
.B(n_289),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_317),
.B(n_187),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_322),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_352),
.B(n_354),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_305),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_382),
.A2(n_299),
.B1(n_303),
.B2(n_302),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_322),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_357),
.B(n_187),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_358),
.B(n_287),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_319),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_319),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_325),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

AND2x2_ASAP7_75t_SL g448 ( 
.A(n_393),
.B(n_222),
.Y(n_448)
);

AND3x2_ASAP7_75t_L g449 ( 
.A(n_355),
.B(n_304),
.C(n_290),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_334),
.B(n_189),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_310),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_325),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_320),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_359),
.B(n_222),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_326),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_321),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_326),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_321),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_347),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_361),
.B(n_243),
.Y(n_460)
);

CKINVDCx8_ASAP7_75t_R g461 ( 
.A(n_327),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_333),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_366),
.B(n_367),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_SL g467 ( 
.A1(n_448),
.A2(n_351),
.B(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_332),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_411),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_376),
.C(n_341),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_337),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

BUFx4f_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

BUFx4f_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_397),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_343),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_399),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_407),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_306),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_435),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_310),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_314),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_362),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_438),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_372),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_410),
.B(n_340),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_314),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_439),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_448),
.B(n_335),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_400),
.A2(n_395),
.B1(n_394),
.B2(n_391),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_328),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_434),
.B(n_328),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_434),
.B(n_329),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_381),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_450),
.B(n_329),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_410),
.B(n_312),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_428),
.A2(n_380),
.B1(n_363),
.B2(n_378),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_440),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_398),
.B(n_353),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_432),
.B(n_353),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_429),
.B(n_364),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_400),
.A2(n_383),
.B1(n_318),
.B2(n_346),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_431),
.B(n_244),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_450),
.B(n_460),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_407),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_330),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_483),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_497),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_490),
.B(n_451),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_492),
.B(n_396),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_467),
.A2(n_418),
.B(n_417),
.C(n_398),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_468),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_417),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_474),
.B(n_396),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_483),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_485),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_483),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_484),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g552 ( 
.A(n_529),
.B(n_451),
.C(n_438),
.Y(n_552)
);

AND2x6_ASAP7_75t_SL g553 ( 
.A(n_494),
.B(n_441),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_418),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_459),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_469),
.B(n_396),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_459),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_467),
.A2(n_443),
.B1(n_431),
.B2(n_454),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_497),
.B(n_432),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_473),
.B(n_432),
.C(n_441),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_484),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_404),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_497),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_497),
.B(n_491),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_491),
.B(n_459),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_404),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_480),
.B(n_501),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_475),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_475),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_498),
.B(n_459),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_498),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_L g584 ( 
.A1(n_493),
.A2(n_461),
.B1(n_403),
.B2(n_373),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_500),
.B(n_504),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_515),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_503),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_L g588 ( 
.A(n_502),
.B(n_509),
.C(n_508),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_459),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_504),
.B(n_459),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_506),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_517),
.B(n_459),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_396),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_402),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_503),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_512),
.B(n_431),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_518),
.B(n_402),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_499),
.B(n_402),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_507),
.B(n_402),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_520),
.B(n_431),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_506),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_520),
.B(n_443),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_536),
.B(n_461),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_512),
.B(n_330),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_525),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_524),
.B(n_443),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_479),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_525),
.B(n_414),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_525),
.B(n_461),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_L g614 ( 
.A(n_496),
.B(n_348),
.C(n_331),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_510),
.B(n_331),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_533),
.B(n_443),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_533),
.B(n_454),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_481),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_513),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_516),
.B(n_360),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_454),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_476),
.A2(n_414),
.B(n_387),
.C(n_454),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_526),
.B(n_506),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_526),
.B(n_416),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_530),
.B(n_522),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_522),
.B(n_356),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_522),
.B(n_360),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_530),
.B(n_375),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_521),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_416),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_526),
.B(n_416),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_476),
.B(n_414),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_576),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_608),
.A2(n_477),
.B1(n_476),
.B2(n_308),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

BUFx4f_ASAP7_75t_L g638 ( 
.A(n_540),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_624),
.A2(n_477),
.B(n_476),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_545),
.A2(n_477),
.B(n_489),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_608),
.B(n_477),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_543),
.B(n_526),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_611),
.A2(n_535),
.B(n_527),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_554),
.A2(n_470),
.B(n_531),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_611),
.A2(n_527),
.B(n_515),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_625),
.A2(n_470),
.B(n_531),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_576),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_632),
.A2(n_470),
.B(n_531),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_558),
.A2(n_530),
.B1(n_495),
.B2(n_403),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_633),
.A2(n_470),
.B(n_531),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_575),
.B(n_526),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_540),
.B(n_628),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_561),
.A2(n_521),
.B(n_530),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_583),
.B(n_526),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_562),
.A2(n_528),
.B(n_471),
.Y(n_656)
);

INVx11_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_613),
.A2(n_436),
.B(n_465),
.C(n_514),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g660 ( 
.A1(n_626),
.A2(n_528),
.B(n_514),
.C(n_478),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_583),
.B(n_466),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_576),
.B(n_403),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g663 ( 
.A1(n_557),
.A2(n_412),
.B(n_409),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_561),
.A2(n_521),
.B(n_471),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_560),
.B(n_462),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_562),
.A2(n_471),
.B(n_466),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_466),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_558),
.A2(n_307),
.B(n_368),
.C(n_374),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_615),
.A2(n_316),
.B1(n_339),
.B2(n_373),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_R g670 ( 
.A(n_553),
.B(n_368),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_623),
.A2(n_634),
.B(n_538),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_596),
.B(n_466),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_588),
.A2(n_374),
.B1(n_379),
.B2(n_478),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_634),
.A2(n_521),
.B(n_478),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_577),
.B(n_602),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_550),
.B(n_379),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_537),
.Y(n_677)
);

OAI21xp33_ASAP7_75t_L g678 ( 
.A1(n_574),
.A2(n_294),
.B(n_293),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_577),
.Y(n_679)
);

INVx11_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_559),
.B(n_189),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_577),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_539),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_574),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_568),
.A2(n_521),
.B(n_478),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_630),
.A2(n_505),
.B(n_471),
.Y(n_686)
);

NOR3xp33_ASAP7_75t_L g687 ( 
.A(n_605),
.B(n_465),
.C(n_436),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_577),
.Y(n_688)
);

O2A1O1Ixp5_ASAP7_75t_L g689 ( 
.A1(n_585),
.A2(n_505),
.B(n_419),
.C(n_416),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_555),
.A2(n_521),
.B(n_505),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_577),
.B(n_190),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_601),
.A2(n_505),
.B(n_472),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_606),
.B(n_462),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_541),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_596),
.B(n_449),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_560),
.A2(n_298),
.B1(n_192),
.B2(n_197),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_602),
.B(n_246),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_591),
.A2(n_190),
.B1(n_295),
.B2(n_192),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_607),
.B(n_449),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_603),
.A2(n_412),
.B(n_409),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_616),
.A2(n_472),
.B(n_413),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_607),
.B(n_453),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_544),
.B(n_419),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_604),
.A2(n_250),
.B1(n_252),
.B2(n_257),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_548),
.B(n_419),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_537),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_552),
.B(n_464),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_548),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_609),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_565),
.B(n_419),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_586),
.A2(n_472),
.B(n_413),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_572),
.A2(n_589),
.B(n_581),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_453),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_609),
.A2(n_602),
.B1(n_591),
.B2(n_622),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_627),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_617),
.A2(n_597),
.B(n_593),
.C(n_594),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_590),
.A2(n_472),
.B(n_413),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_566),
.A2(n_412),
.B(n_409),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_592),
.A2(n_472),
.B(n_413),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_566),
.B(n_453),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_602),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_630),
.A2(n_472),
.B(n_407),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_547),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_564),
.B(n_553),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_630),
.A2(n_407),
.B(n_421),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_629),
.B(n_464),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_557),
.A2(n_422),
.B(n_421),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_570),
.B(n_453),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_546),
.A2(n_457),
.B(n_455),
.C(n_452),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_570),
.A2(n_422),
.B(n_421),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_578),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_578),
.B(n_422),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_582),
.A2(n_426),
.B(n_425),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_706),
.B(n_717),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_654),
.A2(n_651),
.B(n_639),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_683),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_638),
.B(n_602),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_641),
.A2(n_556),
.B1(n_542),
.B2(n_599),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_SL g741 ( 
.A(n_670),
.B(n_614),
.C(n_673),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_693),
.B(n_629),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_684),
.A2(n_600),
.B1(n_621),
.B2(n_584),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_647),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_638),
.B(n_567),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_641),
.A2(n_582),
.B1(n_631),
.B2(n_618),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_652),
.B(n_631),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_640),
.A2(n_549),
.B(n_547),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_677),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_598),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_728),
.B(n_598),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_636),
.A2(n_620),
.B1(n_618),
.B2(n_612),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_647),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_653),
.Y(n_754)
);

CKINVDCx14_ASAP7_75t_R g755 ( 
.A(n_669),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_676),
.B(n_452),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_SL g757 ( 
.A(n_718),
.B(n_681),
.C(n_668),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_694),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_662),
.B(n_610),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_655),
.A2(n_551),
.B(n_549),
.Y(n_760)
);

AO21x1_ASAP7_75t_L g761 ( 
.A1(n_642),
.A2(n_612),
.B(n_610),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_655),
.B(n_567),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_695),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_726),
.B(n_455),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_649),
.B(n_197),
.Y(n_765)
);

BUFx2_ASAP7_75t_SL g766 ( 
.A(n_647),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_708),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_725),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_696),
.B(n_620),
.Y(n_769)
);

AOI21x1_ASAP7_75t_L g770 ( 
.A1(n_642),
.A2(n_563),
.B(n_551),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_709),
.B(n_457),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_710),
.B(n_563),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_733),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_644),
.A2(n_571),
.B(n_569),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_716),
.B(n_595),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_665),
.B(n_569),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_665),
.B(n_458),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_734),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_734),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_671),
.B(n_571),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_635),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_700),
.B(n_573),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_657),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_678),
.B(n_458),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_658),
.B(n_573),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_697),
.B(n_423),
.C(n_425),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_579),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_635),
.B(n_579),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_674),
.A2(n_595),
.B(n_587),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_664),
.A2(n_587),
.B(n_580),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_667),
.B(n_580),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_646),
.A2(n_426),
.B(n_259),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_648),
.A2(n_426),
.B(n_261),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_682),
.B(n_408),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_637),
.B(n_423),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_686),
.A2(n_427),
.B(n_447),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_680),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_SL g798 ( 
.A1(n_714),
.A2(n_427),
.B(n_447),
.C(n_445),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_682),
.B(n_258),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_637),
.B(n_408),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_659),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_659),
.B(n_269),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_679),
.B(n_415),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_650),
.A2(n_273),
.B(n_276),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_731),
.A2(n_415),
.B(n_447),
.C(n_445),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_679),
.B(n_437),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_748),
.A2(n_663),
.B(n_656),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_757),
.A2(n_643),
.B(n_691),
.C(n_660),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_761),
.A2(n_729),
.A3(n_685),
.B(n_735),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_776),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_796),
.A2(n_666),
.B(n_690),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_774),
.A2(n_645),
.B(n_689),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_742),
.A2(n_661),
.B1(n_730),
.B2(n_715),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_737),
.A2(n_732),
.A3(n_661),
.B(n_704),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_781),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_738),
.B(n_741),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_753),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_765),
.A2(n_705),
.B(n_699),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_785),
.A2(n_675),
.B(n_701),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_764),
.B(n_711),
.C(n_698),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_780),
.A2(n_720),
.B(n_692),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_758),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_738),
.B(n_688),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_789),
.A2(n_719),
.B(n_721),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_736),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_790),
.A2(n_702),
.B(n_727),
.Y(n_827)
);

AO31x2_ASAP7_75t_L g828 ( 
.A1(n_740),
.A2(n_730),
.A3(n_704),
.B(n_707),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_780),
.A2(n_703),
.B(n_722),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_757),
.A2(n_722),
.B(n_715),
.C(n_707),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_762),
.A2(n_712),
.B(n_723),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_756),
.B(n_688),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_743),
.A2(n_712),
.B(n_723),
.C(n_437),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_783),
.B(n_797),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_763),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_777),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_743),
.A2(n_437),
.B(n_456),
.C(n_445),
.Y(n_837)
);

OAI22x1_ASAP7_75t_L g838 ( 
.A1(n_771),
.A2(n_773),
.B1(n_745),
.B2(n_739),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_741),
.A2(n_713),
.B(n_724),
.C(n_295),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_762),
.A2(n_456),
.B(n_444),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_755),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_SL g842 ( 
.A1(n_802),
.A2(n_456),
.B(n_444),
.C(n_122),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_444),
.B(n_303),
.C(n_302),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_751),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_781),
.Y(n_845)
);

AO31x2_ASAP7_75t_L g846 ( 
.A1(n_746),
.A2(n_793),
.A3(n_792),
.B(n_750),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_769),
.B(n_747),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_778),
.B(n_199),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_SL g849 ( 
.A1(n_802),
.A2(n_113),
.B(n_183),
.C(n_181),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_781),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_749),
.Y(n_851)
);

OA22x2_ASAP7_75t_L g852 ( 
.A1(n_759),
.A2(n_297),
.B1(n_294),
.B2(n_293),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_760),
.A2(n_279),
.B(n_298),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_801),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_770),
.A2(n_109),
.B(n_180),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_779),
.B(n_776),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_787),
.A2(n_430),
.B(n_296),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_806),
.A2(n_107),
.B(n_179),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_767),
.Y(n_859)
);

OAI22x1_ASAP7_75t_L g860 ( 
.A1(n_745),
.A2(n_297),
.B1(n_201),
.B2(n_202),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_775),
.A2(n_430),
.B(n_296),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_753),
.B(n_781),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_768),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_791),
.A2(n_430),
.B(n_292),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_798),
.A2(n_788),
.B(n_799),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_819),
.A2(n_786),
.B1(n_784),
.B2(n_759),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_847),
.B(n_801),
.Y(n_867)
);

INVx6_ASAP7_75t_L g868 ( 
.A(n_810),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_862),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_815),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_819),
.A2(n_759),
.B1(n_799),
.B2(n_803),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_815),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_828),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_817),
.A2(n_803),
.B1(n_800),
.B2(n_794),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_820),
.A2(n_798),
.B(n_788),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_852),
.A2(n_797),
.B1(n_783),
.B2(n_766),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_SL g878 ( 
.A1(n_821),
.A2(n_794),
.B1(n_753),
.B2(n_800),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_SL g879 ( 
.A1(n_821),
.A2(n_753),
.B1(n_772),
.B2(n_202),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_828),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

CKINVDCx6p67_ASAP7_75t_R g882 ( 
.A(n_834),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_809),
.Y(n_883)
);

CKINVDCx14_ASAP7_75t_R g884 ( 
.A(n_841),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_828),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_844),
.B(n_795),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_836),
.A2(n_782),
.B1(n_804),
.B2(n_752),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_823),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_835),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_818),
.Y(n_890)
);

OAI22xp33_ASAP7_75t_L g891 ( 
.A1(n_848),
.A2(n_199),
.B1(n_201),
.B2(n_206),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_837),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_816),
.B(n_744),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_838),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_851),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_854),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_818),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_859),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_860),
.A2(n_752),
.B1(n_744),
.B2(n_292),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_853),
.A2(n_279),
.B1(n_210),
.B2(n_206),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_SL g902 ( 
.A1(n_853),
.A2(n_210),
.B1(n_9),
.B2(n_10),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_856),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_863),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_832),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_809),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_855),
.Y(n_907)
);

OAI22x1_ASAP7_75t_L g908 ( 
.A1(n_824),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_816),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_818),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_845),
.Y(n_911)
);

INVx3_ASAP7_75t_SL g912 ( 
.A(n_834),
.Y(n_912)
);

CKINVDCx11_ASAP7_75t_R g913 ( 
.A(n_814),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_833),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_814),
.A2(n_861),
.B1(n_865),
.B2(n_831),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_809),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_807),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_845),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_850),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_850),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_812),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_849),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_857),
.A2(n_805),
.B1(n_11),
.B2(n_12),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_864),
.A2(n_840),
.B1(n_829),
.B2(n_822),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_858),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_916),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_875),
.A2(n_825),
.B(n_827),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_916),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_925),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_894),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_883),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_873),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_873),
.Y(n_933)
);

CKINVDCx14_ASAP7_75t_R g934 ( 
.A(n_884),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_873),
.A2(n_811),
.B(n_843),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_880),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_880),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_917),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_897),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_925),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_918),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_880),
.A2(n_846),
.B(n_808),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_902),
.A2(n_7),
.B1(n_11),
.B2(n_14),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_894),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_917),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_885),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_870),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_885),
.B(n_846),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_882),
.B(n_839),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_870),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_872),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_885),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_883),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_872),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_925),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_872),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_883),
.B(n_846),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_921),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_921),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_883),
.B(n_830),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_906),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_906),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_930),
.B(n_881),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_943),
.A2(n_866),
.B(n_879),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_958),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_930),
.B(n_881),
.Y(n_966)
);

OR2x2_ASAP7_75t_SL g967 ( 
.A(n_934),
.B(n_868),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_943),
.A2(n_915),
.B(n_923),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_930),
.B(n_881),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_930),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_944),
.B(n_929),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_959),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_944),
.B(n_905),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_944),
.B(n_867),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_944),
.B(n_906),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_927),
.A2(n_924),
.B(n_907),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_960),
.B(n_867),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_949),
.A2(n_891),
.B(n_900),
.C(n_901),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_945),
.B(n_906),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_945),
.B(n_876),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_929),
.B(n_876),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_938),
.B(n_888),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_934),
.A2(n_877),
.B1(n_903),
.B2(n_874),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_938),
.B(n_888),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_958),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_960),
.B(n_889),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_949),
.B(n_913),
.C(n_871),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_939),
.A2(n_908),
.B1(n_903),
.B2(n_878),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_955),
.A2(n_886),
.B(n_889),
.C(n_919),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_960),
.B(n_909),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_929),
.B(n_909),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_926),
.A2(n_904),
.B(n_895),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_939),
.B(n_912),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_938),
.B(n_895),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_941),
.B(n_911),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_929),
.B(n_907),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_941),
.B(n_911),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_942),
.A2(n_914),
.B(n_892),
.C(n_887),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_927),
.A2(n_914),
.B(n_892),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_955),
.A2(n_899),
.B(n_904),
.C(n_908),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_948),
.B(n_899),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_948),
.A2(n_922),
.B1(n_882),
.B2(n_912),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_929),
.B(n_920),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_955),
.A2(n_842),
.B(n_912),
.C(n_869),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_958),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_1001),
.B(n_957),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_971),
.B(n_948),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_965),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_986),
.B(n_926),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_996),
.B(n_929),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_972),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_971),
.B(n_929),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_982),
.B(n_957),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_985),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_986),
.B(n_926),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_981),
.B(n_929),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_981),
.B(n_929),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_964),
.A2(n_922),
.B1(n_896),
.B2(n_868),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_977),
.B(n_940),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1005),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_996),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_974),
.B(n_940),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_990),
.B(n_940),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_988),
.A2(n_922),
.B1(n_957),
.B2(n_896),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_984),
.B(n_942),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_964),
.A2(n_940),
.B1(n_868),
.B2(n_896),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_999),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_994),
.B(n_942),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_992),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_980),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_996),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_973),
.B(n_928),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1019),
.B(n_970),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1029),
.A2(n_989),
.B(n_968),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1019),
.B(n_991),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1020),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1010),
.B(n_991),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_1024),
.A2(n_968),
.B1(n_987),
.B2(n_983),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1020),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1025),
.B(n_979),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1010),
.B(n_1003),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1008),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_1021),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1011),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1010),
.B(n_1003),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1011),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1010),
.B(n_940),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1029),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1031),
.B(n_940),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1008),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1031),
.B(n_940),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1031),
.B(n_940),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1025),
.B(n_975),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_1014),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1055),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1048),
.B(n_1021),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1043),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.B(n_1012),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1034),
.B(n_1030),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1043),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1045),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1051),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1048),
.B(n_1044),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1035),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1044),
.B(n_1012),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_1065),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1059),
.Y(n_1069)
);

AND2x4_ASAP7_75t_SL g1070 ( 
.A(n_1065),
.B(n_1018),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1066),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1059),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1062),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1066),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1062),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1070),
.B(n_1061),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1069),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1072),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_1073),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_1060),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1077),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1076),
.A2(n_1039),
.B1(n_1070),
.B2(n_1024),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1078),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_1081),
.B(n_1034),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1081),
.A2(n_1018),
.B1(n_987),
.B2(n_983),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1080),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1079),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1079),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1077),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1076),
.B(n_1060),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_1076),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1077),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1088),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1092),
.B(n_1049),
.Y(n_1095)
);

OAI322xp33_ASAP7_75t_L g1096 ( 
.A1(n_1089),
.A2(n_1049),
.A3(n_1057),
.B1(n_1056),
.B2(n_1074),
.C1(n_1071),
.C2(n_988),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_1082),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1084),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1085),
.Y(n_1099)
);

OAI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_1083),
.A2(n_1086),
.B1(n_1085),
.B2(n_1091),
.C(n_1087),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1090),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_978),
.B(n_1026),
.Y(n_1102)
);

AOI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1092),
.A2(n_1063),
.B1(n_1056),
.B2(n_1057),
.C1(n_1058),
.C2(n_1074),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1088),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1086),
.A2(n_1071),
.B(n_993),
.Y(n_1105)
);

OAI321xp33_ASAP7_75t_L g1106 ( 
.A1(n_1092),
.A2(n_1002),
.A3(n_1058),
.B1(n_1067),
.B2(n_1064),
.C(n_1004),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1088),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1092),
.B(n_1067),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1092),
.B(n_1064),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1092),
.B(n_1000),
.C(n_998),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1097),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1097),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1094),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1104),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1107),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1099),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1099),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1108),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1109),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1100),
.B(n_967),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1110),
.A2(n_997),
.B(n_995),
.C(n_1002),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1095),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1103),
.A2(n_1052),
.B(n_1050),
.Y(n_1124)
);

AOI33xp33_ASAP7_75t_L g1125 ( 
.A1(n_1098),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.B3(n_18),
.Y(n_1125)
);

OAI211xp5_ASAP7_75t_L g1126 ( 
.A1(n_1101),
.A2(n_1053),
.B(n_1052),
.C(n_1050),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1096),
.A2(n_1066),
.B1(n_1030),
.B2(n_1051),
.C(n_1052),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1102),
.B(n_1033),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1106),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1094),
.B(n_1033),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1122),
.B(n_1036),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1120),
.A2(n_1053),
.B1(n_1050),
.B2(n_1038),
.Y(n_1132)
);

BUFx8_ASAP7_75t_SL g1133 ( 
.A(n_1117),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1111),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1116),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1112),
.B(n_1032),
.C(n_898),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1118),
.B(n_1036),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1129),
.B(n_1047),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1123),
.B(n_1035),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1130),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1113),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1114),
.B(n_1035),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1121),
.A2(n_1053),
.B(n_1038),
.C(n_1046),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_1120),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1125),
.B(n_1033),
.Y(n_1145)
);

AND2x4_ASAP7_75t_SL g1146 ( 
.A(n_1115),
.B(n_1038),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1119),
.B(n_1121),
.C(n_1128),
.D(n_1127),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1124),
.A2(n_940),
.B1(n_1038),
.B2(n_969),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1134),
.B(n_1125),
.C(n_1144),
.Y(n_1149)
);

NOR4xp25_ASAP7_75t_L g1150 ( 
.A(n_1135),
.B(n_1126),
.C(n_16),
.D(n_17),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1147),
.A2(n_1037),
.B1(n_1032),
.B2(n_1040),
.C(n_1042),
.Y(n_1151)
);

OAI211xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1138),
.A2(n_1054),
.B(n_1041),
.C(n_19),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1141),
.B(n_898),
.C(n_890),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1145),
.A2(n_1137),
.B1(n_1146),
.B2(n_1132),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1140),
.A2(n_1046),
.B(n_1042),
.Y(n_1155)
);

AOI211x1_ASAP7_75t_SL g1156 ( 
.A1(n_1136),
.A2(n_1139),
.B(n_1142),
.C(n_1143),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1142),
.A2(n_15),
.B(n_18),
.Y(n_1157)
);

AOI222xp33_ASAP7_75t_L g1158 ( 
.A1(n_1139),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.C1(n_26),
.C2(n_27),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1131),
.B(n_1148),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1133),
.A2(n_1027),
.B1(n_969),
.B2(n_955),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1144),
.A2(n_1054),
.B1(n_1041),
.B2(n_1040),
.Y(n_1161)
);

OAI211xp5_ASAP7_75t_L g1162 ( 
.A1(n_1147),
.A2(n_890),
.B(n_898),
.C(n_910),
.Y(n_1162)
);

NAND5xp2_ASAP7_75t_L g1163 ( 
.A(n_1144),
.B(n_1046),
.C(n_1042),
.D(n_966),
.E(n_1017),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1135),
.B(n_1040),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1134),
.Y(n_1165)
);

XNOR2xp5_ASAP7_75t_L g1166 ( 
.A(n_1147),
.B(n_22),
.Y(n_1166)
);

OAI211xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1144),
.A2(n_23),
.B(n_26),
.C(n_28),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1135),
.A2(n_1037),
.B(n_963),
.C(n_32),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1135),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1135),
.B(n_890),
.C(n_910),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_L g1171 ( 
.A(n_1144),
.B(n_910),
.C(n_1009),
.Y(n_1171)
);

OAI211xp5_ASAP7_75t_L g1172 ( 
.A1(n_1147),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1165),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1149),
.A2(n_1027),
.B(n_869),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1157),
.Y(n_1175)
);

OAI211xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1156),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_1176)
);

OAI221xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1172),
.A2(n_1016),
.B1(n_1017),
.B2(n_1022),
.C(n_1028),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1169),
.Y(n_1178)
);

AOI21xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1150),
.A2(n_33),
.B(n_34),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1167),
.A2(n_1158),
.B(n_1152),
.C(n_1168),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_1166),
.A2(n_1027),
.B1(n_1014),
.B2(n_1015),
.C(n_1009),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1154),
.B(n_36),
.Y(n_1182)
);

OAI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1158),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1151),
.A2(n_1015),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1184)
);

OAI221xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1162),
.A2(n_1016),
.B1(n_1022),
.B2(n_1028),
.C(n_1023),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1159),
.Y(n_1186)
);

OAI31xp33_ASAP7_75t_L g1187 ( 
.A1(n_1153),
.A2(n_869),
.A3(n_1023),
.B(n_45),
.Y(n_1187)
);

AOI21xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1170),
.A2(n_37),
.B(n_40),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1164),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1171),
.A2(n_47),
.B1(n_48),
.B2(n_920),
.C(n_893),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1155),
.A2(n_47),
.B(n_976),
.C(n_942),
.Y(n_1191)
);

AOI221xp5_ASAP7_75t_L g1192 ( 
.A1(n_1160),
.A2(n_893),
.B1(n_1007),
.B2(n_928),
.C(n_1006),
.Y(n_1192)
);

OAI211xp5_ASAP7_75t_L g1193 ( 
.A1(n_1161),
.A2(n_51),
.B(n_56),
.C(n_57),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1163),
.A2(n_893),
.B(n_935),
.Y(n_1194)
);

OAI31xp33_ASAP7_75t_L g1195 ( 
.A1(n_1172),
.A2(n_893),
.A3(n_1007),
.B(n_1006),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1150),
.A2(n_928),
.B1(n_1013),
.B2(n_959),
.C(n_961),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1186),
.B(n_1013),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1175),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1178),
.B(n_65),
.Y(n_1199)
);

XOR2x1_ASAP7_75t_L g1200 ( 
.A(n_1173),
.B(n_66),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_L g1201 ( 
.A(n_1188),
.B(n_68),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1189),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1182),
.B(n_959),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1179),
.B(n_70),
.Y(n_1204)
);

XNOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_1183),
.B(n_76),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1180),
.Y(n_1206)
);

XNOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1190),
.B(n_78),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1184),
.B(n_81),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1176),
.A2(n_868),
.B1(n_896),
.B2(n_959),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1194),
.Y(n_1210)
);

NAND4xp75_ASAP7_75t_L g1211 ( 
.A(n_1187),
.B(n_84),
.C(n_86),
.D(n_93),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1195),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1177),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1196),
.B(n_1181),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1193),
.B(n_962),
.C(n_961),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1193),
.A2(n_868),
.B1(n_896),
.B2(n_962),
.Y(n_1216)
);

XNOR2xp5_ASAP7_75t_L g1217 ( 
.A(n_1174),
.B(n_98),
.Y(n_1217)
);

NOR2x1_ASAP7_75t_L g1218 ( 
.A(n_1191),
.B(n_1185),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1206),
.B(n_1192),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_L g1220 ( 
.A(n_1202),
.B(n_99),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1201),
.B(n_102),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1204),
.B(n_110),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1198),
.A2(n_962),
.B1(n_961),
.B2(n_946),
.C(n_952),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1198),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_L g1225 ( 
.A(n_1199),
.B(n_111),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1200),
.B(n_119),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1197),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1205),
.B(n_123),
.Y(n_1228)
);

XNOR2x1_ASAP7_75t_SL g1229 ( 
.A(n_1208),
.B(n_126),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1213),
.B(n_1212),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1209),
.A2(n_953),
.B1(n_937),
.B2(n_932),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1216),
.B(n_935),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1214),
.A2(n_932),
.B1(n_946),
.B2(n_936),
.C(n_952),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1225),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1222),
.Y(n_1235)
);

AOI221xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1230),
.A2(n_1224),
.B1(n_1210),
.B2(n_1219),
.C(n_1227),
.Y(n_1236)
);

XNOR2x1_ASAP7_75t_L g1237 ( 
.A(n_1229),
.B(n_1207),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1221),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1228),
.A2(n_1218),
.B1(n_1211),
.B2(n_1217),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1220),
.B(n_1215),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1226),
.B(n_1203),
.Y(n_1241)
);

XNOR2x1_ASAP7_75t_L g1242 ( 
.A(n_1231),
.B(n_1203),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1232),
.B(n_127),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1233),
.B(n_130),
.Y(n_1244)
);

NAND3x1_ASAP7_75t_L g1245 ( 
.A(n_1223),
.B(n_131),
.C(n_132),
.Y(n_1245)
);

AOI211x1_ASAP7_75t_L g1246 ( 
.A1(n_1230),
.A2(n_952),
.B(n_946),
.C(n_937),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1230),
.A2(n_932),
.B1(n_933),
.B2(n_936),
.C(n_937),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1220),
.B(n_135),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1248),
.Y(n_1249)
);

AO22x2_ASAP7_75t_L g1250 ( 
.A1(n_1237),
.A2(n_1239),
.B1(n_1235),
.B2(n_1238),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1236),
.A2(n_1240),
.B1(n_1234),
.B2(n_1241),
.Y(n_1251)
);

AO22x2_ASAP7_75t_L g1252 ( 
.A1(n_1242),
.A2(n_933),
.B1(n_936),
.B2(n_954),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1243),
.A2(n_933),
.B1(n_138),
.B2(n_141),
.C(n_142),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1244),
.A2(n_953),
.B1(n_935),
.B2(n_931),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_1246),
.A2(n_954),
.B1(n_931),
.B2(n_951),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1245),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1247),
.A2(n_953),
.B1(n_935),
.B2(n_931),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1237),
.A2(n_954),
.B1(n_931),
.B2(n_951),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1250),
.A2(n_931),
.B1(n_951),
.B2(n_950),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1256),
.A2(n_137),
.B1(n_144),
.B2(n_145),
.C(n_151),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1249),
.A2(n_931),
.B1(n_951),
.B2(n_950),
.Y(n_1261)
);

XNOR2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1251),
.B(n_1254),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1253),
.A2(n_956),
.B1(n_950),
.B2(n_947),
.Y(n_1263)
);

XOR2x2_ASAP7_75t_L g1264 ( 
.A(n_1257),
.B(n_156),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1264),
.Y(n_1265)
);

XNOR2x1_ASAP7_75t_L g1266 ( 
.A(n_1262),
.B(n_1258),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1260),
.A2(n_1252),
.B1(n_1255),
.B2(n_956),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1259),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1268),
.A2(n_1263),
.B1(n_1261),
.B2(n_956),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_1266),
.B(n_1265),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1270),
.B(n_1267),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_927),
.B(n_159),
.Y(n_1272)
);

AOI221xp5_ASAP7_75t_L g1273 ( 
.A1(n_1272),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.C(n_163),
.Y(n_1273)
);

AOI211xp5_ASAP7_75t_L g1274 ( 
.A1(n_1273),
.A2(n_165),
.B(n_168),
.C(n_169),
.Y(n_1274)
);


endmodule