module fake_aes_7141_n_1078 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_1078);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_1078;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_560;
wire n_517;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_230;
wire n_209;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_235;
wire n_482;
wire n_243;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_788;
wire n_1035;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_937;
wire n_217;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_695;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g209 ( .A(n_114), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_30), .Y(n_210) );
NOR2xp67_ASAP7_75t_L g211 ( .A(n_179), .B(n_132), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_84), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_202), .Y(n_213) );
INVx4_ASAP7_75t_R g214 ( .A(n_86), .Y(n_214) );
INVxp33_ASAP7_75t_SL g215 ( .A(n_163), .Y(n_215) );
CKINVDCx14_ASAP7_75t_R g216 ( .A(n_47), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_204), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_43), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_89), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_181), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_156), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_17), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_28), .B(n_13), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_144), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_27), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_51), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_198), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_47), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_20), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_147), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_141), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_96), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_27), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_46), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_17), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_95), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_56), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_58), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_60), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_52), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_97), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_94), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_172), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_120), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_177), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_79), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_16), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_62), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_46), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_136), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_29), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_158), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_149), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_29), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_189), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_123), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_45), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_152), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_155), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_137), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_206), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_199), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_32), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_145), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_99), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_151), .Y(n_269) );
CKINVDCx16_ASAP7_75t_R g270 ( .A(n_57), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_13), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_153), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_115), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g275 ( .A(n_0), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_164), .Y(n_276) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_148), .Y(n_277) );
BUFx2_ASAP7_75t_SL g278 ( .A(n_10), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_201), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_107), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_105), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_19), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_23), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_142), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_169), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_150), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_166), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_167), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_18), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_135), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_100), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_208), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_55), .Y(n_293) );
CKINVDCx16_ASAP7_75t_R g294 ( .A(n_121), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_38), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_207), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_28), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_22), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_108), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_146), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_11), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_51), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_35), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_143), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_134), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_76), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_165), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_70), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_71), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_191), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_69), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_203), .Y(n_313) );
CKINVDCx16_ASAP7_75t_R g314 ( .A(n_194), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_101), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_66), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_117), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_109), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_39), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_124), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_43), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_154), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_185), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_192), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_106), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_171), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_40), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_129), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_219), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_217), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_248), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_217), .B(n_1), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_217), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_219), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_216), .B(n_1), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_219), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_322), .B(n_2), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_219), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_232), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_232), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_275), .B(n_2), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_232), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_234), .B(n_85), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_232), .Y(n_345) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_221), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_306), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_240), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_275), .B(n_263), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_271), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
INVx5_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_322), .B(n_3), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_223), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_246), .B(n_4), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_271), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_230), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_258), .B(n_6), .Y(n_359) );
INVx6_ASAP7_75t_L g360 ( .A(n_288), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_274), .B(n_7), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_289), .B(n_8), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_210), .B(n_8), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_236), .B(n_9), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_349), .B(n_277), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_349), .B(n_279), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_349), .B(n_294), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_330), .B(n_331), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
NAND2xp33_ASAP7_75t_R g373 ( .A(n_344), .B(n_215), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_364), .B(n_314), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_330), .B(n_218), .Y(n_376) );
INVx6_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_332), .B(n_221), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_329), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_332), .B(n_253), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_346), .B(n_247), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_228), .B1(n_239), .B2(n_235), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_332), .B(n_248), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
INVx4_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_330), .B(n_222), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_329), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_338), .B(n_289), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
INVx4_ASAP7_75t_L g392 ( .A(n_344), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_331), .B(n_218), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_331), .Y(n_394) );
AND2x6_ASAP7_75t_L g395 ( .A(n_338), .B(n_288), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_338), .B(n_310), .Y(n_396) );
INVx5_ASAP7_75t_L g397 ( .A(n_360), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
INVx4_ASAP7_75t_SL g399 ( .A(n_344), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_336), .B(n_226), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_363), .B(n_212), .C(n_209), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_364), .A2(n_241), .B1(n_249), .B2(n_242), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_336), .A2(n_270), .B1(n_321), .B2(n_231), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_338), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_342), .Y(n_407) );
NOR2x1p5_ASAP7_75t_L g408 ( .A(n_346), .B(n_226), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_364), .B(n_327), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_342), .B(n_237), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_377), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_385), .B(n_354), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_376), .B(n_346), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_366), .B(n_359), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_385), .B(n_354), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_407), .B(n_354), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
NOR2x1p5_ASAP7_75t_L g418 ( .A(n_409), .B(n_359), .Y(n_418) );
INVx5_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_383), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_407), .B(n_354), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_390), .Y(n_423) );
NOR2x1p5_ASAP7_75t_L g424 ( .A(n_409), .B(n_361), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_368), .B(n_393), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_385), .B(n_213), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_385), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_405), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_392), .B(n_220), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_392), .B(n_229), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_400), .B(n_344), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_378), .B(n_356), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_410), .B(n_344), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_380), .B(n_363), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_392), .A2(n_348), .B1(n_351), .B2(n_334), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_348), .B1(n_351), .B2(n_334), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_371), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_384), .A2(n_357), .B1(n_252), .B2(n_257), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_403), .B(n_237), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_369), .B(n_215), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_377), .Y(n_446) );
AND2x6_ASAP7_75t_SL g447 ( .A(n_381), .B(n_250), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_399), .B(n_233), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_403), .B(n_254), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_382), .B(n_255), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_395), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_373), .A2(n_358), .B1(n_355), .B2(n_225), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_396), .B(n_256), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_395), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_395), .B(n_256), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_395), .B(n_259), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_406), .A2(n_358), .B(n_355), .C(n_282), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_367), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_399), .B(n_238), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_399), .B(n_245), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_395), .B(n_259), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_383), .B(n_269), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_367), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_406), .A2(n_227), .B(n_222), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_371), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_391), .B(n_269), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_388), .A2(n_283), .B1(n_293), .B2(n_266), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_388), .B(n_311), .Y(n_470) );
NAND2x1_ASAP7_75t_L g471 ( .A(n_388), .B(n_214), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_388), .B(n_286), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_372), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_404), .B(n_401), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_402), .B(n_254), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_372), .Y(n_476) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_408), .B(n_224), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_375), .A2(n_299), .B1(n_304), .B2(n_302), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_387), .B(n_308), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_394), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_394), .Y(n_481) );
NAND3xp33_ASAP7_75t_SL g482 ( .A(n_370), .B(n_305), .C(n_301), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_398), .B(n_313), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_397), .B(n_323), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_397), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_397), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_397), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_397), .A2(n_295), .B1(n_303), .B2(n_298), .Y(n_488) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_365), .B(n_316), .C(n_303), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_414), .B(n_309), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_418), .B(n_307), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_412), .A2(n_261), .B(n_365), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_SL g493 ( .A1(n_413), .A2(n_337), .B(n_339), .C(n_335), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_424), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_459), .A2(n_312), .B(n_310), .C(n_251), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_452), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_477), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_482), .B(n_278), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_426), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_419), .B(n_243), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_417), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_415), .A2(n_389), .B(n_386), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_428), .A2(n_264), .B(n_262), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_445), .B(n_244), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_428), .A2(n_273), .B(n_272), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_432), .A2(n_280), .B(n_276), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_432), .A2(n_285), .B(n_284), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_444), .B(n_260), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_420), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_438), .A2(n_291), .B(n_292), .C(n_287), .Y(n_510) );
INVx3_ASAP7_75t_SL g511 ( .A(n_475), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_433), .A2(n_300), .B(n_296), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_442), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_423), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_441), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_433), .A2(n_325), .B(n_317), .Y(n_516) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_434), .A2(n_328), .B(n_326), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_429), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_474), .A2(n_281), .B(n_267), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_436), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_451), .A2(n_281), .B(n_320), .C(n_290), .Y(n_522) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_477), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_429), .B(n_265), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_479), .B(n_360), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_438), .A2(n_360), .B1(n_260), .B2(n_319), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_429), .B(n_464), .Y(n_527) );
OR2x6_ASAP7_75t_L g528 ( .A(n_429), .B(n_260), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_471), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_445), .B(n_268), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_455), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_437), .A2(n_320), .B1(n_290), .B2(n_319), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_416), .A2(n_297), .B(n_324), .C(n_318), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_422), .A2(n_297), .B(n_324), .C(n_318), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_449), .B(n_453), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_441), .Y(n_536) );
OR2x6_ASAP7_75t_L g537 ( .A(n_442), .B(n_260), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_435), .B(n_211), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_489), .B(n_319), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_454), .A2(n_335), .B(n_339), .C(n_337), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_442), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_469), .B(n_319), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_460), .A2(n_353), .B(n_341), .Y(n_543) );
BUFx12f_ASAP7_75t_L g544 ( .A(n_447), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_470), .A2(n_340), .B1(n_347), .B2(n_343), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_469), .B(n_9), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_465), .A2(n_353), .B(n_343), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_439), .A2(n_440), .B1(n_443), .B2(n_468), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_467), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_467), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_466), .A2(n_340), .B(n_352), .C(n_347), .Y(n_552) );
BUFx12f_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_470), .A2(n_352), .B1(n_315), .B2(n_345), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_411), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_439), .A2(n_352), .B1(n_315), .B2(n_353), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_473), .A2(n_315), .B1(n_345), .B2(n_329), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_450), .A2(n_15), .B(n_12), .C(n_14), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_431), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_446), .Y(n_560) );
BUFx10_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_472), .A2(n_353), .B(n_379), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_478), .B(n_20), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_480), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_457), .B(n_315), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_480), .A2(n_350), .B1(n_345), .B2(n_329), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_478), .A2(n_483), .B1(n_458), .B2(n_463), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_481), .B(n_21), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_448), .A2(n_353), .B1(n_345), .B2(n_350), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_484), .B(n_329), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_448), .B(n_22), .Y(n_572) );
OAI22x1_ASAP7_75t_L g573 ( .A1(n_461), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_461), .A2(n_24), .B(n_25), .C(n_26), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_462), .B(n_30), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_462), .B(n_31), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_485), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_426), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_414), .B(n_32), .Y(n_579) );
AO22x1_ASAP7_75t_L g580 ( .A1(n_421), .A2(n_33), .B1(n_34), .B2(n_36), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_412), .A2(n_379), .B(n_350), .Y(n_581) );
CKINVDCx8_ASAP7_75t_R g582 ( .A(n_447), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_421), .Y(n_583) );
BUFx8_ASAP7_75t_SL g584 ( .A(n_425), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_459), .A2(n_33), .B(n_34), .C(n_36), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_430), .B(n_37), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_430), .B(n_37), .Y(n_587) );
INVx6_ASAP7_75t_L g588 ( .A(n_418), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_421), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_417), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_412), .A2(n_379), .B(n_350), .Y(n_591) );
INVx3_ASAP7_75t_SL g592 ( .A(n_430), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_417), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_417), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_418), .B(n_38), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_430), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_519), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_519), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_568), .A2(n_88), .B(n_87), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_528), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_528), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_495), .A2(n_379), .B(n_41), .C(n_42), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_549), .A2(n_40), .B1(n_41), .B2(n_44), .Y(n_603) );
BUFx12f_ASAP7_75t_L g604 ( .A(n_544), .Y(n_604) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_573), .A2(n_552), .A3(n_510), .B(n_581), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_518), .A2(n_48), .B(n_49), .C(n_50), .Y(n_606) );
AO31x2_ASAP7_75t_L g607 ( .A1(n_591), .A2(n_49), .A3(n_50), .B(n_53), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_568), .A2(n_91), .B(n_90), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_583), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_492), .A2(n_93), .B(n_92), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_563), .A2(n_102), .B(n_98), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_528), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_579), .Y(n_613) );
BUFx2_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_523), .B(n_54), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_571), .A2(n_104), .B(n_103), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_502), .A2(n_527), .B(n_566), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_508), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_585), .A2(n_59), .B(n_60), .C(n_61), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_523), .Y(n_620) );
AO32x2_ASAP7_75t_L g621 ( .A1(n_556), .A2(n_59), .A3(n_61), .B1(n_63), .B2(n_64), .Y(n_621) );
BUFx3_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_589), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_564), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_535), .A2(n_65), .B1(n_67), .B2(n_68), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_501), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_497), .B(n_72), .Y(n_627) );
AO32x2_ASAP7_75t_L g628 ( .A1(n_570), .A2(n_72), .A3(n_73), .B1(n_74), .B2(n_75), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_537), .B(n_110), .Y(n_629) );
INVx3_ASAP7_75t_SL g630 ( .A(n_588), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_509), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_522), .A2(n_77), .B(n_78), .C(n_80), .Y(n_632) );
CKINVDCx11_ASAP7_75t_R g633 ( .A(n_582), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_537), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_514), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_490), .B(n_81), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_521), .Y(n_637) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_520), .A2(n_157), .B(n_200), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_511), .B(n_82), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_548), .A2(n_83), .B1(n_111), .B2(n_112), .Y(n_640) );
AO21x1_ASAP7_75t_L g641 ( .A1(n_533), .A2(n_160), .B(n_113), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_561), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_588), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_561), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_537), .Y(n_645) );
BUFx10_ASAP7_75t_L g646 ( .A(n_595), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_595), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_519), .Y(n_648) );
AO31x2_ASAP7_75t_L g649 ( .A1(n_575), .A2(n_116), .A3(n_118), .B(n_119), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_541), .B(n_122), .Y(n_650) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_496), .Y(n_651) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_542), .A2(n_125), .A3(n_126), .B(n_127), .Y(n_652) );
AO31x2_ASAP7_75t_L g653 ( .A1(n_569), .A2(n_128), .A3(n_130), .B(n_131), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_531), .Y(n_654) );
OAI22xp33_ASAP7_75t_SL g655 ( .A1(n_546), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_590), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_593), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_594), .Y(n_658) );
AOI221xp5_ASAP7_75t_SL g659 ( .A1(n_558), .A2(n_534), .B1(n_540), .B2(n_526), .C(n_574), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_586), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_494), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_532), .A2(n_159), .B(n_161), .C(n_162), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_555), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_524), .A2(n_507), .B(n_506), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_503), .A2(n_168), .B(n_170), .Y(n_665) );
BUFx8_ASAP7_75t_L g666 ( .A(n_587), .Y(n_666) );
CKINVDCx11_ASAP7_75t_R g667 ( .A(n_491), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_559), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_504), .B(n_174), .Y(n_669) );
INVx3_ASAP7_75t_SL g670 ( .A(n_529), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_505), .A2(n_512), .B(n_516), .C(n_538), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_577), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_565), .A2(n_175), .B1(n_176), .B2(n_178), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_530), .B(n_182), .Y(n_674) );
BUFx10_ASAP7_75t_L g675 ( .A(n_539), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_498), .Y(n_676) );
O2A1O1Ixp5_ASAP7_75t_L g677 ( .A1(n_539), .A2(n_183), .B(n_184), .C(n_186), .Y(n_677) );
AO31x2_ASAP7_75t_L g678 ( .A1(n_560), .A2(n_187), .A3(n_188), .B(n_190), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_541), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_580), .A2(n_193), .B1(n_195), .B2(n_197), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_562), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_499), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_550), .Y(n_683) );
INVx8_ASAP7_75t_L g684 ( .A(n_496), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_515), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_536), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_496), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_578), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_513), .B(n_551), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_572), .B(n_576), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_500), .A2(n_543), .B(n_547), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_545), .A2(n_554), .B(n_557), .C(n_567), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_554), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_517), .A2(n_535), .B1(n_549), .B2(n_373), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_568), .A2(n_474), .B(n_427), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_535), .A2(n_425), .B1(n_449), .B2(n_444), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g698 ( .A1(n_568), .A2(n_474), .B(n_427), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_519), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_596), .B(n_414), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_SL g701 ( .A1(n_493), .A2(n_552), .B(n_510), .C(n_525), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_495), .A2(n_518), .B(n_585), .C(n_414), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_592), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_701), .A2(n_702), .B(n_617), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_633), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_656), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_700), .B(n_697), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_696), .A2(n_698), .B(n_613), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_664), .A2(n_671), .B(n_691), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_623), .B(n_609), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_624), .B(n_626), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_703), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_631), .B(n_635), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_658), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_637), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_620), .B(n_639), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_654), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_647), .B(n_646), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_657), .B(n_660), .Y(n_719) );
CKINVDCx8_ASAP7_75t_R g720 ( .A(n_614), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_646), .B(n_627), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_629), .A2(n_636), .B(n_674), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_682), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_681), .B(n_672), .Y(n_724) );
AND2x6_ASAP7_75t_L g725 ( .A(n_690), .B(n_597), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_663), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_630), .B(n_622), .Y(n_727) );
BUFx4f_ASAP7_75t_SL g728 ( .A(n_604), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_668), .Y(n_729) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_634), .B(n_645), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_695), .A2(n_640), .B1(n_692), .B2(n_680), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_618), .B(n_695), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_685), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_625), .A2(n_615), .B1(n_632), .B2(n_619), .C(n_606), .Y(n_734) );
AO31x2_ASAP7_75t_L g735 ( .A1(n_602), .A2(n_694), .A3(n_693), .B(n_662), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_643), .B(n_670), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_688), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_607), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_666), .B(n_687), .Y(n_739) );
BUFx12f_ASAP7_75t_L g740 ( .A(n_667), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_686), .B(n_675), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_676), .A2(n_661), .B1(n_669), .B2(n_612), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_679), .B(n_601), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_679), .B(n_600), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_621), .B(n_628), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_677), .A2(n_659), .B(n_610), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_621), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_689), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_605), .B(n_659), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_605), .B(n_683), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_684), .Y(n_751) );
BUFx3_ASAP7_75t_L g752 ( .A(n_684), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_597), .B(n_598), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_665), .A2(n_611), .B(n_616), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_651), .B(n_598), .Y(n_755) );
AO21x1_ASAP7_75t_L g756 ( .A1(n_655), .A2(n_650), .B(n_673), .Y(n_756) );
AO31x2_ASAP7_75t_L g757 ( .A1(n_649), .A2(n_605), .A3(n_653), .B(n_652), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_648), .B(n_699), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_628), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_648), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_628), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_649), .B(n_653), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_678), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_652), .A2(n_701), .B(n_702), .Y(n_764) );
BUFx12f_ASAP7_75t_L g765 ( .A(n_678), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_678), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_652), .B(n_696), .Y(n_767) );
AO31x2_ASAP7_75t_L g768 ( .A1(n_641), .A2(n_702), .A3(n_602), .B(n_603), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_656), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_656), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_659), .B(n_619), .C(n_702), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_656), .Y(n_772) );
INVx3_ASAP7_75t_L g773 ( .A(n_634), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_700), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g775 ( .A1(n_702), .A2(n_613), .B(n_585), .C(n_495), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_703), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_700), .B(n_535), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_656), .Y(n_778) );
CKINVDCx6p67_ASAP7_75t_R g779 ( .A(n_703), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_642), .B(n_644), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_703), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_633), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_700), .B(n_592), .Y(n_783) );
OA21x2_ASAP7_75t_L g784 ( .A1(n_599), .A2(n_608), .B(n_638), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_642), .B(n_644), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_703), .Y(n_786) );
BUFx8_ASAP7_75t_SL g787 ( .A(n_604), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_696), .A2(n_698), .B(n_702), .Y(n_788) );
AO31x2_ASAP7_75t_L g789 ( .A1(n_641), .A2(n_702), .A3(n_602), .B(n_603), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_656), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_700), .B(n_535), .Y(n_791) );
INVx1_ASAP7_75t_SL g792 ( .A(n_623), .Y(n_792) );
AO21x2_ASAP7_75t_L g793 ( .A1(n_764), .A2(n_762), .B(n_709), .Y(n_793) );
INVx4_ASAP7_75t_L g794 ( .A(n_725), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_738), .Y(n_795) );
OR2x6_ASAP7_75t_L g796 ( .A(n_731), .B(n_708), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_783), .Y(n_797) );
AO21x2_ASAP7_75t_L g798 ( .A1(n_767), .A2(n_746), .B(n_704), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_707), .B(n_706), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_775), .A2(n_771), .B(n_734), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_714), .B(n_769), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_759), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_748), .B(n_777), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_770), .B(n_772), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_752), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_791), .B(n_774), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_732), .A2(n_788), .B1(n_756), .B2(n_742), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_747), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_778), .B(n_790), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_716), .B(n_792), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_724), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_765), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_750), .Y(n_813) );
OA21x2_ASAP7_75t_L g814 ( .A1(n_763), .A2(n_766), .B(n_749), .Y(n_814) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_711), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_711), .B(n_715), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_750), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_719), .B(n_713), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_745), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_758), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_726), .B(n_729), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_717), .B(n_744), .Y(n_822) );
OR2x6_ASAP7_75t_L g823 ( .A(n_773), .B(n_722), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_725), .Y(n_824) );
INVxp67_ASAP7_75t_L g825 ( .A(n_786), .Y(n_825) );
BUFx2_ASAP7_75t_L g826 ( .A(n_758), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_723), .B(n_737), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_733), .B(n_773), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_761), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_730), .B(n_743), .Y(n_830) );
AOI31xp33_ASAP7_75t_L g831 ( .A1(n_705), .A2(n_782), .A3(n_721), .B(n_739), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_761), .Y(n_832) );
NOR2x1_ASAP7_75t_R g833 ( .A(n_740), .B(n_728), .Y(n_833) );
AO21x2_ASAP7_75t_L g834 ( .A1(n_754), .A2(n_753), .B(n_757), .Y(n_834) );
NOR2x1_ASAP7_75t_SL g835 ( .A(n_760), .B(n_751), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g836 ( .A1(n_776), .A2(n_781), .B1(n_712), .B2(n_741), .C(n_718), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_743), .B(n_735), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_735), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_780), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_785), .Y(n_840) );
BUFx3_ASAP7_75t_L g841 ( .A(n_725), .Y(n_841) );
BUFx2_ASAP7_75t_L g842 ( .A(n_725), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_735), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_727), .B(n_736), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_768), .B(n_789), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_768), .B(n_789), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_784), .A2(n_755), .B(n_768), .Y(n_847) );
OAI21xp33_ASAP7_75t_L g848 ( .A1(n_789), .A2(n_720), .B(n_779), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_787), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_707), .B(n_706), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_707), .B(n_706), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_707), .B(n_706), .Y(n_852) );
OR2x2_ASAP7_75t_L g853 ( .A(n_748), .B(n_707), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_738), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_710), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_707), .B(n_706), .Y(n_856) );
INVx4_ASAP7_75t_L g857 ( .A(n_725), .Y(n_857) );
INVx1_ASAP7_75t_SL g858 ( .A(n_805), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_819), .B(n_796), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_806), .B(n_818), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_795), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_795), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_855), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_819), .B(n_796), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_796), .B(n_799), .Y(n_865) );
INVx5_ASAP7_75t_L g866 ( .A(n_794), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_818), .B(n_799), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_839), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_796), .B(n_850), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_796), .B(n_850), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_851), .B(n_852), .Y(n_871) );
OR2x6_ASAP7_75t_L g872 ( .A(n_794), .B(n_857), .Y(n_872) );
OR2x2_ASAP7_75t_L g873 ( .A(n_853), .B(n_815), .Y(n_873) );
INVx2_ASAP7_75t_SL g874 ( .A(n_842), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_851), .B(n_852), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_856), .B(n_845), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_856), .B(n_845), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_846), .B(n_802), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_803), .B(n_827), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_840), .Y(n_880) );
INVx1_ASAP7_75t_SL g881 ( .A(n_805), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_803), .B(n_820), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_820), .B(n_826), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_844), .B(n_797), .Y(n_884) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_800), .B(n_807), .C(n_848), .Y(n_885) );
INVx1_ASAP7_75t_SL g886 ( .A(n_826), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_846), .B(n_802), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_808), .B(n_854), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_830), .A2(n_857), .B1(n_824), .B2(n_841), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_808), .B(n_854), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_837), .B(n_813), .Y(n_891) );
AND2x4_ASAP7_75t_L g892 ( .A(n_837), .B(n_817), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_823), .B(n_829), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_814), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_811), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_814), .Y(n_896) );
AOI22x1_ASAP7_75t_L g897 ( .A1(n_857), .A2(n_842), .B1(n_812), .B2(n_828), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_836), .A2(n_848), .B1(n_810), .B2(n_830), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_827), .B(n_809), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_801), .B(n_809), .Y(n_900) );
INVx1_ASAP7_75t_SL g901 ( .A(n_858), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_895), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_876), .B(n_843), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_871), .B(n_811), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_876), .B(n_843), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_877), .B(n_838), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_861), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_871), .B(n_822), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_861), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_875), .B(n_822), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_862), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_875), .B(n_816), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_877), .B(n_838), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_899), .B(n_804), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_862), .Y(n_915) );
INVx4_ASAP7_75t_L g916 ( .A(n_866), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_878), .B(n_832), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_878), .B(n_832), .Y(n_918) );
INVx5_ASAP7_75t_L g919 ( .A(n_872), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_882), .B(n_798), .Y(n_920) );
INVx1_ASAP7_75t_SL g921 ( .A(n_881), .Y(n_921) );
INVx1_ASAP7_75t_SL g922 ( .A(n_900), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_887), .B(n_847), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_882), .B(n_798), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_873), .B(n_798), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_887), .B(n_847), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_899), .B(n_804), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_900), .B(n_801), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_866), .Y(n_929) );
CKINVDCx16_ASAP7_75t_R g930 ( .A(n_884), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_886), .Y(n_931) );
AND2x4_ASAP7_75t_L g932 ( .A(n_859), .B(n_823), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_859), .B(n_847), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_864), .B(n_834), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_867), .B(n_821), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_883), .B(n_793), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_864), .B(n_834), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_860), .B(n_849), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_879), .B(n_793), .Y(n_939) );
INVx3_ASAP7_75t_L g940 ( .A(n_872), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_863), .B(n_821), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_886), .B(n_793), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_923), .B(n_865), .Y(n_943) );
INVx2_ASAP7_75t_SL g944 ( .A(n_919), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_923), .B(n_869), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_907), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_907), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_926), .B(n_869), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_922), .B(n_868), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_908), .B(n_880), .Y(n_950) );
OR2x2_ASAP7_75t_L g951 ( .A(n_920), .B(n_891), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_920), .B(n_891), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_924), .B(n_891), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_924), .B(n_891), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_909), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_909), .Y(n_956) );
INVx1_ASAP7_75t_SL g957 ( .A(n_901), .Y(n_957) );
INVx2_ASAP7_75t_SL g958 ( .A(n_919), .Y(n_958) );
NAND2x1p5_ASAP7_75t_L g959 ( .A(n_916), .B(n_866), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_926), .B(n_870), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_911), .Y(n_961) );
OAI21x1_ASAP7_75t_SL g962 ( .A1(n_916), .A2(n_897), .B(n_898), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_903), .B(n_870), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_925), .B(n_892), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_925), .B(n_892), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_905), .B(n_888), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_910), .B(n_888), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_940), .B(n_893), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_906), .B(n_890), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_906), .B(n_890), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_913), .B(n_894), .Y(n_971) );
NAND2x1p5_ASAP7_75t_L g972 ( .A(n_919), .B(n_866), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_913), .B(n_912), .Y(n_973) );
INVx2_ASAP7_75t_SL g974 ( .A(n_919), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_915), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_933), .B(n_894), .Y(n_976) );
INVxp67_ASAP7_75t_L g977 ( .A(n_902), .Y(n_977) );
INVxp67_ASAP7_75t_L g978 ( .A(n_938), .Y(n_978) );
AND2x4_ASAP7_75t_SL g979 ( .A(n_940), .B(n_872), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_933), .B(n_896), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_943), .B(n_934), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_943), .B(n_934), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_946), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_946), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_966), .B(n_939), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g986 ( .A(n_957), .B(n_930), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_945), .B(n_937), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_973), .B(n_939), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_947), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_945), .B(n_937), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_947), .Y(n_991) );
OAI332xp33_ASAP7_75t_L g992 ( .A1(n_950), .A2(n_941), .A3(n_904), .B1(n_935), .B2(n_921), .B3(n_936), .C1(n_927), .C2(n_914), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_948), .B(n_917), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_948), .B(n_917), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_962), .A2(n_919), .B(n_897), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_955), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_976), .B(n_936), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_955), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_956), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_956), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_966), .B(n_928), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_960), .B(n_918), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_969), .B(n_931), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_978), .B(n_831), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_961), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_968), .B(n_940), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_960), .B(n_918), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_977), .B(n_885), .C(n_825), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_992), .B(n_969), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_983), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_983), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_993), .B(n_970), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_981), .B(n_963), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g1014 ( .A(n_986), .Y(n_1014) );
A2O1A1Ixp33_ASAP7_75t_L g1015 ( .A1(n_1004), .A2(n_979), .B(n_944), .C(n_974), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_981), .B(n_963), .Y(n_1016) );
NAND2x1p5_ASAP7_75t_L g1017 ( .A(n_995), .B(n_929), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_988), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_993), .B(n_970), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_988), .Y(n_1020) );
AOI221x1_ASAP7_75t_SL g1021 ( .A1(n_1008), .A2(n_949), .B1(n_967), .B2(n_968), .C(n_975), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_994), .B(n_976), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_989), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_1001), .B(n_833), .Y(n_1024) );
INVxp67_ASAP7_75t_L g1025 ( .A(n_1003), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_989), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_991), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_994), .B(n_980), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_991), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1009), .B(n_1002), .Y(n_1030) );
INVxp67_ASAP7_75t_L g1031 ( .A(n_1014), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1018), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1021), .B(n_1002), .Y(n_1033) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_1017), .A2(n_959), .B1(n_974), .B2(n_944), .Y(n_1034) );
INVxp67_ASAP7_75t_SL g1035 ( .A(n_1017), .Y(n_1035) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_1017), .A2(n_958), .B1(n_972), .B2(n_929), .Y(n_1036) );
O2A1O1Ixp5_ASAP7_75t_L g1037 ( .A1(n_1015), .A2(n_1006), .B(n_985), .C(n_999), .Y(n_1037) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_1015), .A2(n_962), .B(n_972), .Y(n_1038) );
AOI321xp33_ASAP7_75t_L g1039 ( .A1(n_1024), .A2(n_1006), .A3(n_968), .B1(n_987), .B2(n_982), .C(n_990), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_1012), .A2(n_997), .B1(n_958), .B2(n_1007), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1020), .B(n_1007), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1025), .A2(n_980), .B1(n_968), .B2(n_971), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_1019), .A2(n_997), .B1(n_965), .B2(n_964), .Y(n_1043) );
NOR3xp33_ASAP7_75t_L g1044 ( .A(n_1037), .B(n_1011), .C(n_1026), .Y(n_1044) );
AOI21xp5_ASAP7_75t_L g1045 ( .A1(n_1036), .A2(n_1022), .B(n_1028), .Y(n_1045) );
AOI211xp5_ASAP7_75t_L g1046 ( .A1(n_1036), .A2(n_1013), .B(n_1016), .C(n_1026), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_1033), .A2(n_1031), .B1(n_1030), .B2(n_1043), .C(n_1040), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1042), .Y(n_1048) );
NAND4xp25_ASAP7_75t_SL g1049 ( .A(n_1038), .B(n_889), .C(n_990), .D(n_987), .Y(n_1049) );
AOI211xp5_ASAP7_75t_L g1050 ( .A1(n_1034), .A2(n_1029), .B(n_1027), .C(n_1023), .Y(n_1050) );
NOR2xp33_ASAP7_75t_SL g1051 ( .A(n_1035), .B(n_866), .Y(n_1051) );
OAI311xp33_ASAP7_75t_L g1052 ( .A1(n_1039), .A2(n_965), .A3(n_964), .B1(n_951), .C1(n_954), .Y(n_1052) );
AND4x1_ASAP7_75t_L g1053 ( .A(n_1047), .B(n_1032), .C(n_1041), .D(n_982), .Y(n_1053) );
NOR2x1p5_ASAP7_75t_L g1054 ( .A(n_1049), .B(n_824), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1044), .B(n_1010), .Y(n_1055) );
AOI211x1_ASAP7_75t_L g1056 ( .A1(n_1045), .A2(n_984), .B(n_998), .C(n_1005), .Y(n_1056) );
OAI321xp33_ASAP7_75t_L g1057 ( .A1(n_1046), .A2(n_874), .A3(n_942), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1048), .B(n_1010), .Y(n_1058) );
NOR3xp33_ASAP7_75t_SL g1059 ( .A(n_1057), .B(n_1052), .C(n_1051), .Y(n_1059) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_1058), .A2(n_1050), .B(n_1000), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1056), .B(n_996), .Y(n_1061) );
NOR2x1_ASAP7_75t_L g1062 ( .A(n_1054), .B(n_857), .Y(n_1062) );
OR2x6_ASAP7_75t_L g1063 ( .A(n_1062), .B(n_1055), .Y(n_1063) );
CKINVDCx16_ASAP7_75t_R g1064 ( .A(n_1061), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1059), .Y(n_1065) );
XNOR2xp5_ASAP7_75t_L g1066 ( .A(n_1060), .B(n_1053), .Y(n_1066) );
INVx3_ASAP7_75t_L g1067 ( .A(n_1063), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1063), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_1065), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1068), .B(n_1064), .Y(n_1070) );
AND2x4_ASAP7_75t_L g1071 ( .A(n_1067), .B(n_1055), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_1067), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1071), .A2(n_1066), .B1(n_1069), .B2(n_1068), .Y(n_1073) );
OAI21x1_ASAP7_75t_SL g1074 ( .A1(n_1071), .A2(n_1067), .B(n_835), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1073), .B(n_1070), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1076 ( .A1(n_1074), .A2(n_1072), .B(n_835), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_1075), .A2(n_828), .B(n_841), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_1077), .A2(n_1076), .B1(n_932), .B2(n_971), .Y(n_1078) );
endmodule