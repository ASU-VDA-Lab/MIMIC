module fake_jpeg_27465_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_29),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_40),
.B1(n_28),
.B2(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_17),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_30),
.B1(n_21),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_16),
.B1(n_33),
.B2(n_34),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_29),
.B1(n_31),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_61),
.B1(n_16),
.B2(n_33),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_77),
.Y(n_113)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_70),
.B(n_74),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_87),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_86),
.B1(n_98),
.B2(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_40),
.B1(n_43),
.B2(n_42),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_103),
.B1(n_42),
.B2(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_26),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_86)
);

OA22x2_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_92),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

OA22x2_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_43),
.B1(n_42),
.B2(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_44),
.C(n_41),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_119),
.C(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_111),
.B1(n_126),
.B2(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_23),
.B1(n_32),
.B2(n_28),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_36),
.B1(n_41),
.B2(n_44),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_44),
.B1(n_41),
.B2(n_73),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_104),
.C(n_67),
.Y(n_119)
);

AOI22x1_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_36),
.B1(n_27),
.B2(n_26),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_136),
.B(n_137),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_23),
.B1(n_32),
.B2(n_24),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_19),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_32),
.B(n_24),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_152),
.B1(n_117),
.B2(n_122),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_87),
.B1(n_96),
.B2(n_83),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_148),
.B1(n_114),
.B2(n_128),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_69),
.B1(n_80),
.B2(n_106),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_145),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_149),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_87),
.B1(n_78),
.B2(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_155),
.B1(n_118),
.B2(n_126),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_150),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_44),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_160),
.B(n_163),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_108),
.B1(n_121),
.B2(n_113),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_36),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_72),
.B1(n_24),
.B2(n_78),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_161),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_26),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_44),
.C(n_41),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_100),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_129),
.B1(n_116),
.B2(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_115),
.B1(n_121),
.B2(n_120),
.Y(n_169)
);

OAI22x1_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_180),
.B1(n_159),
.B2(n_14),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_189),
.B1(n_198),
.B2(n_143),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_118),
.B1(n_123),
.B2(n_117),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_182),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_111),
.B(n_128),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_190),
.B(n_0),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_173),
.B1(n_183),
.B2(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_193),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_165),
.C(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_114),
.B1(n_123),
.B2(n_131),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_133),
.B(n_1),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_75),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_133),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_130),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_138),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_171),
.B1(n_189),
.B2(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_206),
.B1(n_216),
.B2(n_168),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_145),
.B(n_151),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_207),
.B(n_210),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_211),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_147),
.B1(n_150),
.B2(n_163),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_147),
.B(n_153),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_44),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_168),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_222),
.Y(n_231)
);

AOI22x1_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_3),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_13),
.B(n_12),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_178),
.B(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_14),
.B(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_9),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_2),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_0),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_0),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_206),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_1),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_207),
.B(n_214),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_186),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_253),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_179),
.C(n_175),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_239),
.C(n_230),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_179),
.C(n_170),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_228),
.B(n_223),
.C(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_208),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_195),
.Y(n_253)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_258),
.B(n_232),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_210),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_267),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_234),
.B(n_246),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_245),
.C(n_233),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_274),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_242),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_230),
.C(n_210),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_275),
.C(n_240),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_202),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_240),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_226),
.B1(n_204),
.B2(n_201),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_233),
.B1(n_209),
.B2(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_208),
.C(n_207),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_276),
.A2(n_260),
.B1(n_268),
.B2(n_265),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_238),
.CI(n_235),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_281),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_258),
.B(n_262),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_195),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_284),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_264),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_243),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_260),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_241),
.C(n_209),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_289),
.C(n_227),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_241),
.C(n_222),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_262),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_263),
.CI(n_275),
.CON(n_299),
.SN(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_270),
.CI(n_273),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_304),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_261),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_277),
.B(n_227),
.CI(n_252),
.CON(n_305),
.SN(n_305)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_282),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_287),
.B1(n_276),
.B2(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_289),
.C(n_283),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_314),
.C(n_310),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_284),
.B1(n_290),
.B2(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_315),
.B1(n_299),
.B2(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_297),
.C(n_307),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_318),
.B(n_319),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_298),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_322),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_295),
.B(n_300),
.Y(n_321)
);

O2A1O1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_324),
.B(n_312),
.C(n_317),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_310),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_320),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_299),
.B(n_303),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_326),
.A2(n_314),
.B(n_305),
.C(n_309),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_286),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_330),
.B(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_277),
.C(n_4),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_7),
.B(n_4),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_3),
.B(n_5),
.Y(n_336)
);


endmodule