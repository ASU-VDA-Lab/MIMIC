module fake_jpeg_2217_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_9),
.C(n_5),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_37),
.B1(n_50),
.B2(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_66),
.B1(n_48),
.B2(n_42),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_50),
.B1(n_49),
.B2(n_43),
.Y(n_66)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_55),
.C(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_68),
.B1(n_61),
.B2(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_56),
.B1(n_53),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_92),
.B1(n_96),
.B2(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_98),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_8),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

CKINVDCx10_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_105),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_23),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_92),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_19),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_116),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_20),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_10),
.B1(n_11),
.B2(n_17),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_21),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_130),
.C(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_36),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_113),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_133),
.B(n_127),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_115),
.B(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_137),
.A2(n_140),
.B1(n_118),
.B2(n_117),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_129),
.B1(n_119),
.B2(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_128),
.C(n_134),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_139),
.B1(n_131),
.B2(n_125),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_124),
.B(n_104),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_26),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_28),
.B(n_30),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_32),
.Y(n_149)
);


endmodule