module fake_jpeg_30585_n_174 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_78),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_0),
.CON(n_71),
.SN(n_71)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_0),
.Y(n_88)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_57),
.B1(n_43),
.B2(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_93),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_52),
.B1(n_62),
.B2(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_63),
.B1(n_61),
.B2(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_99),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_103),
.Y(n_126)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_77),
.B1(n_65),
.B2(n_46),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_76),
.B1(n_73),
.B2(n_47),
.Y(n_120)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_77),
.B1(n_72),
.B2(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_129),
.B1(n_135),
.B2(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_66),
.B(n_60),
.C(n_48),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_52),
.B1(n_51),
.B2(n_3),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_133),
.B1(n_139),
.B2(n_11),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_102),
.B1(n_98),
.B2(n_101),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_52),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_13),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_42),
.B1(n_22),
.B2(n_23),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_40),
.B1(n_24),
.B2(n_25),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_7),
.C(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_10),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_132),
.C(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_14),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_153),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_128),
.B1(n_120),
.B2(n_136),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_15),
.B(n_16),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_15),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_139),
.B1(n_131),
.B2(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_142),
.C(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_165),
.C(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_142),
.A3(n_153),
.B1(n_156),
.B2(n_158),
.C1(n_157),
.C2(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_152),
.B(n_144),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_133),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_140),
.C(n_135),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_17),
.C(n_18),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_21),
.Y(n_174)
);


endmodule