module fake_jpeg_12762_n_581 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_581);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_581;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g185 ( 
.A(n_64),
.Y(n_185)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_71),
.B(n_106),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_74),
.Y(n_150)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_2),
.C(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_81),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_80),
.B(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_22),
.B(n_2),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_82),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_97),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_22),
.B(n_3),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_94),
.B(n_108),
.Y(n_167)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_104),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_30),
.B(n_5),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_18),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_114),
.Y(n_159)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_118),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_5),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_123),
.Y(n_153)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_5),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_56),
.B(n_17),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_126),
.Y(n_166)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_6),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_6),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_49),
.B1(n_36),
.B2(n_40),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_131),
.B(n_141),
.C(n_165),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_51),
.B1(n_45),
.B2(n_40),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_147),
.B1(n_107),
.B2(n_23),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_137),
.B(n_143),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_45),
.B1(n_35),
.B2(n_21),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_51),
.B1(n_35),
.B2(n_21),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_75),
.A2(n_51),
.B1(n_54),
.B2(n_28),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_151),
.A2(n_162),
.B1(n_158),
.B2(n_200),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_54),
.B1(n_46),
.B2(n_39),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_154),
.A2(n_160),
.B1(n_158),
.B2(n_210),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_155),
.B(n_172),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_101),
.A2(n_46),
.B1(n_39),
.B2(n_38),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_84),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_87),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_173),
.B(n_177),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_37),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_31),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_178),
.B(n_180),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_31),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_63),
.B(n_29),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_182),
.B(n_183),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_70),
.B(n_29),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_64),
.A2(n_28),
.B(n_26),
.C(n_67),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_23),
.B(n_8),
.C(n_10),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_91),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_200),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_73),
.B(n_7),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_196),
.B(n_201),
.CI(n_193),
.CON(n_248),
.SN(n_248)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_83),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_88),
.B(n_35),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_206),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_98),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_105),
.B(n_21),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_161),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_212),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_213),
.Y(n_289)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_215),
.B(n_217),
.C(n_226),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_216),
.B(n_223),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_137),
.A2(n_116),
.B1(n_112),
.B2(n_109),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_220),
.Y(n_339)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_153),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_222),
.B(n_230),
.C(n_235),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_159),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_224),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_227),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_143),
.A2(n_23),
.B1(n_8),
.B2(n_9),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_229),
.A2(n_245),
.B(n_250),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_7),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_10),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_234),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_155),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_144),
.B(n_10),
.Y(n_235)
);

AOI22x1_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_23),
.B1(n_12),
.B2(n_13),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_236),
.A2(n_275),
.B1(n_169),
.B2(n_150),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_11),
.B(n_12),
.C(n_14),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_237),
.B(n_272),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_171),
.Y(n_238)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_239),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_131),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_240),
.A2(n_242),
.B1(n_261),
.B2(n_266),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_132),
.A2(n_167),
.B1(n_141),
.B2(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_169),
.A2(n_190),
.B1(n_138),
.B2(n_149),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_244),
.A2(n_253),
.B1(n_256),
.B2(n_279),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_157),
.A2(n_184),
.B1(n_181),
.B2(n_190),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_146),
.B(n_163),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_276),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_248),
.B(n_252),
.Y(n_316)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_157),
.A2(n_181),
.B1(n_190),
.B2(n_188),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_176),
.A2(n_210),
.B1(n_160),
.B2(n_179),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_254),
.Y(n_310)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_135),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_255),
.Y(n_326)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_257),
.B(n_269),
.Y(n_299)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_258),
.B(n_259),
.Y(n_329)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_170),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_175),
.C(n_150),
.Y(n_292)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_175),
.Y(n_262)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_263),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_152),
.A2(n_204),
.B1(n_193),
.B2(n_201),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_267),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_152),
.A2(n_204),
.B1(n_202),
.B2(n_198),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_271),
.A2(n_280),
.B1(n_130),
.B2(n_171),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_179),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_192),
.A2(n_202),
.B1(n_209),
.B2(n_145),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_172),
.B(n_199),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_209),
.A2(n_170),
.B1(n_148),
.B2(n_140),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_142),
.A2(n_195),
.B1(n_187),
.B2(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_142),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_282),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_130),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_285),
.A2(n_301),
.B1(n_317),
.B2(n_320),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_305),
.C(n_306),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_256),
.A2(n_187),
.B1(n_186),
.B2(n_148),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_SL g305 ( 
.A(n_222),
.B(n_211),
.C(n_164),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_234),
.B(n_186),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_211),
.C(n_135),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_312),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_264),
.B(n_233),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_314),
.A2(n_337),
.B1(n_231),
.B2(n_255),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_223),
.A2(n_156),
.B1(n_189),
.B2(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_235),
.B(n_156),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_319),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_189),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_248),
.A2(n_274),
.B1(n_242),
.B2(n_236),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_229),
.A2(n_248),
.B1(n_230),
.B2(n_236),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_323),
.B1(n_213),
.B2(n_215),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_230),
.A2(n_276),
.B1(n_237),
.B2(n_259),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_270),
.A3(n_246),
.B1(n_237),
.B2(n_265),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_325),
.B(n_287),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_251),
.B1(n_275),
.B2(n_225),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_327),
.A2(n_333),
.B1(n_335),
.B2(n_285),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_214),
.B(n_220),
.C(n_243),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_331),
.B(n_217),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_247),
.A2(n_282),
.B(n_212),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_284),
.B(n_315),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_250),
.A2(n_258),
.B1(n_245),
.B2(n_252),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_263),
.A2(n_267),
.B1(n_257),
.B2(n_278),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_260),
.A2(n_277),
.B1(n_281),
.B2(n_283),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_221),
.B(n_249),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_335),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_216),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_340),
.B(n_347),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_341),
.A2(n_343),
.B1(n_361),
.B2(n_366),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_342),
.B(n_367),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_239),
.B1(n_254),
.B2(n_227),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_382),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_260),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_346),
.B(n_351),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_224),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_349),
.Y(n_391)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_226),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_286),
.B(n_232),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_360),
.Y(n_386)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_357),
.Y(n_398)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

INVx6_ASAP7_75t_SL g359 ( 
.A(n_289),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_359),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_238),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_311),
.A2(n_321),
.B1(n_323),
.B2(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_286),
.B(n_238),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_363),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_306),
.B(n_312),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_300),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_365),
.Y(n_406)
);

INVx2_ASAP7_75t_R g365 ( 
.A(n_325),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_311),
.A2(n_307),
.B1(n_320),
.B2(n_324),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_287),
.B(n_338),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_381),
.Y(n_410)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_309),
.B(n_319),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_376),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_318),
.B(n_324),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_378),
.A2(n_303),
.B1(n_310),
.B2(n_326),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_314),
.A2(n_302),
.B1(n_296),
.B2(n_301),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_379),
.A2(n_336),
.B1(n_322),
.B2(n_294),
.Y(n_418)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_334),
.Y(n_382)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_385),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_377),
.A2(n_333),
.B1(n_292),
.B2(n_303),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_403),
.B1(n_409),
.B2(n_379),
.Y(n_434)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_401),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_295),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_407),
.C(n_412),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_326),
.B(n_294),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_404),
.A2(n_374),
.B(n_382),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_290),
.C(n_293),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_377),
.A2(n_295),
.B1(n_334),
.B2(n_330),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_290),
.C(n_293),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_360),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_418),
.A2(n_345),
.B1(n_354),
.B2(n_358),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_414),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_422),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_404),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_372),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_431),
.C(n_436),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_424),
.B(n_442),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_378),
.B(n_369),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_425),
.A2(n_438),
.B(n_439),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_416),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_443),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_340),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_429),
.B(n_430),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_364),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_353),
.C(n_366),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_432),
.A2(n_409),
.B1(n_392),
.B2(n_400),
.Y(n_455)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_353),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_417),
.A2(n_351),
.B(n_365),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_417),
.A2(n_365),
.B(n_352),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_408),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_441),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_380),
.B1(n_362),
.B2(n_347),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_384),
.A2(n_355),
.B(n_361),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_384),
.A2(n_406),
.B(n_387),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_446),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_418),
.B1(n_406),
.B2(n_411),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_388),
.B(n_341),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_413),
.C(n_386),
.Y(n_468)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_349),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_390),
.A2(n_343),
.B1(n_373),
.B2(n_375),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_449),
.A2(n_394),
.B1(n_402),
.B2(n_391),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_436),
.B(n_383),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_463),
.Y(n_485)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_455),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_475),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_386),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_464),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_469),
.C(n_471),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_412),
.C(n_410),
.Y(n_469)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_394),
.C(n_375),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_392),
.Y(n_472)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_473),
.A2(n_446),
.B1(n_441),
.B2(n_462),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_396),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_447),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_396),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_477),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_429),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_426),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_478),
.B(n_480),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_479),
.A2(n_450),
.B1(n_467),
.B2(n_494),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_471),
.B(n_420),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_442),
.Y(n_481)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_443),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_492),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_487),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_419),
.C(n_423),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_495),
.C(n_469),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_465),
.Y(n_489)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_489),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_461),
.A2(n_444),
.B1(n_434),
.B2(n_425),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_491),
.A2(n_500),
.B1(n_501),
.B2(n_467),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_432),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_445),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_475),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_419),
.C(n_447),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_502),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_457),
.A2(n_421),
.B(n_438),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_457),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_461),
.A2(n_449),
.B1(n_422),
.B2(n_443),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_450),
.A2(n_424),
.B1(n_439),
.B2(n_437),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_448),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_477),
.B1(n_494),
.B2(n_497),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_505),
.A2(n_510),
.B1(n_497),
.B2(n_451),
.Y(n_537)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_507),
.Y(n_526)
);

INVx13_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_479),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_511),
.A2(n_500),
.B1(n_491),
.B2(n_483),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_499),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_498),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_514),
.B(n_485),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_483),
.B(n_468),
.CI(n_458),
.CON(n_516),
.SN(n_516)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_519),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_474),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_485),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_454),
.C(n_458),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_520),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_462),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_459),
.C(n_473),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_459),
.C(n_451),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_502),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_525),
.B(n_532),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_SL g527 ( 
.A(n_514),
.B(n_487),
.C(n_486),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_527),
.A2(n_536),
.B(n_512),
.Y(n_547)
);

FAx1_ASAP7_75t_SL g528 ( 
.A(n_518),
.B(n_482),
.CI(n_492),
.CON(n_528),
.SN(n_528)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_528),
.A2(n_535),
.B1(n_516),
.B2(n_470),
.Y(n_551)
);

CKINVDCx14_ASAP7_75t_R g548 ( 
.A(n_530),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_521),
.Y(n_531)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_531),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_534),
.A2(n_538),
.B(n_520),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_482),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_511),
.B1(n_507),
.B2(n_490),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_504),
.A2(n_493),
.B(n_501),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_542),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_504),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_517),
.C(n_522),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_545),
.C(n_550),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_533),
.A2(n_515),
.B(n_519),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_506),
.C(n_510),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_549),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_506),
.C(n_533),
.Y(n_550)
);

AOI322xp5_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_528),
.A3(n_508),
.B1(n_535),
.B2(n_526),
.C1(n_516),
.C2(n_524),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_552),
.A2(n_553),
.B1(n_560),
.B2(n_398),
.Y(n_565)
);

AOI322xp5_ASAP7_75t_L g553 ( 
.A1(n_546),
.A2(n_548),
.A3(n_539),
.B1(n_456),
.B2(n_542),
.C1(n_550),
.C2(n_524),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_546),
.A2(n_549),
.B1(n_531),
.B2(n_543),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_558),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_456),
.C(n_427),
.Y(n_558)
);

AOI322xp5_ASAP7_75t_L g560 ( 
.A1(n_542),
.A2(n_466),
.A3(n_464),
.B1(n_541),
.B2(n_433),
.C1(n_400),
.C2(n_399),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_466),
.B1(n_464),
.B2(n_445),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_393),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_445),
.B1(n_399),
.B2(n_401),
.Y(n_563)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_563),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_564),
.A2(n_565),
.B(n_554),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_555),
.B(n_398),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_566),
.A2(n_567),
.B(n_568),
.Y(n_570)
);

AOI31xp67_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_356),
.A3(n_350),
.B(n_357),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_357),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_555),
.B(n_336),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_569),
.A2(n_568),
.B(n_567),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_572),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_562),
.A2(n_554),
.B(n_342),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_342),
.C(n_322),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_573),
.B(n_322),
.Y(n_575)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_575),
.Y(n_579)
);

OAI211xp5_ASAP7_75t_L g578 ( 
.A1(n_576),
.A2(n_570),
.B(n_342),
.C(n_328),
.Y(n_578)
);

OAI211xp5_ASAP7_75t_L g580 ( 
.A1(n_578),
.A2(n_342),
.B(n_577),
.C(n_288),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_579),
.Y(n_581)
);


endmodule