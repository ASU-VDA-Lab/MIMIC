module real_aes_18265_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_781;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_0), .Y(n_249) );
AND2x4_ASAP7_75t_L g115 ( .A(n_1), .B(n_116), .Y(n_115) );
XNOR2x2_ASAP7_75t_L g859 ( .A(n_2), .B(n_860), .Y(n_859) );
BUFx3_ASAP7_75t_L g190 ( .A(n_3), .Y(n_190) );
INVx1_ASAP7_75t_L g116 ( .A(n_4), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_5), .B(n_902), .Y(n_901) );
XNOR2xp5_ASAP7_75t_L g878 ( .A(n_6), .B(n_29), .Y(n_878) );
AOI22x1_ASAP7_75t_SL g881 ( .A1(n_6), .A2(n_29), .B1(n_882), .B2(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_6), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_7), .B(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g119 ( .A(n_8), .Y(n_119) );
OR2x2_ASAP7_75t_L g130 ( .A(n_8), .B(n_23), .Y(n_130) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_9), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_10), .B(n_184), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_11), .B(n_184), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_12), .B(n_209), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_13), .A2(n_83), .B1(n_159), .B2(n_184), .Y(n_258) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_14), .A2(n_38), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_15), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_16), .B(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_17), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_18), .Y(n_545) );
AO32x2_ASAP7_75t_L g255 ( .A1(n_19), .A2(n_176), .A3(n_177), .B1(n_256), .B2(n_259), .Y(n_255) );
AO32x1_ASAP7_75t_L g293 ( .A1(n_19), .A2(n_176), .A3(n_177), .B1(n_256), .B2(n_259), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_20), .B(n_530), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_21), .B(n_176), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_22), .Y(n_558) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_23), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_24), .A2(n_44), .B1(n_187), .B2(n_199), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_25), .A2(n_91), .B1(n_159), .B2(n_167), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_26), .B(n_166), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_27), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_28), .B(n_222), .Y(n_282) );
INVx1_ASAP7_75t_L g883 ( .A(n_29), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_30), .A2(n_63), .B1(n_167), .B2(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_31), .B(n_184), .Y(n_600) );
INVx2_ASAP7_75t_L g868 ( .A(n_32), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_33), .B(n_163), .Y(n_631) );
INVx1_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
BUFx3_ASAP7_75t_L g871 ( .A(n_34), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_35), .B(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g891 ( .A(n_35), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_36), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_37), .B(n_536), .Y(n_637) );
AND2x2_ASAP7_75t_L g551 ( .A(n_39), .B(n_536), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_40), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_41), .B(n_221), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_42), .B(n_530), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_43), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_45), .B(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_46), .A2(n_78), .B1(n_221), .B2(n_222), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_47), .B(n_264), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_48), .A2(n_200), .B(n_247), .C(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_49), .A2(n_80), .B1(n_159), .B2(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g155 ( .A(n_50), .Y(n_155) );
AND2x4_ASAP7_75t_L g173 ( .A(n_51), .B(n_174), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_52), .A2(n_53), .B1(n_167), .B2(n_187), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_54), .B(n_176), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_55), .B(n_536), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_56), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_57), .B(n_167), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_58), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g174 ( .A(n_59), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_60), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_61), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g171 ( .A(n_62), .B(n_159), .C(n_169), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_64), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_65), .B(n_176), .Y(n_604) );
INVx1_ASAP7_75t_L g875 ( .A(n_66), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_67), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g252 ( .A(n_68), .B(n_253), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_69), .Y(n_268) );
AND2x2_ASAP7_75t_L g909 ( .A(n_70), .B(n_910), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_71), .B(n_163), .C(n_199), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_72), .A2(n_95), .B1(n_184), .B2(n_221), .Y(n_225) );
INVx2_ASAP7_75t_L g164 ( .A(n_73), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_74), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_75), .B(n_528), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_76), .B(n_184), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_77), .B(n_224), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_79), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_81), .B(n_203), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_82), .A2(n_90), .B1(n_530), .B2(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_84), .B(n_184), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_85), .B(n_169), .Y(n_168) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_86), .B(n_162), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_87), .B(n_197), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_88), .A2(n_102), .B1(n_167), .B2(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_89), .B(n_222), .Y(n_279) );
INVx1_ASAP7_75t_SL g860 ( .A(n_92), .Y(n_860) );
INVx1_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_93), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_94), .B(n_209), .Y(n_285) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_96), .B(n_162), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_97), .B(n_536), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_98), .B(n_162), .C(n_224), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_99), .B(n_528), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_100), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_101), .B(n_530), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_122), .B(n_909), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_117), .Y(n_107) );
OR2x6_ASAP7_75t_L g910 ( .A(n_108), .B(n_117), .Y(n_910) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_131), .Y(n_122) );
INVxp67_ASAP7_75t_L g885 ( .A(n_123), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g876 ( .A(n_125), .Y(n_876) );
CKINVDCx8_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g900 ( .A(n_126), .Y(n_900) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_127), .B(n_129), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_129), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2x1_ASAP7_75t_L g908 ( .A(n_130), .B(n_871), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_888), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_863), .B1(n_872), .B2(n_886), .Y(n_132) );
INVx1_ASAP7_75t_L g889 ( .A(n_133), .Y(n_889) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_859), .B1(n_861), .B2(n_862), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B(n_515), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_135), .B(n_139), .Y(n_861) );
INVx8_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx12f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_138), .Y(n_137) );
BUFx8_ASAP7_75t_SL g858 ( .A(n_138), .Y(n_858) );
AND2x2_ASAP7_75t_L g907 ( .A(n_138), .B(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_140), .B(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g884 ( .A(n_140), .Y(n_884) );
OR2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_425), .Y(n_140) );
NAND4xp25_ASAP7_75t_L g141 ( .A(n_142), .B(n_330), .C(n_357), .D(n_393), .Y(n_141) );
AOI221x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_235), .B1(n_269), .B2(n_305), .C(n_309), .Y(n_142) );
NAND3xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_211), .C(n_233), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_178), .Y(n_146) );
INVx2_ASAP7_75t_L g270 ( .A(n_147), .Y(n_270) );
AND2x2_ASAP7_75t_L g443 ( .A(n_147), .B(n_387), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_147), .B(n_234), .Y(n_452) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g458 ( .A(n_148), .Y(n_458) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g303 ( .A(n_149), .Y(n_303) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g386 ( .A(n_150), .B(n_232), .Y(n_386) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_156), .B(n_175), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_151), .A2(n_156), .B(n_175), .Y(n_315) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_151), .A2(n_525), .B(n_535), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_151), .A2(n_556), .B(n_564), .Y(n_555) );
OAI21x1_ASAP7_75t_L g654 ( .A1(n_151), .A2(n_556), .B(n_564), .Y(n_654) );
OAI21xp33_ASAP7_75t_SL g745 ( .A1(n_151), .A2(n_525), .B(n_535), .Y(n_745) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g536 ( .A(n_152), .Y(n_536) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
INVx2_ASAP7_75t_L g230 ( .A(n_153), .Y(n_230) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_165), .B(n_172), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_163), .Y(n_157) );
INVx2_ASAP7_75t_SL g222 ( .A(n_159), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_159), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_160), .Y(n_162) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx1_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
INVx1_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
INVx1_ASAP7_75t_L g247 ( .A(n_160), .Y(n_247) );
INVx3_ASAP7_75t_L g528 ( .A(n_160), .Y(n_528) );
INVx1_ASAP7_75t_L g531 ( .A(n_160), .Y(n_531) );
INVx2_ASAP7_75t_L g563 ( .A(n_162), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_163), .A2(n_183), .B1(n_185), .B2(n_186), .Y(n_182) );
INVx6_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_163), .A2(n_200), .B1(n_257), .B2(n_258), .Y(n_256) );
O2A1O1Ixp5_ASAP7_75t_L g557 ( .A1(n_163), .A2(n_196), .B(n_558), .C(n_559), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_163), .A2(n_602), .B(n_603), .Y(n_601) );
BUFx8_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
INVx2_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_171), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_167), .A2(n_528), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g608 ( .A(n_167), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_167), .A2(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx4f_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
AOI31xp67_ASAP7_75t_L g180 ( .A1(n_172), .A2(n_181), .A3(n_182), .B(n_188), .Y(n_180) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_172), .A2(n_194), .B(n_201), .Y(n_193) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_172), .A2(n_526), .B(n_532), .Y(n_525) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_172), .A2(n_557), .B(n_560), .Y(n_556) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_172), .A2(n_569), .B(n_572), .Y(n_568) );
AND2x4_ASAP7_75t_SL g588 ( .A(n_172), .B(n_177), .Y(n_588) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_172), .A2(n_598), .B(n_601), .Y(n_597) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_172), .A2(n_630), .B(n_633), .Y(n_629) );
BUFx10_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
INVx1_ASAP7_75t_L g251 ( .A(n_173), .Y(n_251) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_173), .A2(n_218), .A3(n_262), .B(n_267), .Y(n_261) );
BUFx10_ASAP7_75t_L g541 ( .A(n_173), .Y(n_541) );
INVx2_ASAP7_75t_L g181 ( .A(n_176), .Y(n_181) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_177), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
BUFx3_ASAP7_75t_L g218 ( .A(n_177), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_177), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g276 ( .A(n_177), .Y(n_276) );
INVx1_ASAP7_75t_SL g567 ( .A(n_177), .Y(n_567) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_178), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_178), .B(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g456 ( .A(n_178), .Y(n_456) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
AND2x2_ASAP7_75t_L g234 ( .A(n_179), .B(n_217), .Y(n_234) );
INVx2_ASAP7_75t_L g312 ( .A(n_179), .Y(n_312) );
AND2x2_ASAP7_75t_L g377 ( .A(n_179), .B(n_315), .Y(n_377) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g232 ( .A(n_180), .Y(n_232) );
INVx3_ASAP7_75t_L g284 ( .A(n_184), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_184), .A2(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g636 ( .A(n_184), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_185), .A2(n_220), .B1(n_223), .B2(n_225), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_185), .A2(n_263), .B1(n_265), .B2(n_266), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_185), .A2(n_282), .B(n_283), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_185), .A2(n_547), .B1(n_607), .B2(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_187), .A2(n_199), .B1(n_243), .B2(n_244), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g304 ( .A(n_191), .Y(n_304) );
AND2x2_ASAP7_75t_L g314 ( .A(n_191), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g376 ( .A(n_191), .B(n_217), .Y(n_376) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_208), .Y(n_191) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_192), .A2(n_193), .B(n_208), .Y(n_214) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_192), .A2(n_597), .B(n_604), .Y(n_596) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_192), .A2(n_629), .B(n_637), .Y(n_628) );
OA21x2_ASAP7_75t_L g640 ( .A1(n_192), .A2(n_629), .B(n_637), .Y(n_640) );
OAI21x1_ASAP7_75t_L g643 ( .A1(n_192), .A2(n_597), .B(n_604), .Y(n_643) );
O2A1O1Ixp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_198), .C(n_200), .Y(n_194) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_200), .A2(n_527), .B(n_529), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_200), .A2(n_573), .B(n_574), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_200), .A2(n_582), .B(n_583), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_200), .A2(n_599), .B(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B1(n_206), .B2(n_207), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_203), .A2(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_204), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_584) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx3_ASAP7_75t_L g250 ( .A(n_205), .Y(n_250) );
INVx2_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
NOR2xp67_ASAP7_75t_SL g539 ( .A(n_209), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_210), .A2(n_541), .A3(n_606), .B(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g341 ( .A(n_211), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_213), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_213), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_213), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_213), .B(n_411), .Y(n_418) );
INVx2_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g387 ( .A(n_214), .B(n_362), .Y(n_387) );
OR2x2_ASAP7_75t_L g389 ( .A(n_214), .B(n_315), .Y(n_389) );
INVx1_ASAP7_75t_L g448 ( .A(n_214), .Y(n_448) );
BUFx2_ASAP7_75t_L g462 ( .A(n_214), .Y(n_462) );
OR2x2_ASAP7_75t_L g490 ( .A(n_214), .B(n_217), .Y(n_490) );
INVx1_ASAP7_75t_L g509 ( .A(n_215), .Y(n_509) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g356 ( .A(n_216), .Y(n_356) );
OR2x2_ASAP7_75t_L g369 ( .A(n_216), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g388 ( .A(n_216), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_231), .Y(n_216) );
INVx2_ASAP7_75t_L g308 ( .A(n_217), .Y(n_308) );
AND2x2_ASAP7_75t_L g324 ( .A(n_217), .B(n_231), .Y(n_324) );
INVx1_ASAP7_75t_L g362 ( .A(n_217), .Y(n_362) );
INVx1_ASAP7_75t_L g405 ( .A(n_217), .Y(n_405) );
AND2x2_ASAP7_75t_L g447 ( .A(n_217), .B(n_448), .Y(n_447) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .A3(n_226), .B(n_228), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_221), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g245 ( .A(n_224), .Y(n_245) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_SL g259 ( .A(n_227), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g253 ( .A(n_230), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_230), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g503 ( .A(n_233), .Y(n_503) );
AND2x4_ASAP7_75t_L g441 ( .A(n_234), .B(n_301), .Y(n_441) );
INVx2_ASAP7_75t_L g470 ( .A(n_234), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_234), .B(n_462), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_235), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_254), .Y(n_235) );
AND2x2_ASAP7_75t_L g381 ( .A(n_236), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g402 ( .A(n_236), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g273 ( .A(n_237), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g297 ( .A(n_237), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
AND2x2_ASAP7_75t_L g368 ( .A(n_237), .B(n_260), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_237), .B(n_352), .Y(n_409) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g321 ( .A(n_238), .Y(n_321) );
AOI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_252), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_246), .B(n_251), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_242), .B(n_245), .Y(n_241) );
AOI21x1_ASAP7_75t_L g633 ( .A1(n_245), .A2(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g586 ( .A(n_247), .Y(n_586) );
INVx2_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
INVx2_ASAP7_75t_L g547 ( .A(n_250), .Y(n_547) );
INVx3_ASAP7_75t_L g287 ( .A(n_254), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_254), .B(n_327), .Y(n_332) );
AND2x2_ASAP7_75t_L g487 ( .A(n_254), .B(n_291), .Y(n_487) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_260), .Y(n_254) );
INVx1_ASAP7_75t_L g338 ( .A(n_255), .Y(n_338) );
AND2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_274), .Y(n_366) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_259), .A2(n_278), .B(n_281), .Y(n_277) );
AND2x4_ASAP7_75t_L g319 ( .A(n_260), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g329 ( .A(n_261), .B(n_293), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_261), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_261), .B(n_274), .Y(n_391) );
AND2x2_ASAP7_75t_L g397 ( .A(n_261), .B(n_321), .Y(n_397) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_266), .A2(n_279), .B(n_280), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_266), .A2(n_533), .B(n_534), .Y(n_532) );
OAI21xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B(n_288), .Y(n_269) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_270), .A2(n_431), .B(n_435), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_270), .B(n_461), .Y(n_508) );
NAND2x1_ASAP7_75t_SL g271 ( .A(n_272), .B(n_286), .Y(n_271) );
INVx1_ASAP7_75t_L g514 ( .A(n_272), .Y(n_514) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
INVx2_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
INVxp67_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
AND2x2_ASAP7_75t_L g337 ( .A(n_274), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g348 ( .A(n_274), .B(n_349), .Y(n_348) );
INVx3_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
INVx1_ASAP7_75t_L g370 ( .A(n_274), .Y(n_370) );
OR2x2_ASAP7_75t_L g403 ( .A(n_274), .B(n_338), .Y(n_403) );
INVx1_ASAP7_75t_L g474 ( .A(n_274), .Y(n_474) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B(n_285), .Y(n_275) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B(n_299), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_290), .A2(n_413), .B1(n_415), .B2(n_418), .Y(n_412) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_291), .B(n_339), .Y(n_373) );
BUFx2_ASAP7_75t_L g432 ( .A(n_291), .Y(n_432) );
INVx2_ASAP7_75t_L g382 ( .A(n_292), .Y(n_382) );
OR2x2_ASAP7_75t_L g466 ( .A(n_292), .B(n_296), .Y(n_466) );
INVx1_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
INVx1_ASAP7_75t_L g347 ( .A(n_293), .Y(n_347) );
NOR2x1p5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_296), .Y(n_417) );
OR2x2_ASAP7_75t_L g501 ( .A(n_296), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g504 ( .A(n_296), .B(n_339), .Y(n_504) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_297), .Y(n_467) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_301), .B(n_361), .Y(n_423) );
AND2x2_ASAP7_75t_L g513 ( .A(n_301), .B(n_311), .Y(n_513) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g422 ( .A(n_302), .B(n_311), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g379 ( .A(n_303), .B(n_312), .Y(n_379) );
AND2x2_ASAP7_75t_L g414 ( .A(n_303), .B(n_308), .Y(n_414) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g333 ( .A(n_306), .B(n_314), .Y(n_333) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g473 ( .A(n_308), .B(n_474), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_316), .B1(n_322), .B2(n_325), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_310), .A2(n_511), .B(n_512), .C(n_514), .Y(n_510) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g361 ( .A(n_312), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g429 ( .A(n_312), .Y(n_429) );
OR2x2_ASAP7_75t_L g476 ( .A(n_313), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g331 ( .A(n_317), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g434 ( .A(n_320), .Y(n_434) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_321), .Y(n_349) );
INVx1_ASAP7_75t_L g421 ( .A(n_321), .Y(n_421) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g477 ( .A(n_324), .Y(n_477) );
AND2x2_ASAP7_75t_L g499 ( .A(n_324), .B(n_462), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_325), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g351 ( .A(n_329), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g407 ( .A(n_329), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g502 ( .A(n_329), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B1(n_334), .B2(n_341), .C(n_342), .Y(n_330) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx2_ASAP7_75t_L g424 ( .A(n_337), .Y(n_424) );
BUFx2_ASAP7_75t_L g444 ( .A(n_339), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_350), .B(n_353), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
AND2x2_ASAP7_75t_L g486 ( .A(n_345), .B(n_408), .Y(n_486) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
AND2x2_ASAP7_75t_L g482 ( .A(n_347), .B(n_352), .Y(n_482) );
INVx1_ASAP7_75t_L g365 ( .A(n_349), .Y(n_365) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B(n_371), .C(n_383), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_367), .B2(n_369), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
BUFx2_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
AND2x2_ASAP7_75t_L g492 ( .A(n_366), .B(n_434), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_367), .A2(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_378), .B2(n_380), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_374), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g446 ( .A(n_379), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g433 ( .A(n_382), .B(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_382), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_388), .B(n_390), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g460 ( .A(n_385), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g497 ( .A(n_385), .B(n_462), .Y(n_497) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
OR2x2_ASAP7_75t_L g489 ( .A(n_386), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g404 ( .A(n_389), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
OR2x2_ASAP7_75t_L g469 ( .A(n_389), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g440 ( .A(n_390), .Y(n_440) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_412), .C(n_419), .Y(n_393) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .A3(n_400), .B1(n_402), .B2(n_404), .C1(n_406), .C2(n_410), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_396), .A2(n_436), .B(n_472), .C(n_475), .Y(n_471) );
BUFx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g416 ( .A(n_397), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g453 ( .A(n_397), .Y(n_453) );
AND2x4_ASAP7_75t_L g481 ( .A(n_397), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI32xp33_ASAP7_75t_L g450 ( .A1(n_399), .A2(n_437), .A3(n_451), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_405), .B(n_458), .Y(n_457) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_423), .C(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_426), .B(n_483), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_430), .B(n_438), .C(n_463), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_431), .A2(n_506), .B(n_507), .C(n_509), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
OAI31xp33_ASAP7_75t_L g485 ( .A1(n_433), .A2(n_486), .A3(n_487), .B(n_488), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g445 ( .A(n_437), .Y(n_445) );
NAND4xp25_ASAP7_75t_SL g438 ( .A(n_439), .B(n_442), .C(n_450), .D(n_459), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AOI32xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .A3(n_445), .B1(n_446), .B2(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g494 ( .A(n_446), .Y(n_494) );
INVx1_ASAP7_75t_L g506 ( .A(n_449), .Y(n_506) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_471), .C(n_478), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B(n_468), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_472), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_495), .C(n_505), .D(n_510), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_486), .A2(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_503), .B2(n_504), .Y(n_498) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_502), .Y(n_511) );
INVxp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_515), .B(n_859), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_858), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_517), .B(n_753), .Y(n_516) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_518), .B(n_688), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_612), .C(n_661), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_552), .B(n_576), .C(n_593), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g827 ( .A(n_521), .B(n_746), .Y(n_827) );
OR2x2_ASAP7_75t_L g838 ( .A(n_521), .B(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_522), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g729 ( .A(n_522), .B(n_619), .Y(n_729) );
AND2x2_ASAP7_75t_L g850 ( .A(n_522), .B(n_660), .Y(n_850) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_537), .Y(n_522) );
INVx2_ASAP7_75t_L g680 ( .A(n_523), .Y(n_680) );
AND2x2_ASAP7_75t_L g695 ( .A(n_523), .B(n_647), .Y(n_695) );
AND2x2_ASAP7_75t_L g704 ( .A(n_523), .B(n_578), .Y(n_704) );
AND2x2_ASAP7_75t_L g773 ( .A(n_523), .B(n_659), .Y(n_773) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g744 ( .A(n_537), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g592 ( .A(n_538), .B(n_566), .Y(n_592) );
INVx2_ASAP7_75t_L g617 ( .A(n_538), .Y(n_617) );
AOI21x1_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .B(n_551), .Y(n_538) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g781 ( .A(n_552), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_565), .Y(n_553) );
INVx1_ASAP7_75t_L g801 ( .A(n_554), .Y(n_801) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g639 ( .A(n_555), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g722 ( .A(n_555), .B(n_628), .Y(n_722) );
AND2x2_ASAP7_75t_L g648 ( .A(n_565), .B(n_591), .Y(n_648) );
INVxp67_ASAP7_75t_L g797 ( .A(n_565), .Y(n_797) );
OR2x2_ASAP7_75t_L g839 ( .A(n_565), .B(n_578), .Y(n_839) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_575), .Y(n_566) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_589), .Y(n_576) );
INVx1_ASAP7_75t_L g694 ( .A(n_577), .Y(n_694) );
AND2x2_ASAP7_75t_L g848 ( .A(n_577), .B(n_744), .Y(n_848) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g620 ( .A(n_578), .Y(n_620) );
INVx4_ASAP7_75t_L g659 ( .A(n_578), .Y(n_659) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B(n_588), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
AND2x2_ASAP7_75t_L g675 ( .A(n_590), .B(n_658), .Y(n_675) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g712 ( .A(n_591), .B(n_660), .Y(n_712) );
INVx2_ASAP7_75t_L g678 ( .A(n_592), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_592), .B(n_683), .Y(n_846) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_595), .B(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g831 ( .A(n_595), .Y(n_831) );
AND2x2_ASAP7_75t_L g845 ( .A(n_595), .B(n_667), .Y(n_845) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_605), .Y(n_595) );
INVx1_ASAP7_75t_L g626 ( .A(n_596), .Y(n_626) );
AND2x2_ASAP7_75t_L g780 ( .A(n_596), .B(n_687), .Y(n_780) );
OR2x2_ASAP7_75t_L g817 ( .A(n_596), .B(n_605), .Y(n_817) );
AND2x2_ASAP7_75t_L g627 ( .A(n_605), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_605), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g687 ( .A(n_605), .Y(n_687) );
OR2x2_ASAP7_75t_L g700 ( .A(n_605), .B(n_640), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_605), .B(n_640), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_622), .B(n_644), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI31xp33_ASAP7_75t_L g690 ( .A1(n_614), .A2(n_691), .A3(n_693), .B(n_696), .Y(n_690) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
AND2x2_ASAP7_75t_L g703 ( .A(n_615), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g713 ( .A(n_616), .Y(n_713) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_616), .Y(n_719) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g647 ( .A(n_617), .Y(n_647) );
AND2x2_ASAP7_75t_L g676 ( .A(n_617), .B(n_660), .Y(n_676) );
INVx2_ASAP7_75t_L g726 ( .A(n_617), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_618), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g751 ( .A(n_619), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g800 ( .A(n_619), .B(n_801), .Y(n_800) );
AOI33xp33_ASAP7_75t_L g855 ( .A1(n_619), .A2(n_685), .A3(n_695), .B1(n_722), .B2(n_831), .B3(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g660 ( .A(n_621), .Y(n_660) );
INVx1_ASAP7_75t_L g747 ( .A(n_621), .Y(n_747) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_638), .Y(n_623) );
INVx2_ASAP7_75t_L g655 ( .A(n_624), .Y(n_655) );
AND2x2_ASAP7_75t_L g736 ( .A(n_624), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g698 ( .A(n_625), .Y(n_698) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g766 ( .A(n_626), .B(n_653), .Y(n_766) );
AND2x2_ASAP7_75t_L g716 ( .A(n_627), .B(n_710), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_627), .B(n_734), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_627), .B(n_766), .Y(n_815) );
AND2x2_ASAP7_75t_L g652 ( .A(n_628), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g671 ( .A(n_628), .B(n_666), .Y(n_671) );
INVx1_ASAP7_75t_L g686 ( .A(n_628), .Y(n_686) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g741 ( .A(n_639), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_639), .B(n_834), .Y(n_836) );
AND2x2_ASAP7_75t_L g849 ( .A(n_639), .B(n_665), .Y(n_849) );
AND2x2_ASAP7_75t_L g667 ( .A(n_640), .B(n_653), .Y(n_667) );
INVx2_ASAP7_75t_L g649 ( .A(n_641), .Y(n_649) );
AND2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g822 ( .A(n_641), .B(n_734), .Y(n_822) );
BUFx2_ASAP7_75t_L g804 ( .A(n_642), .Y(n_804) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx3_ASAP7_75t_L g666 ( .A(n_643), .Y(n_666) );
OAI32xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .A3(n_650), .B1(n_655), .B2(n_656), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g752 ( .A(n_647), .Y(n_752) );
AND2x2_ASAP7_75t_L g782 ( .A(n_647), .B(n_704), .Y(n_782) );
AND2x2_ASAP7_75t_L g724 ( .A(n_648), .B(n_725), .Y(n_724) );
AND3x2_ASAP7_75t_L g731 ( .A(n_648), .B(n_658), .C(n_726), .Y(n_731) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_651), .A2(n_673), .B1(n_682), .B2(n_684), .Y(n_681) );
OAI322xp33_ASAP7_75t_L g829 ( .A1(n_651), .A2(n_750), .A3(n_830), .B1(n_831), .B2(n_832), .C1(n_833), .C2(n_836), .Y(n_829) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g851 ( .A(n_652), .B(n_834), .Y(n_851) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_653), .Y(n_670) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_653), .Y(n_710) );
BUFx3_ASAP7_75t_L g734 ( .A(n_653), .Y(n_734) );
INVx1_ASAP7_75t_L g760 ( .A(n_653), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_653), .Y(n_764) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g718 ( .A(n_657), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g769 ( .A(n_658), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_658), .B(n_726), .Y(n_820) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2x1_ASAP7_75t_L g679 ( .A(n_659), .B(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g683 ( .A(n_659), .Y(n_683) );
AND2x2_ASAP7_75t_L g725 ( .A(n_659), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g746 ( .A(n_659), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_660), .B(n_773), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_668), .B(n_672), .C(n_681), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI31xp33_ASAP7_75t_L g823 ( .A1(n_663), .A2(n_824), .A3(n_826), .B(n_827), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
AND2x4_ASAP7_75t_L g776 ( .A(n_664), .B(n_685), .Y(n_776) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_665), .Y(n_708) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g792 ( .A(n_666), .B(n_686), .Y(n_792) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_677), .Y(n_672) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g832 ( .A(n_675), .Y(n_832) );
AND2x2_ASAP7_75t_L g692 ( .A(n_676), .B(n_683), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_677), .A2(n_762), .B1(n_765), .B2(n_767), .Y(n_761) );
OR2x6_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g819 ( .A(n_680), .Y(n_819) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g789 ( .A(n_685), .B(n_734), .Y(n_789) );
INVx2_ASAP7_75t_L g835 ( .A(n_685), .Y(n_835) );
AND2x4_ASAP7_75t_L g843 ( .A(n_685), .B(n_764), .Y(n_843) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_705), .C(n_735), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_701), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_692), .B(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x4_ASAP7_75t_L g756 ( .A(n_694), .B(n_711), .Y(n_756) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_697), .B(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g787 ( .A(n_699), .B(n_766), .Y(n_787) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_700), .Y(n_707) );
INVx1_ASAP7_75t_L g825 ( .A(n_700), .Y(n_825) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g854 ( .A(n_703), .Y(n_854) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_704), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .B(n_714), .C(n_727), .Y(n_705) );
NOR3x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .C(n_709), .Y(n_706) );
NAND2x1_ASAP7_75t_L g775 ( .A(n_709), .B(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2x1p5_ASAP7_75t_SL g711 ( .A(n_712), .B(n_713), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_720), .B2(n_723), .Y(n_714) );
INVxp67_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g808 ( .A(n_719), .Y(n_808) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g803 ( .A(n_722), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g857 ( .A(n_725), .Y(n_857) );
AOI21xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B(n_732), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g811 ( .A(n_732), .Y(n_811) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx2_ASAP7_75t_L g738 ( .A(n_734), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_734), .B(n_792), .Y(n_791) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_739), .B(n_740), .Y(n_735) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_738), .B(n_825), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_748), .B2(n_750), .Y(n_740) );
OR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g793 ( .A(n_743), .Y(n_793) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g768 ( .A(n_744), .B(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g785 ( .A(n_745), .Y(n_785) );
INVx1_ASAP7_75t_L g805 ( .A(n_746), .Y(n_805) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_754), .B(n_809), .Y(n_753) );
NAND3xp33_ASAP7_75t_SL g754 ( .A(n_755), .B(n_770), .C(n_783), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g816 ( .A(n_759), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2x1p5_ASAP7_75t_L g813 ( .A(n_768), .B(n_796), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_774), .B1(n_777), .B2(n_781), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g826 ( .A(n_776), .Y(n_826) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI21xp33_ASAP7_75t_L g798 ( .A1(n_778), .A2(n_799), .B(n_802), .Y(n_798) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_794), .B1(n_798), .B2(n_806), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B(n_788), .Y(n_784) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_793), .Y(n_788) );
INVx1_ASAP7_75t_L g853 ( .A(n_789), .Y(n_853) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g842 ( .A(n_792), .Y(n_842) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx2_ASAP7_75t_L g834 ( .A(n_804), .Y(n_834) );
INVxp67_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_828), .Y(n_809) );
AOI211xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B(n_814), .C(n_823), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_818), .C(n_821), .Y(n_814) );
OR2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_837), .C(n_852), .Y(n_828) );
OR2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_840), .B1(n_844), .B2(n_846), .C(n_847), .Y(n_837) );
NOR2xp67_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_847) );
OAI21xp33_ASAP7_75t_SL g852 ( .A1(n_853), .A2(n_854), .B(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_864), .B(n_891), .Y(n_890) );
BUFx4f_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx6_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x6_ASAP7_75t_SL g866 ( .A(n_867), .B(n_869), .Y(n_866) );
BUFx3_ASAP7_75t_L g887 ( .A(n_867), .Y(n_887) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx3_ASAP7_75t_L g896 ( .A(n_868), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_868), .B(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_879), .B(n_885), .Y(n_872) );
NAND2xp5_ASAP7_75t_R g873 ( .A(n_874), .B(n_877), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_875), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g898 ( .A(n_877), .Y(n_898) );
OAI21x1_ASAP7_75t_L g897 ( .A1(n_879), .A2(n_898), .B(n_899), .Y(n_897) );
AND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_884), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B(n_892), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_897), .B(n_901), .Y(n_892) );
CKINVDCx11_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx12f_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
BUFx10_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
endmodule