module fake_netlist_6_4505_n_78 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_78);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_78;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_27;
wire n_38;
wire n_61;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

AND2x6_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_16),
.B1(n_9),
.B2(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_7),
.B(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp67_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_25),
.B(n_31),
.C(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_46),
.Y(n_48)
);

AO31x2_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_33),
.A3(n_25),
.B(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_24),
.B(n_22),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_22),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_34),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_29),
.B(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_34),
.B1(n_29),
.B2(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

OR2x6_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_49),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_61),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_60),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_58),
.B(n_46),
.C(n_40),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_66),
.C(n_67),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_66),
.B(n_57),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_70),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI22x1_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_35),
.B1(n_29),
.B2(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_21),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);


endmodule