module fake_jpeg_7699_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_24),
.B1(n_28),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_70),
.B1(n_25),
.B2(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_24),
.B1(n_33),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_41),
.B1(n_30),
.B2(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_24),
.B1(n_33),
.B2(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_40),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_90),
.B(n_30),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_31),
.B1(n_25),
.B2(n_29),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_77),
.B(n_17),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_25),
.B1(n_23),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_41),
.B1(n_29),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_98),
.B1(n_51),
.B2(n_63),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_85),
.B1(n_83),
.B2(n_18),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_40),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_46),
.B1(n_45),
.B2(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_103),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_16),
.Y(n_147)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_117),
.B1(n_119),
.B2(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_47),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_116),
.C(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_121),
.B1(n_51),
.B2(n_91),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_19),
.B(n_18),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_47),
.C(n_39),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_19),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_18),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_72),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_82),
.A3(n_86),
.B1(n_45),
.B2(n_46),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_135),
.B(n_138),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_56),
.B(n_39),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_126),
.B1(n_110),
.B2(n_117),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_118),
.Y(n_163)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_45),
.A3(n_46),
.B1(n_39),
.B2(n_43),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_39),
.B1(n_53),
.B2(n_64),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_141),
.B1(n_143),
.B2(n_150),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_56),
.B1(n_81),
.B2(n_89),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_147),
.B(n_149),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_96),
.B1(n_92),
.B2(n_72),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_46),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_111),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_84),
.B1(n_45),
.B2(n_60),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_104),
.B1(n_119),
.B2(n_110),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_43),
.B(n_66),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_19),
.B1(n_32),
.B2(n_17),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_43),
.C(n_21),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_109),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_32),
.B1(n_17),
.B2(n_8),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_174),
.B(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_161),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_160),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_132),
.Y(n_161)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_74),
.B1(n_20),
.B2(n_27),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_140),
.C(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_121),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_112),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_126),
.A3(n_104),
.B1(n_107),
.B2(n_102),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_184),
.B1(n_128),
.B2(n_21),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_120),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_123),
.B(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_176),
.Y(n_197)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_124),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_136),
.A3(n_151),
.B1(n_142),
.B2(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_43),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_149),
.B1(n_155),
.B2(n_147),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_147),
.B1(n_153),
.B2(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_187),
.B(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_140),
.B1(n_117),
.B2(n_128),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_194),
.C(n_201),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_175),
.B1(n_178),
.B2(n_168),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_128),
.B1(n_60),
.B2(n_74),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_34),
.B1(n_26),
.B2(n_27),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_171),
.B1(n_166),
.B2(n_165),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_43),
.C(n_66),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_213),
.B1(n_177),
.B2(n_164),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_209),
.B1(n_174),
.B2(n_176),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_169),
.C(n_183),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_210),
.C(n_184),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_0),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_27),
.C(n_21),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_233),
.C(n_236),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_228),
.B(n_234),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_167),
.B(n_181),
.C(n_20),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_231),
.B(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_195),
.B(n_22),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_167),
.C(n_27),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_34),
.B1(n_26),
.B2(n_27),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_10),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_34),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_201),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_247),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_190),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_236),
.C(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_208),
.C(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_189),
.C(n_193),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_189),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_260),
.C(n_238),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_254),
.B(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_267),
.B(n_262),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_225),
.B(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_223),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_273),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_214),
.B1(n_196),
.B2(n_187),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_228),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_276),
.C(n_241),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_239),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_185),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_277),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_186),
.B1(n_216),
.B2(n_234),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_279),
.B1(n_246),
.B2(n_261),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_228),
.C(n_237),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_280),
.C(n_259),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_248),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_287),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_247),
.C(n_252),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_291),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_6),
.B(n_11),
.Y(n_305)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_292),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_240),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_295),
.C(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_253),
.C(n_21),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_21),
.C(n_8),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_34),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_276),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_7),
.C(n_11),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_278),
.B1(n_263),
.B2(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_268),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_279),
.B1(n_7),
.B2(n_8),
.Y(n_301)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_1),
.C(n_2),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_308),
.C(n_6),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_286),
.C(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_6),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_1),
.C(n_2),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_1),
.B(n_2),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_7),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_9),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_316),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_310),
.A2(n_300),
.B1(n_298),
.B2(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_311),
.B(n_312),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_322),
.A2(n_307),
.B(n_12),
.Y(n_327)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_325),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

OAI211xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_326),
.B(n_320),
.C(n_307),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_320),
.B(n_3),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_331),
.A3(n_328),
.B1(n_329),
.B2(n_4),
.C(n_3),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_3),
.B(n_4),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_3),
.B(n_4),
.Y(n_337)
);


endmodule