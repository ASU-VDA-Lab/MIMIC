module fake_jpeg_13434_n_448 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_48),
.B(n_55),
.Y(n_131)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_54),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_8),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_66),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_11),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_22),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_85),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_11),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_35),
.Y(n_115)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_91),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_35),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_22),
.C(n_20),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_94),
.B(n_38),
.C(n_37),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_22),
.B1(n_30),
.B2(n_46),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_92),
.B1(n_91),
.B2(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_39),
.B1(n_45),
.B2(n_36),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_132),
.B1(n_27),
.B2(n_1),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_122),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_109),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_85),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_30),
.B1(n_45),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_122),
.A2(n_128),
.B1(n_141),
.B2(n_41),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_33),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_42),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_57),
.A2(n_39),
.B1(n_45),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_76),
.B1(n_50),
.B2(n_67),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_144),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_63),
.A2(n_68),
.B1(n_70),
.B2(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_46),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_34),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_151),
.B(n_162),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

OR2x4_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_31),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_153),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_174),
.Y(n_197)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_163),
.B(n_166),
.Y(n_228)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_41),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_58),
.B1(n_53),
.B2(n_54),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g231 ( 
.A1(n_167),
.A2(n_136),
.B1(n_98),
.B2(n_101),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_168),
.B(n_172),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_179),
.C(n_137),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_97),
.B(n_40),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_100),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_176),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_27),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_10),
.C(n_9),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_10),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_9),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_99),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_185),
.B1(n_187),
.B2(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_117),
.B(n_138),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_191),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_4),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_114),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_178),
.B1(n_171),
.B2(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_105),
.B(n_6),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_96),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_217),
.B1(n_221),
.B2(n_190),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_189),
.B1(n_153),
.B2(n_154),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_154),
.A2(n_128),
.B1(n_141),
.B2(n_101),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_145),
.B(n_136),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_238),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_SL g273 ( 
.A1(n_231),
.A2(n_239),
.B(n_221),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_98),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_154),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_149),
.B(n_134),
.Y(n_238)
);

XNOR2x2_ASAP7_75t_SL g239 ( 
.A(n_151),
.B(n_111),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_192),
.C(n_170),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_134),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_152),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_241),
.A2(n_254),
.B1(n_281),
.B2(n_199),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_244),
.B(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_271),
.C(n_201),
.Y(n_282)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_248),
.B(n_250),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_185),
.B(n_183),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_250),
.A2(n_216),
.B(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_148),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_167),
.B1(n_195),
.B2(n_135),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_152),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_256),
.B(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_233),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_261),
.A2(n_262),
.B(n_252),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_212),
.A2(n_146),
.B(n_158),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_196),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_147),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_161),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_267),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_268),
.B(n_272),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_212),
.A2(n_111),
.B1(n_135),
.B2(n_123),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_273),
.B1(n_226),
.B2(n_199),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_157),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_270),
.B(n_274),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_6),
.C(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_222),
.B(n_225),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_200),
.B(n_214),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_207),
.B(n_202),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_208),
.B(n_203),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_269),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_202),
.A2(n_231),
.B1(n_219),
.B2(n_205),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_297),
.C(n_308),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_253),
.B(n_231),
.CI(n_226),
.CON(n_284),
.SN(n_284)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_312),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_286),
.A2(n_296),
.B1(n_310),
.B2(n_267),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_289),
.A2(n_295),
.B(n_303),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_201),
.B1(n_205),
.B2(n_209),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_300),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_291),
.B(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_241),
.A2(n_248),
.B1(n_281),
.B2(n_254),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_203),
.C(n_235),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_216),
.B1(n_235),
.B2(n_206),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_243),
.C(n_244),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_262),
.A2(n_247),
.B1(n_251),
.B2(n_257),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_314),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_316),
.B(n_263),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_246),
.B(n_276),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_272),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_333),
.C(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_326),
.B1(n_329),
.B2(n_334),
.Y(n_348)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_268),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_328),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_249),
.B1(n_260),
.B2(n_259),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_294),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_286),
.A2(n_259),
.B1(n_312),
.B2(n_310),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_300),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_292),
.B1(n_284),
.B2(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_292),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_283),
.B(n_317),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_338),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_316),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_301),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_302),
.C(n_305),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_299),
.Y(n_347)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_284),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_345),
.Y(n_368)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_366),
.C(n_339),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_295),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_358),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_352),
.Y(n_377)
);

NAND2x1p5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_289),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_290),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_313),
.B1(n_285),
.B2(n_304),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_360),
.A2(n_367),
.B1(n_370),
.B2(n_346),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_313),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_320),
.A2(n_285),
.B1(n_304),
.B2(n_311),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_311),
.B1(n_337),
.B2(n_324),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_366),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_345),
.B1(n_325),
.B2(n_322),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_372),
.A2(n_375),
.B1(n_370),
.B2(n_378),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_350),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_373),
.B(n_355),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_335),
.B1(n_343),
.B2(n_321),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_334),
.C(n_329),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_379),
.Y(n_394)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_319),
.C(n_342),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_382),
.A2(n_377),
.B(n_352),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_327),
.C(n_331),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_336),
.C(n_344),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_367),
.C(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_335),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_395),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_403),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_376),
.B(n_351),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_406),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_356),
.B(n_372),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_356),
.B(n_393),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_407),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_404),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_412),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_399),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_385),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_402),
.B(n_374),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_416),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_381),
.Y(n_415)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_383),
.C(n_371),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_398),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_417),
.A2(n_361),
.B1(n_362),
.B2(n_369),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_405),
.B(n_392),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_419),
.A2(n_426),
.B(n_420),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_420),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_395),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_424),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_423),
.B(n_400),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_376),
.C(n_394),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_394),
.B(n_396),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_414),
.Y(n_429)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_429),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_408),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_434),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_408),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_425),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_435),
.B(n_428),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_436),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_418),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_421),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_442),
.B(n_432),
.Y(n_443)
);

AOI211xp5_ASAP7_75t_L g445 ( 
.A1(n_443),
.A2(n_444),
.B(n_433),
.C(n_386),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_439),
.C(n_433),
.Y(n_444)
);

BUFx24_ASAP7_75t_SL g446 ( 
.A(n_445),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_447),
.A2(n_380),
.B(n_397),
.Y(n_448)
);


endmodule