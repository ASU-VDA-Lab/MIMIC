module fake_jpeg_31574_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_0),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_67),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_68),
.Y(n_90)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_19),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_92),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx11_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_68),
.B1(n_63),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_103),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_61),
.B(n_52),
.C(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_51),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_75),
.B1(n_66),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_95),
.B1(n_96),
.B2(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_53),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_121),
.B1(n_122),
.B2(n_32),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_21),
.C(n_47),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_126),
.C(n_16),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_125),
.Y(n_140)
);

OAI21x1_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_3),
.B(n_5),
.Y(n_119)
);

BUFx12f_ASAP7_75t_SL g135 ( 
.A(n_119),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_20),
.B1(n_44),
.B2(n_43),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_130),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_108),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_22),
.C(n_39),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_17),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_129),
.B(n_131),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NAND4xp25_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.D(n_144),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_141),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_10),
.C(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_139),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_13),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_14),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_49),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_120),
.A3(n_128),
.B1(n_123),
.B2(n_37),
.C1(n_38),
.C2(n_36),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_136),
.B1(n_135),
.B2(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.C(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_146),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_146),
.C(n_151),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_152),
.B(n_147),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_147),
.B(n_117),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_114),
.Y(n_160)
);


endmodule