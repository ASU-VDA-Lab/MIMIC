module real_jpeg_23598_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_80),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_41),
.B(n_88),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_1),
.A2(n_103),
.B1(n_194),
.B2(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_36),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_27),
.B1(n_36),
.B2(n_73),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_70),
.B1(n_78),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_27),
.B1(n_36),
.B2(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_83),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_83),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_27),
.B1(n_36),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_27),
.B1(n_36),
.B2(n_95),
.Y(n_124)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_27),
.B1(n_36),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_26),
.B1(n_64),
.B2(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_64),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_214)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_19),
.B(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_84),
.C(n_101),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_20),
.A2(n_21),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_22),
.B(n_54),
.C(n_68),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_23),
.A2(n_37),
.B1(n_38),
.B2(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_23),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_27),
.A2(n_36),
.B1(n_57),
.B2(n_61),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_27),
.B(n_34),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_30),
.A2(n_31),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_33),
.A2(n_34),
.B(n_70),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_34),
.A2(n_59),
.B(n_90),
.C(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_34),
.B(n_91),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_34),
.B(n_44),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_36),
.A2(n_57),
.A3(n_59),
.B1(n_212),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_39),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_39),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_40),
.A2(n_41),
.B1(n_88),
.B2(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_40),
.B(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_43),
.Y(n_153)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_46),
.A2(n_128),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_63),
.B(n_65),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_63),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_55),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_55),
.A2(n_99),
.B1(n_100),
.B2(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_56),
.A2(n_122),
.B1(n_149),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_59),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_58),
.B(n_61),
.Y(n_219)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_66),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_74),
.B1(n_80),
.B2(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_76),
.B1(n_82),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_84),
.B(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_96),
.C(n_98),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_98),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_93),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_86),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_86),
.A2(n_167),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_86),
.A2(n_175),
.B1(n_176),
.B2(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_111),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_91),
.A2(n_133),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_92),
.B(n_175),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_110),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_103),
.A2(n_129),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_103),
.A2(n_184),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_103),
.A2(n_105),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_114),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_126),
.CI(n_135),
.CON(n_114),
.SN(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_133),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_157),
.B(n_247),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_154),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_140),
.B(n_154),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_141),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_147),
.B(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_150),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_241),
.B(n_246),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_225),
.B(n_240),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_205),
.B(n_224),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_180),
.B(n_204),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_170),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_162),
.B(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_177),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_177),
.C(n_178),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B(n_203),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_188),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_197),
.B(n_202),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_217),
.B1(n_222),
.B2(n_223),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_216),
.C(n_222),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_220),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_235),
.C(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule