module fake_jpeg_18505_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_58),
.B1(n_36),
.B2(n_19),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_24),
.B2(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_45),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_42),
.B1(n_38),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_97),
.B1(n_85),
.B2(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_20),
.B1(n_37),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_75),
.A2(n_78),
.B1(n_87),
.B2(n_89),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_37),
.B1(n_42),
.B2(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_47),
.Y(n_111)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_80),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_24),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_22),
.B(n_19),
.C(n_35),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_29),
.B(n_32),
.C(n_31),
.Y(n_116)
);

AOI22x1_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_48),
.B1(n_41),
.B2(n_39),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_96),
.B1(n_102),
.B2(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_30),
.B1(n_21),
.B2(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_94),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_98),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_30),
.B1(n_36),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_95),
.B1(n_101),
.B2(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_22),
.B1(n_35),
.B2(n_19),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_36),
.B1(n_22),
.B2(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_32),
.B1(n_29),
.B2(n_17),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_32),
.B1(n_29),
.B2(n_17),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_111),
.B1(n_124),
.B2(n_23),
.Y(n_160)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_77),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_85),
.B1(n_94),
.B2(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_120),
.B1(n_132),
.B2(n_90),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_133),
.B1(n_83),
.B2(n_88),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_34),
.C(n_46),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_86),
.Y(n_150)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_25),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_131),
.B(n_134),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_47),
.B1(n_46),
.B2(n_23),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_68),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_10),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_160),
.B(n_108),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_154),
.B1(n_157),
.B2(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_84),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_148),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_144),
.B1(n_111),
.B2(n_115),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_68),
.B1(n_74),
.B2(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_91),
.B(n_71),
.C(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_70),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_156),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_73),
.B1(n_76),
.B2(n_23),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_34),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_76),
.B1(n_23),
.B2(n_17),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_103),
.B(n_16),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_119),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_122),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_168),
.B(n_177),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_186),
.B1(n_172),
.B2(n_168),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_181),
.B1(n_188),
.B2(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_123),
.C(n_116),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_116),
.B(n_111),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_189),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_118),
.B1(n_103),
.B2(n_123),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_131),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_113),
.C(n_126),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_137),
.C(n_145),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_154),
.B1(n_146),
.B2(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_107),
.B1(n_132),
.B2(n_113),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_126),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_142),
.B(n_115),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_126),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_136),
.B(n_138),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_172),
.B(n_173),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_213),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_204),
.C(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_210),
.B1(n_217),
.B2(n_182),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_141),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_147),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_135),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_208),
.B(n_211),
.Y(n_243)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_146),
.B1(n_144),
.B2(n_153),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_165),
.B(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_161),
.B(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_125),
.B1(n_162),
.B2(n_133),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_1),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_184),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_138),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_119),
.C(n_129),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_176),
.B1(n_164),
.B2(n_188),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_163),
.A2(n_121),
.B(n_122),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_228),
.B1(n_233),
.B2(n_240),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_164),
.B1(n_180),
.B2(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_170),
.B1(n_193),
.B2(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_171),
.B1(n_119),
.B2(n_183),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_197),
.A2(n_114),
.B1(n_106),
.B2(n_121),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_114),
.C(n_106),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_0),
.B(n_1),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_250),
.B(n_213),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_121),
.B1(n_3),
.B2(n_4),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_3),
.B(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_15),
.B(n_14),
.Y(n_251)
);

AOI21x1_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_250),
.B(n_247),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_263),
.B(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_207),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_266),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_198),
.B(n_199),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_238),
.B1(n_239),
.B2(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_198),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_236),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_204),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_203),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_231),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_271),
.B(n_272),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_195),
.B(n_201),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_217),
.B(n_222),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_245),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_275),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_234),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_233),
.B1(n_244),
.B2(n_246),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_290),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_257),
.B1(n_253),
.B2(n_256),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_230),
.B1(n_229),
.B2(n_235),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_237),
.C(n_230),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_229),
.C(n_235),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_206),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_226),
.C(n_248),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_258),
.A2(n_226),
.B1(n_255),
.B2(n_216),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_225),
.C(n_265),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_249),
.B(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_261),
.CI(n_265),
.CON(n_294),
.SN(n_294)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_218),
.B(n_241),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_299),
.B1(n_306),
.B2(n_11),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_225),
.B(n_252),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_14),
.C(n_13),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_304),
.C(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_13),
.C(n_12),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_287),
.C(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_13),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_273),
.C(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_273),
.C(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.C(n_304),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_294),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_296),
.C(n_300),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_294),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_312),
.B(n_302),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_299),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_301),
.B1(n_317),
.B2(n_300),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_309),
.B(n_303),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_330),
.C(n_323),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_315),
.C(n_318),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_334),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_329),
.B1(n_321),
.B2(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_328),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_331),
.B(n_336),
.Y(n_340)
);

AOI332xp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_337),
.A3(n_11),
.B1(n_5),
.B2(n_6),
.B3(n_3),
.C1(n_8),
.C2(n_9),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_4),
.B(n_5),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_7),
.B(n_9),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_9),
.Y(n_345)
);


endmodule