module real_jpeg_33857_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_705, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_705;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_703;
wire n_110;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_586;
wire n_120;
wire n_155;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_699;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_694;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_0),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_0),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_2),
.A2(n_194),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_2),
.A2(n_194),
.B1(n_392),
.B2(n_396),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_2),
.A2(n_194),
.B1(n_499),
.B2(n_502),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_3),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_3),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_3),
.A2(n_288),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_3),
.A2(n_288),
.B1(n_469),
.B2(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_3),
.A2(n_288),
.B1(n_559),
.B2(n_562),
.Y(n_558)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_4),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_132),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_4),
.A2(n_132),
.B1(n_234),
.B2(n_239),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_4),
.A2(n_132),
.B1(n_384),
.B2(n_386),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_5),
.A2(n_72),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_5),
.A2(n_293),
.B1(n_438),
.B2(n_442),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_5),
.A2(n_293),
.B1(n_530),
.B2(n_533),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_5),
.A2(n_293),
.B1(n_630),
.B2(n_632),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_75),
.B1(n_119),
.B2(n_124),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_75),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_6),
.A2(n_75),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_8),
.B(n_140),
.Y(n_415)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_8),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_8),
.B(n_67),
.Y(n_504)
);

OAI32xp33_ASAP7_75t_L g537 ( 
.A1(n_8),
.A2(n_538),
.A3(n_541),
.B1(n_543),
.B2(n_548),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_8),
.A2(n_465),
.B1(n_580),
.B2(n_583),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_L g611 ( 
.A1(n_8),
.A2(n_251),
.B(n_612),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_11),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_12),
.A2(n_139),
.B1(n_223),
.B2(n_226),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_12),
.A2(n_139),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_12),
.A2(n_139),
.B1(n_426),
.B2(n_429),
.Y(n_425)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_14),
.B(n_212),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_15),
.Y(n_123)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_16),
.A2(n_374),
.B1(n_375),
.B2(n_378),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_16),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_16),
.A2(n_374),
.B1(n_479),
.B2(n_485),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_16),
.A2(n_374),
.B1(n_586),
.B2(n_588),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_16),
.A2(n_374),
.B1(n_600),
.B2(n_604),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_17),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_18),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_18),
.A2(n_64),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_18),
.A2(n_64),
.B1(n_244),
.B2(n_248),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_214),
.B1(n_694),
.B2(n_699),
.C(n_700),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_181),
.Y(n_20)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_21),
.A2(n_22),
.B1(n_701),
.B2(n_702),
.C(n_703),
.Y(n_700)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_22),
.B(n_695),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_180),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_84),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_24),
.B(n_84),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_54),
.B1(n_65),
.B2(n_68),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_26),
.A2(n_66),
.B1(n_129),
.B2(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_26),
.A2(n_55),
.B1(n_66),
.B2(n_129),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_26),
.A2(n_66),
.B1(n_135),
.B2(n_193),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_27),
.B(n_292),
.Y(n_291)
);

NAND2x1_ASAP7_75t_SL g318 ( 
.A(n_27),
.B(n_286),
.Y(n_318)
);

AO22x1_ASAP7_75t_L g372 ( 
.A1(n_27),
.A2(n_67),
.B1(n_292),
.B2(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_27),
.B(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_29),
.Y(n_197)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_33),
.Y(n_411)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_34),
.Y(n_421)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_35),
.Y(n_196)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_36),
.Y(n_296)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_37),
.Y(n_141)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_46),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_51),
.Y(n_418)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_53),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_53),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_59),
.Y(n_414)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_59),
.Y(n_464)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_64),
.A2(n_306),
.B(n_310),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_64),
.B(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_67),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_67),
.B(n_193),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_67),
.B(n_373),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_74),
.Y(n_379)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_81),
.Y(n_377)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_177),
.C(n_179),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_85),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_127),
.C(n_142),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_87),
.B1(n_142),
.B2(n_143),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_86),
.A2(n_199),
.B(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_87),
.B(n_199),
.C(n_211),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_87),
.B(n_200),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_116),
.B(n_118),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_88),
.A2(n_116),
.B1(n_118),
.B2(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_88),
.A2(n_468),
.B1(n_474),
.B2(n_475),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_88),
.B(n_662),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_88),
.A2(n_116),
.B1(n_468),
.B2(n_672),
.Y(n_671)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_89),
.A2(n_222),
.B1(n_232),
.B2(n_233),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_89),
.A2(n_232),
.B1(n_233),
.B2(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_89),
.A2(n_222),
.B1(n_232),
.B2(n_391),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_SL g528 ( 
.A1(n_89),
.A2(n_529),
.B(n_535),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_89),
.A2(n_232),
.B1(n_529),
.B2(n_585),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_104),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

OAI22x1_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_98),
.B2(n_101),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_92),
.Y(n_606)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_97),
.Y(n_647)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_99),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_101),
.Y(n_563)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_103),
.Y(n_561)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_103),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_105),
.Y(n_542)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_106),
.Y(n_473)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_112),
.Y(n_241)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_112),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_112),
.Y(n_534)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_116),
.B(n_468),
.Y(n_535)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_117),
.B(n_465),
.Y(n_597)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_123),
.Y(n_238)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_123),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_123),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_138),
.Y(n_290)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_152),
.B1(n_168),
.B2(n_169),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_152),
.B1(n_201),
.B2(n_209),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_148),
.Y(n_282)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_148),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_149),
.Y(n_170)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_168),
.B(n_169),
.Y(n_178)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_152),
.A2(n_168),
.B1(n_201),
.B2(n_278),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_152),
.A2(n_209),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_152),
.B(n_510),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_156),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_161),
.B1(n_163),
.B2(n_167),
.Y(n_160)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_161),
.Y(n_442)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_168),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_168),
.B(n_363),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_168),
.B(n_478),
.Y(n_507)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_175),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_176),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_176),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_212),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_183),
.B(n_696),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_184),
.B(n_187),
.Y(n_698)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.C(n_198),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_189),
.B(n_211),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_192),
.B(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_198),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22x1_ASAP7_75t_L g361 ( 
.A1(n_210),
.A2(n_268),
.B1(n_269),
.B2(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_210),
.B(n_465),
.Y(n_673)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_212),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_212),
.B(n_698),
.Y(n_702)
);

INVxp33_ASAP7_75t_SL g699 ( 
.A(n_214),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_344),
.B(n_688),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_336),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_329),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_218),
.B(n_329),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_R g218 ( 
.A(n_219),
.B(n_297),
.C(n_323),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_219),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_267),
.C(n_283),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_220),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_242),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_221),
.B(n_242),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_225),
.Y(n_396)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_230),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_231),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g653 ( 
.A(n_231),
.Y(n_653)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_232),
.Y(n_474)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx4f_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_251),
.B1(n_258),
.B2(n_265),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_243),
.A2(n_251),
.B1(n_382),
.B2(n_387),
.Y(n_381)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_246),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_247),
.Y(n_385)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_247),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

OAI22x1_ASAP7_75t_L g493 ( 
.A1(n_251),
.A2(n_425),
.B1(n_494),
.B2(n_498),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_251),
.A2(n_612),
.B(n_629),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_259),
.B(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_252),
.A2(n_259),
.B(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_252),
.A2(n_266),
.B1(n_383),
.B2(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_252),
.B(n_558),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_252),
.A2(n_388),
.B1(n_627),
.B2(n_628),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

BUFx4f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_257),
.Y(n_609)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_263),
.Y(n_386)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_263),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_264),
.Y(n_428)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_264),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_264),
.Y(n_503)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_267),
.A2(n_283),
.B1(n_284),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_276),
.B2(n_277),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_268),
.A2(n_437),
.B(n_443),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_268),
.A2(n_443),
.B(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

BUFx4f_ASAP7_75t_L g409 ( 
.A(n_282),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_285),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_324),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_314),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_299),
.A2(n_320),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_300),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_301),
.Y(n_556)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_319),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g587 ( 
.A(n_309),
.Y(n_587)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_318),
.B(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_322),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_322),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_327),
.B(n_328),
.Y(n_324)
);

NAND2x1_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_327),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_342),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_336),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_337),
.B(n_339),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B(n_343),
.Y(n_339)
);

NAND2x1_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_518),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_444),
.B(n_514),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_347),
.B(n_685),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_350),
.B(n_397),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g516 ( 
.A(n_348),
.B(n_350),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_348),
.B(n_350),
.Y(n_517)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.C(n_358),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_359),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_371),
.C(n_380),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_372),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_362),
.Y(n_510)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_367),
.Y(n_550)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_403),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_390),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_381),
.B(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_389),
.Y(n_620)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_398),
.B(n_400),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.C(n_405),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_401),
.A2(n_402),
.B1(n_404),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_404),
.Y(n_449)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_432),
.C(n_435),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_SL g451 ( 
.A(n_406),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_422),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_407),
.A2(n_408),
.B1(n_422),
.B2(n_423),
.Y(n_511)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI32xp33_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.A3(n_412),
.B1(n_415),
.B2(n_416),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_430),
.Y(n_634)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_432),
.A2(n_433),
.B1(n_436),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_450),
.C(n_487),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_446),
.A2(n_686),
.B(n_687),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_450),
.Y(n_686)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.C(n_456),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_451),
.B(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_457),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_467),
.C(n_476),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_458),
.B(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_465),
.B(n_466),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_544),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_465),
.B(n_620),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_465),
.B(n_650),
.Y(n_649)
);

OAI21xp33_ASAP7_75t_SL g662 ( 
.A1(n_465),
.A2(n_649),
.B(n_663),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_476),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_471),
.Y(n_592)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_512),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_488),
.B(n_512),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.C(n_511),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_489),
.B(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_492),
.A2(n_511),
.B1(n_566),
.B2(n_567),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_504),
.B1(n_505),
.B2(n_508),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_504),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_504),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_493),
.A2(n_504),
.B1(n_505),
.B2(n_508),
.Y(n_568)
);

INVx3_ASAP7_75t_SL g494 ( 
.A(n_495),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_498),
.A2(n_556),
.B(n_557),
.Y(n_555)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_509),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B(n_517),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_684),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_569),
.B(n_682),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_564),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_522),
.B(n_683),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_527),
.C(n_536),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_524),
.B(n_572),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_527),
.A2(n_528),
.B1(n_536),
.B2(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_531),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_532),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_555),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_537),
.B(n_555),
.Y(n_576)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_551),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_557),
.A2(n_599),
.B(n_607),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_613),
.Y(n_612)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_564),
.Y(n_683)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_570),
.A2(n_593),
.B(n_681),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_571),
.B(n_574),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_571),
.B(n_574),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_577),
.C(n_584),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_667),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_584),
.Y(n_667)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_585),
.Y(n_672)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

OAI321xp33_ASAP7_75t_L g593 ( 
.A1(n_594),
.A2(n_665),
.A3(n_674),
.B1(n_679),
.B2(n_680),
.C(n_705),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_595),
.A2(n_625),
.B(n_664),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_596),
.A2(n_610),
.B(n_624),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_598),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_597),
.B(n_598),
.Y(n_624)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

BUFx2_ASAP7_75t_SL g602 ( 
.A(n_603),
.Y(n_602)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_611),
.B(n_618),
.Y(n_610)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_619),
.B(n_621),
.Y(n_618)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_635),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_626),
.B(n_635),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_636),
.B(n_660),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_660),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_637),
.A2(n_648),
.B1(n_654),
.B2(n_659),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_638),
.B(n_642),
.Y(n_637)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_638),
.Y(n_659)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx6_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_655),
.B(n_657),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_656),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_666),
.B(n_668),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_668),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_669),
.B(n_670),
.C(n_673),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_669),
.B(n_677),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_670),
.A2(n_671),
.B1(n_673),
.B2(n_678),
.Y(n_677)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_671),
.Y(n_670)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_673),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_675),
.B(n_676),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_SL g679 ( 
.A(n_675),
.B(n_676),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_689),
.A2(n_690),
.B(n_692),
.Y(n_688)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_691),
.Y(n_690)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_693),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_696),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_697),
.B(n_698),
.Y(n_696)
);


endmodule