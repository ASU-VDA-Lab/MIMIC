module fake_jpeg_19807_n_186 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_30),
.B1(n_20),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_50),
.B1(n_33),
.B2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_20),
.B1(n_29),
.B2(n_19),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_22),
.B1(n_29),
.B2(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_15),
.B1(n_56),
.B2(n_28),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_35),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_78),
.C(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_27),
.B1(n_24),
.B2(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_24),
.B1(n_17),
.B2(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_81),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_41),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_40),
.Y(n_80)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_34),
.CI(n_41),
.CON(n_81),
.SN(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_1),
.B1(n_5),
.B2(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_9),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_11),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_58),
.Y(n_112)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_88),
.B1(n_67),
.B2(n_86),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_58),
.B(n_4),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_103),
.B(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_80),
.C(n_63),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_102),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_101),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_1),
.C(n_5),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_70),
.B1(n_82),
.B2(n_81),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_69),
.B(n_68),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_123),
.C(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_81),
.B1(n_74),
.B2(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_95),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_138),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_143),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_92),
.B1(n_108),
.B2(n_100),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_115),
.B(n_117),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_91),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_154),
.C(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_155),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_124),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_129),
.C(n_131),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_134),
.C(n_126),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_154),
.C(n_137),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_147),
.C(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_99),
.C(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_163),
.B1(n_157),
.B2(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_160),
.C(n_122),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.C(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_166),
.B(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_172),
.C(n_94),
.Y(n_179)
);

AOI21x1_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_175),
.B(n_136),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_145),
.B1(n_95),
.B2(n_119),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_181),
.B(n_94),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_101),
.Y(n_186)
);


endmodule