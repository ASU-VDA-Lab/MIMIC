module real_jpeg_11096_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_344, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_344;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_1),
.A2(n_64),
.B1(n_67),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_155),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_155),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_155),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_2),
.A2(n_3),
.B(n_31),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_47),
.B(n_59),
.C(n_86),
.D(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_45),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_3),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_107),
.B(n_109),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_3),
.A2(n_30),
.B(n_41),
.C(n_143),
.D(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_30),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_34),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_124),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_4),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_4),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_4),
.A2(n_127),
.B(n_153),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_9),
.A2(n_22),
.B1(n_64),
.B2(n_67),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_9),
.A2(n_22),
.B1(n_46),
.B2(n_47),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_10),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_11),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_64),
.B1(n_67),
.B2(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_101),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_101),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_12),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_89),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_89),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_89),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_54),
.B1(n_64),
.B2(n_67),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_54),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_15),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_106),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_106),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_106),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_16),
.A2(n_33),
.B1(n_64),
.B2(n_67),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_336),
.B(n_339),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_75),
.B(n_335),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_20),
.B(n_35),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_20),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_20),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_32),
.B2(n_34),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_21),
.A2(n_25),
.B1(n_34),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_23),
.A2(n_27),
.B(n_124),
.C(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_25),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_25),
.B(n_205),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_338)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_26),
.A2(n_29),
.B1(n_219),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_204),
.B(n_242),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_285),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_29),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_29),
.A2(n_220),
.B(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_34),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_70),
.C(n_72),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_36),
.A2(n_37),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_57),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_38),
.A2(n_39),
.B1(n_57),
.B2(n_310),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_40),
.A2(n_49),
.B1(n_164),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_40),
.A2(n_199),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_45),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_41),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_41),
.A2(n_45),
.B1(n_239),
.B2(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_41),
.A2(n_45),
.B1(n_257),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_43),
.B(n_46),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_44),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_47),
.A2(n_143),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_49),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_49),
.A2(n_165),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_51),
.A2(n_52),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_57),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_57),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_58),
.A2(n_68),
.B1(n_100),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_58),
.A2(n_141),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_58),
.A2(n_68),
.B1(n_196),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_58),
.A2(n_68),
.B1(n_214),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_58),
.A2(n_68),
.B1(n_233),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_59),
.A2(n_63),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_67),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_64),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_108),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_67),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_68),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_68),
.A2(n_102),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_69),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_70),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_328),
.B(n_334),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_301),
.A3(n_321),
.B1(n_326),
.B2(n_327),
.C(n_343),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_249),
.A3(n_289),
.B1(n_295),
.B2(n_300),
.C(n_344),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_207),
.C(n_246),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_179),
.B(n_206),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_158),
.B(n_178),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_135),
.B(n_157),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_112),
.B(n_134),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_84),
.B(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_99),
.C(n_104),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_109),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_108),
.B1(n_154),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_107),
.A2(n_108),
.B1(n_169),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_107),
.A2(n_108),
.B1(n_189),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_107),
.A2(n_108),
.B1(n_212),
.B2(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_107),
.A2(n_108),
.B(n_231),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_116),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_124),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_121),
.B(n_133),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_128),
.B(n_132),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_148),
.B2(n_156),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_147),
.C(n_156),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_174),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_175),
.C(n_176),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_173),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_170),
.C(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_181),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_193),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_192),
.C(n_193),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_188),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_208),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_226),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_209),
.B(n_226),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_215),
.CI(n_216),
.CON(n_209),
.SN(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_244),
.B2(n_245),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_234),
.C(n_245),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_240),
.C(n_243),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_267),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_250),
.B(n_267),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_260),
.C(n_266),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_251),
.A2(n_252),
.B1(n_260),
.B2(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_262),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_261),
.A2(n_280),
.B(n_284),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_263),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_287),
.B2(n_288),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_278),
.B2(n_279),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_279),
.C(n_288),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_275),
.B(n_277),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_277),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_277),
.A2(n_303),
.B1(n_312),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_286),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_282),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_314),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_312),
.C(n_313),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_305),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_310),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_316),
.C(n_320),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_333),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_330),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_338),
.B(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);


endmodule