module real_jpeg_32991_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_1),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_1),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_1),
.B(n_286),
.Y(n_285)
);

NAND2x1_ASAP7_75t_L g396 ( 
.A(n_1),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_1),
.B(n_402),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_1),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_1),
.B(n_528),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_2),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_2),
.B(n_36),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_2),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_2),
.B(n_389),
.Y(n_388)
);

AND2x4_ASAP7_75t_SL g499 ( 
.A(n_2),
.B(n_113),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_2),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_2),
.B(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_2),
.B(n_581),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_4),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_4),
.B(n_362),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_4),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_4),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_5),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_5),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_5),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_367),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_R g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_11),
.B1(n_53),
.B2(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_6),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_6),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_6),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_6),
.B(n_297),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_7),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_7),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_9),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_11),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_11),
.B(n_152),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_11),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_11),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_11),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_11),
.B(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_11),
.B(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_11),
.B(n_520),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_12),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g407 ( 
.A(n_12),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_12),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_12),
.B(n_393),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_12),
.B(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_12),
.B(n_536),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_12),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_21),
.B(n_24),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_14),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_87),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_14),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_14),
.Y(n_228)
);

NAND2x1_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_15),
.B(n_36),
.Y(n_154)
);

AND2x4_ASAP7_75t_SL g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_15),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_15),
.B(n_47),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_15),
.B(n_427),
.Y(n_426)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_16),
.B(n_607),
.C(n_617),
.Y(n_616)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_17),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_17),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_18),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_18),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_18),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_18),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_18),
.B(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_19),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_457),
.B(n_566),
.C(n_602),
.D(n_616),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_351),
.B(n_454),
.Y(n_27)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_252),
.B(n_348),
.Y(n_28)
);

AO21x2_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_155),
.B(n_251),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_136),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_31),
.B(n_136),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_83),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_32),
.B(n_346),
.C(n_347),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_50),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_33),
.B(n_51),
.C(n_68),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.C(n_45),
.Y(n_33)
);

XNOR2x2_ASAP7_75t_L g140 ( 
.A(n_34),
.B(n_141),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_35),
.B(n_37),
.Y(n_143)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_40),
.Y(n_215)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_41),
.B(n_46),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_44),
.Y(n_280)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_49),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_49),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_49),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_68),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_63),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_56),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_57),
.Y(n_323)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_62),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_63),
.B(n_307),
.C(n_313),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_63),
.A2(n_313),
.B1(n_314),
.B2(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_63),
.Y(n_339)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_67),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_67),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_69),
.B(n_77),
.C(n_82),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_71),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_71),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_75),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_80),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_120),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_84),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_100),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_85),
.B(n_101),
.C(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_86),
.B(n_94),
.C(n_98),
.Y(n_314)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_89),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_90),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_90),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_90),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_90),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_109),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_120),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_135),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_135),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_131),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_127),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_130),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_131),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_138),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_140),
.B(n_142),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.C(n_149),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_148),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_154),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_245),
.B(n_250),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_195),
.B(n_244),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_187),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_158),
.B(n_187),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_173),
.B(n_186),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_170),
.C(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_181),
.Y(n_412)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_193),
.C(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_208),
.B(n_243),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_206),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.C(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_199),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_223),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_204),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_225),
.B(n_240),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_233),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_232),
.Y(n_409)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_248),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_333),
.B(n_341),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_253),
.B(n_333),
.C(n_349),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_282),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_254),
.B(n_283),
.C(n_451),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_270),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2x2_ASAP7_75t_L g334 ( 
.A(n_256),
.B(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_259),
.A2(n_270),
.B1(n_271),
.B2(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_259),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_263),
.C(n_268),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_264),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2x2_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_305),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_293),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_294),
.C(n_295),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_288),
.C(n_291),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_285),
.B(n_288),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_285),
.B(n_288),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_290),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g430 ( 
.A1(n_291),
.A2(n_360),
.B(n_366),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_296),
.B(n_301),
.C(n_303),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx4f_ASAP7_75t_SL g520 ( 
.A(n_298),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_303),
.B(n_410),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_303),
.B(n_411),
.C(n_420),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_305),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_315),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_306),
.Y(n_444)
);

XOR2x2_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.C(n_311),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_312),
.Y(n_491)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_324),
.B1(n_325),
.B2(n_332),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_316),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_316),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_319),
.C(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_325),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.B(n_330),
.C(n_331),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_329),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.C(n_340),
.Y(n_333)
);

AOI221xp5_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.C(n_345),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_334),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_342),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_340),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_342),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_449),
.Y(n_351)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_352),
.A2(n_455),
.B(n_456),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_438),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_353),
.B(n_438),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_371),
.Y(n_353)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_354),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.C(n_369),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_355),
.A2(n_356),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_357),
.B(n_369),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_365),
.B2(n_366),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_360),
.A2(n_361),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_360),
.B(n_366),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_366),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_360),
.B(n_426),
.C(n_428),
.Y(n_488)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g538 ( 
.A(n_364),
.Y(n_538)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_367),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_368),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_413),
.B1(n_436),
.B2(n_437),
.Y(n_371)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_372),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_399),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_387),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g500 ( 
.A(n_374),
.B(n_387),
.C(n_400),
.Y(n_500)
);

XNOR2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_378),
.Y(n_484)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.C(n_396),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_396),
.Y(n_416)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_405),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_401),
.B(n_406),
.C(n_410),
.Y(n_481)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_406),
.A2(n_407),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_406),
.B(n_473),
.C(n_475),
.Y(n_548)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_422),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_417),
.C(n_418),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_417),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_448),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_431),
.B(n_432),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B(n_435),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.C(n_447),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_447),
.Y(n_453)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.C(n_446),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_452),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NOR3x1_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_505),
.C(n_561),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_501),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_462),
.B(n_501),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_469),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_465),
.B(n_470),
.C(n_486),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.C(n_468),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_486),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_480),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_481),
.C(n_482),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_473),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_473),
.A2(n_474),
.B1(n_524),
.B2(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_474),
.B(n_522),
.C(n_527),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.C(n_485),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_500),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_488),
.B(n_500),
.C(n_555),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_493),
.C(n_499),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_498),
.B2(n_499),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_497),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_499),
.Y(n_498)
);

MAJx2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.C(n_504),
.Y(n_501)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_553),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g596 ( 
.A(n_507),
.B(n_553),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_544),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_517),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_509),
.B(n_544),
.C(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.C(n_514),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_547),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_514),
.Y(n_547)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_517),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_532),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_521),
.B1(n_530),
.B2(n_531),
.Y(n_518)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_519),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_519),
.B(n_572),
.C(n_573),
.Y(n_571)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_521),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_522),
.A2(n_523),
.B1(n_534),
.B2(n_535),
.Y(n_533)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_531),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_539),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_577),
.C(n_578),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_534),
.A2(n_587),
.B1(n_588),
.B2(n_594),
.Y(n_586)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_548),
.C(n_549),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_560),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_548),
.B(n_550),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_556),
.C(n_558),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_554),
.B(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_557),
.B(n_559),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_562),
.A2(n_600),
.B(n_601),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_564),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_SL g566 ( 
.A(n_567),
.B(n_596),
.C(n_597),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_570),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_568),
.B(n_570),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_574),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_571),
.A2(n_595),
.B(n_613),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_595),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_575),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_579),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_579),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_586),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_588),
.C(n_594),
.Y(n_611)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_587),
.A2(n_588),
.B1(n_606),
.B2(n_607),
.Y(n_605)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_589),
.B(n_593),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_593),
.B(n_608),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_598),
.B(n_599),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_614),
.Y(n_602)
);

AOI221xp5_ASAP7_75t_L g603 ( 
.A1(n_604),
.A2(n_605),
.B1(n_610),
.B2(n_611),
.C(n_612),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_604),
.A2(n_605),
.B1(n_610),
.B2(n_611),
.Y(n_618)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_607),
.Y(n_606)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_612),
.B(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);


endmodule