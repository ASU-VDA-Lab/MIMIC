module fake_jpeg_12092_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_46),
.B(n_66),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_18),
.A2(n_5),
.B(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_50),
.B(n_0),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_21),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_21),
.B(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_39),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_0),
.Y(n_77)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_8),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_8),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_33),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_77),
.B(n_90),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_30),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_29),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_79),
.A2(n_87),
.B(n_81),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_82),
.B(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_85),
.B(n_89),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_108),
.B1(n_115),
.B2(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_37),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_107),
.Y(n_128)
);

OR2x4_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_29),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_121),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_1),
.B1(n_13),
.B2(n_88),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_22),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_112),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_48),
.A2(n_34),
.B1(n_25),
.B2(n_36),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_125),
.B1(n_93),
.B2(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_36),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_30),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_124),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_58),
.A2(n_25),
.B1(n_22),
.B2(n_35),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_30),
.B1(n_20),
.B2(n_33),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_13),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_30),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_65),
.B(n_11),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_73),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_141),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_114),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_20),
.B1(n_56),
.B2(n_1),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_1),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_20),
.B1(n_3),
.B2(n_10),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_143),
.A2(n_145),
.B1(n_156),
.B2(n_149),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_155),
.B1(n_138),
.B2(n_139),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_148),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_147),
.B(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_114),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_79),
.A2(n_103),
.B(n_88),
.C(n_124),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_163),
.B1(n_102),
.B2(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_75),
.B(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_84),
.A2(n_125),
.B1(n_100),
.B2(n_93),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_104),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_166),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_164),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_81),
.A2(n_91),
.B1(n_87),
.B2(n_97),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_136),
.B1(n_148),
.B2(n_127),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_74),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_97),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_97),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_175),
.A2(n_176),
.B(n_197),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_102),
.B(n_84),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_181),
.A2(n_206),
.B1(n_186),
.B2(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_195),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_126),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_196),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_192),
.A2(n_199),
.B1(n_205),
.B2(n_183),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_147),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_129),
.B1(n_128),
.B2(n_168),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_161),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_162),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_204),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_152),
.B(n_132),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_137),
.B1(n_153),
.B2(n_151),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_133),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_155),
.A3(n_157),
.B1(n_166),
.B2(n_160),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_174),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_142),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_215),
.B(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_224),
.B1(n_228),
.B2(n_205),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_223),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_133),
.C(n_170),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_225),
.C(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_233),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_175),
.B(n_179),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_230),
.B(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_142),
.B1(n_176),
.B2(n_203),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_188),
.C(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_184),
.B1(n_180),
.B2(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_184),
.B(n_210),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_185),
.B(n_174),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_232),
.A2(n_222),
.B1(n_226),
.B2(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_187),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_238),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_178),
.B(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_241),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_177),
.B(n_186),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_241),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_205),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_225),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_262),
.C(n_245),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_253),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_221),
.B(n_235),
.C(n_236),
.D(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_219),
.B1(n_212),
.B2(n_211),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_256),
.B1(n_267),
.B2(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_213),
.B1(n_217),
.B2(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_214),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_261),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_230),
.C(n_224),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_238),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_233),
.B(n_214),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_283),
.B1(n_259),
.B2(n_250),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_276),
.B(n_255),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_281),
.C(n_289),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_287),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_264),
.B(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_245),
.C(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_285),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_248),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_268),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_250),
.C(n_243),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_258),
.A3(n_244),
.B1(n_255),
.B2(n_253),
.C1(n_268),
.C2(n_243),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_297),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_252),
.C(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_293),
.C(n_300),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_259),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_298),
.B(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_275),
.B(n_289),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_301),
.B(n_278),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_281),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_319),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_275),
.C(n_298),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_317),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_287),
.B(n_272),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_309),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_272),
.B(n_274),
.C(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_286),
.B(n_269),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_315),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_277),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_279),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_295),
.B1(n_303),
.B2(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_325),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_290),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_316),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_307),
.B(n_319),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_313),
.B(n_314),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_335),
.C(n_322),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_334),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_314),
.B1(n_290),
.B2(n_288),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_329),
.C(n_306),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_329),
.B(n_323),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_339),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

AOI321xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_341),
.A3(n_322),
.B1(n_326),
.B2(n_282),
.C(n_321),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_326),
.Y(n_345)
);


endmodule