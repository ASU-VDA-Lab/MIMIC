module real_aes_2149_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g100 ( .A1(n_0), .A2(n_56), .B1(n_90), .B2(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g183 ( .A(n_1), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_2), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g265 ( .A(n_3), .Y(n_265) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_4), .A2(n_15), .B1(n_90), .B2(n_98), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_5), .Y(n_281) );
INVx2_ASAP7_75t_L g198 ( .A(n_6), .Y(n_198) );
INVx1_ASAP7_75t_L g244 ( .A(n_7), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_7), .A2(n_80), .B1(n_160), .B2(n_244), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g83 ( .A1(n_8), .A2(n_36), .B1(n_76), .B2(n_84), .C1(n_102), .C2(n_106), .Y(n_83) );
INVx1_ASAP7_75t_L g241 ( .A(n_9), .Y(n_241) );
INVx1_ASAP7_75t_SL g216 ( .A(n_10), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_11), .B(n_219), .Y(n_325) );
AOI33xp33_ASAP7_75t_L g293 ( .A1(n_12), .A2(n_38), .A3(n_204), .B1(n_212), .B2(n_294), .B3(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g274 ( .A(n_13), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_14), .A2(n_80), .B1(n_160), .B2(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_14), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g175 ( .A1(n_15), .A2(n_56), .B1(n_58), .B2(n_176), .C(n_178), .Y(n_175) );
OR2x2_ASAP7_75t_L g199 ( .A(n_16), .B(n_69), .Y(n_199) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_16), .A2(n_69), .B(n_198), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_17), .A2(n_35), .B1(n_153), .B2(n_156), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_18), .B(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_20), .A2(n_67), .B1(n_112), .B2(n_117), .Y(n_111) );
INVx1_ASAP7_75t_SL g91 ( .A(n_21), .Y(n_91) );
INVx1_ASAP7_75t_L g185 ( .A(n_22), .Y(n_185) );
AND2x2_ASAP7_75t_L g207 ( .A(n_22), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g225 ( .A(n_22), .B(n_183), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_23), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_24), .B(n_202), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_25), .A2(n_44), .B1(n_140), .B2(n_143), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_26), .A2(n_228), .B1(n_234), .B2(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_27), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_28), .B(n_219), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_29), .A2(n_37), .B1(n_122), .B2(n_127), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_30), .A2(n_162), .B1(n_170), .B2(n_171), .Y(n_161) );
INVx1_ASAP7_75t_L g170 ( .A(n_30), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_31), .B(n_262), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_32), .B(n_219), .Y(n_266) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_33), .A2(n_58), .B1(n_90), .B2(n_94), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_34), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_39), .B(n_219), .Y(n_305) );
INVx1_ASAP7_75t_L g205 ( .A(n_40), .Y(n_205) );
INVx1_ASAP7_75t_L g221 ( .A(n_40), .Y(n_221) );
AND2x2_ASAP7_75t_L g306 ( .A(n_41), .B(n_196), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_42), .A2(n_48), .B1(n_146), .B2(n_148), .Y(n_145) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_43), .A2(n_60), .B1(n_202), .B2(n_210), .C(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_45), .B(n_202), .Y(n_257) );
INVx1_ASAP7_75t_L g92 ( .A(n_46), .Y(n_92) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_47), .A2(n_54), .B1(n_132), .B2(n_136), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_49), .B(n_228), .Y(n_283) );
AOI21xp5_ASAP7_75t_SL g253 ( .A1(n_50), .A2(n_210), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_51), .A2(n_80), .B1(n_159), .B2(n_160), .Y(n_79) );
INVx1_ASAP7_75t_L g159 ( .A(n_51), .Y(n_159) );
INVx1_ASAP7_75t_L g237 ( .A(n_52), .Y(n_237) );
INVx1_ASAP7_75t_L g304 ( .A(n_53), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_55), .A2(n_210), .B(n_303), .Y(n_302) );
INVxp33_ASAP7_75t_L g180 ( .A(n_56), .Y(n_180) );
INVx1_ASAP7_75t_L g208 ( .A(n_57), .Y(n_208) );
INVx1_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVxp67_ASAP7_75t_L g179 ( .A(n_58), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_59), .B(n_202), .Y(n_296) );
INVx1_ASAP7_75t_L g167 ( .A(n_60), .Y(n_167) );
AND2x2_ASAP7_75t_L g226 ( .A(n_61), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g238 ( .A(n_62), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_63), .A2(n_210), .B(n_215), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_64), .A2(n_210), .B(n_288), .C(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_65), .B(n_227), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_66), .A2(n_210), .B1(n_291), .B2(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g164 ( .A(n_68), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_70), .A2(n_167), .B1(n_168), .B2(n_169), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_70), .Y(n_168) );
INVx1_ASAP7_75t_L g255 ( .A(n_71), .Y(n_255) );
AND2x2_ASAP7_75t_L g297 ( .A(n_72), .B(n_227), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_73), .A2(n_272), .B(n_273), .C(n_275), .Y(n_271) );
BUFx2_ASAP7_75t_SL g177 ( .A(n_74), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_75), .B(n_219), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_172), .B1(n_186), .B2(n_547), .C(n_550), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_161), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_80), .Y(n_160) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_130), .Y(n_81) );
NAND3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_111), .C(n_121), .Y(n_82) );
INVx4_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
INVx6_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x4_ASAP7_75t_L g104 ( .A(n_87), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_88), .Y(n_116) );
AND2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
OAI22x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_90), .Y(n_101) );
AND2x2_ASAP7_75t_L g109 ( .A(n_93), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
BUFx2_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
AND2x4_ASAP7_75t_L g134 ( .A(n_95), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g142 ( .A(n_95), .B(n_109), .Y(n_142) );
AND2x4_ASAP7_75t_L g155 ( .A(n_95), .B(n_119), .Y(n_155) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x4_ASAP7_75t_L g108 ( .A(n_97), .B(n_99), .Y(n_108) );
AND2x2_ASAP7_75t_L g115 ( .A(n_97), .B(n_100), .Y(n_115) );
INVx1_ASAP7_75t_L g126 ( .A(n_97), .Y(n_126) );
INVxp67_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g129 ( .A(n_100), .B(n_126), .Y(n_129) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g118 ( .A(n_108), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g144 ( .A(n_108), .B(n_135), .Y(n_144) );
AND2x2_ASAP7_75t_L g147 ( .A(n_109), .B(n_129), .Y(n_147) );
AND2x4_ASAP7_75t_L g135 ( .A(n_110), .B(n_120), .Y(n_135) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x4_ASAP7_75t_L g150 ( .A(n_115), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g158 ( .A(n_115), .B(n_135), .Y(n_158) );
BUFx5_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g128 ( .A(n_119), .B(n_129), .Y(n_128) );
BUFx4f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g138 ( .A(n_129), .B(n_135), .Y(n_138) );
NAND4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_139), .C(n_145), .D(n_152), .Y(n_130) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
INVx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx8_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx5_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_162), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_SL g169 ( .A(n_167), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
AND3x1_ASAP7_75t_SL g174 ( .A(n_175), .B(n_181), .C(n_184), .Y(n_174) );
INVxp67_ASAP7_75t_L g557 ( .A(n_175), .Y(n_557) );
CKINVDCx8_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_181), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_181), .A2(n_320), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g203 ( .A(n_182), .B(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_SL g562 ( .A(n_182), .B(n_184), .Y(n_562) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g214 ( .A(n_183), .B(n_205), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_184), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2x1p5_ASAP7_75t_L g211 ( .A(n_185), .B(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR3x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_412), .C(n_483), .Y(n_188) );
NAND3x1_ASAP7_75t_SL g189 ( .A(n_190), .B(n_339), .C(n_361), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_329), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_258), .B1(n_307), .B2(n_311), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_192), .A2(n_515), .B1(n_516), .B2(n_518), .Y(n_514) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_230), .Y(n_192) );
AND2x2_ASAP7_75t_L g330 ( .A(n_193), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_193), .B(n_377), .Y(n_396) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g314 ( .A(n_194), .Y(n_314) );
AND2x2_ASAP7_75t_L g364 ( .A(n_194), .B(n_232), .Y(n_364) );
INVx1_ASAP7_75t_L g403 ( .A(n_194), .Y(n_403) );
OR2x2_ASAP7_75t_L g440 ( .A(n_194), .B(n_250), .Y(n_440) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_194), .Y(n_452) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_194), .Y(n_476) );
AND2x2_ASAP7_75t_L g533 ( .A(n_194), .B(n_360), .Y(n_533) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_200), .B(n_226), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AND2x4_ASAP7_75t_L g234 ( .A(n_198), .B(n_199), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_209), .Y(n_200) );
INVx1_ASAP7_75t_L g284 ( .A(n_202), .Y(n_284) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_206), .Y(n_202) );
INVx1_ASAP7_75t_L g320 ( .A(n_203), .Y(n_320) );
OR2x6_ASAP7_75t_L g217 ( .A(n_204), .B(n_213), .Y(n_217) );
INVxp33_ASAP7_75t_L g294 ( .A(n_204), .Y(n_294) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x4_ASAP7_75t_L g246 ( .A(n_205), .B(n_222), .Y(n_246) );
INVx1_ASAP7_75t_L g321 ( .A(n_206), .Y(n_321) );
BUFx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x6_ASAP7_75t_L g549 ( .A(n_207), .B(n_214), .Y(n_549) );
INVx2_ASAP7_75t_L g213 ( .A(n_208), .Y(n_213) );
AND2x6_ASAP7_75t_L g243 ( .A(n_208), .B(n_220), .Y(n_243) );
INVxp67_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
INVx1_ASAP7_75t_L g295 ( .A(n_212), .Y(n_295) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_217), .B(n_218), .C(n_224), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_217), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_224), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_217), .A2(n_224), .B(n_265), .C(n_266), .Y(n_264) );
INVxp67_ASAP7_75t_L g272 ( .A(n_217), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_217), .A2(n_224), .B(n_304), .C(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g327 ( .A(n_217), .Y(n_327) );
INVx1_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_224), .B(n_234), .Y(n_247) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_224), .A2(n_325), .B(n_326), .Y(n_324) );
INVx5_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_225), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_227), .A2(n_271), .B1(n_276), .B2(n_277), .Y(n_270) );
INVx3_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_228), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx4f_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
NOR2x1_ASAP7_75t_L g230 ( .A(n_231), .B(n_248), .Y(n_230) );
INVx1_ASAP7_75t_L g408 ( .A(n_231), .Y(n_408) );
AND2x2_ASAP7_75t_L g434 ( .A(n_231), .B(n_250), .Y(n_434) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_231), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g331 ( .A(n_232), .B(n_317), .Y(n_331) );
INVx3_ASAP7_75t_L g360 ( .A(n_232), .Y(n_360) );
NOR2x1_ASAP7_75t_SL g479 ( .A(n_232), .B(n_250), .Y(n_479) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_234), .A2(n_253), .B(n_257), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .B(n_247), .Y(n_235) );
OAI222xp33_ASAP7_75t_L g550 ( .A1(n_237), .A2(n_551), .B1(n_552), .B2(n_558), .C1(n_560), .C2(n_563), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_239), .B(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B1(n_244), .B2(n_245), .Y(n_240) );
INVxp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_248), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g358 ( .A(n_249), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_250), .Y(n_373) );
AND2x2_ASAP7_75t_L g445 ( .A(n_250), .B(n_317), .Y(n_445) );
AND2x4_ASAP7_75t_L g462 ( .A(n_250), .B(n_406), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_250), .B(n_404), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_250), .B(n_313), .Y(n_538) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_258), .A2(n_355), .B1(n_426), .B2(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_285), .Y(n_258) );
INVx2_ASAP7_75t_L g428 ( .A(n_259), .Y(n_428) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
BUFx3_ASAP7_75t_L g418 ( .A(n_260), .Y(n_418) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_261), .B(n_287), .Y(n_310) );
INVx2_ASAP7_75t_L g334 ( .A(n_261), .Y(n_334) );
INVx1_ASAP7_75t_L g346 ( .A(n_261), .Y(n_346) );
AND2x4_ASAP7_75t_L g353 ( .A(n_261), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g370 ( .A(n_261), .B(n_269), .Y(n_370) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_261), .Y(n_384) );
INVxp67_ASAP7_75t_L g392 ( .A(n_261), .Y(n_392) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_267), .Y(n_261) );
INVx2_ASAP7_75t_SL g288 ( .A(n_262), .Y(n_288) );
AND2x2_ASAP7_75t_L g421 ( .A(n_268), .B(n_337), .Y(n_421) );
AND2x2_ASAP7_75t_L g437 ( .A(n_268), .B(n_338), .Y(n_437) );
NOR2xp67_ASAP7_75t_L g524 ( .A(n_268), .B(n_337), .Y(n_524) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g333 ( .A(n_269), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g344 ( .A(n_269), .Y(n_344) );
INVx1_ASAP7_75t_L g357 ( .A(n_269), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_269), .B(n_299), .Y(n_394) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_278), .Y(n_269) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_277), .A2(n_300), .B(n_306), .Y(n_299) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_277), .A2(n_300), .B(n_306), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B1(n_283), .B2(n_284), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g517 ( .A(n_285), .Y(n_517) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_298), .Y(n_285) );
AND2x2_ASAP7_75t_L g391 ( .A(n_286), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g420 ( .A(n_286), .Y(n_420) );
AND2x2_ASAP7_75t_L g522 ( .A(n_286), .B(n_337), .Y(n_522) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_287), .B(n_299), .Y(n_382) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_297), .Y(n_287) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_289), .B(n_297), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_290), .B(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g308 ( .A(n_298), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_298), .B(n_418), .Y(n_497) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_299), .Y(n_411) );
AND2x2_ASAP7_75t_L g438 ( .A(n_299), .B(n_384), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g352 ( .A(n_308), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
AND2x2_ASAP7_75t_L g456 ( .A(n_308), .B(n_333), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_308), .B(n_476), .Y(n_481) );
AND2x2_ASAP7_75t_L g491 ( .A(n_308), .B(n_370), .Y(n_491) );
OR2x2_ASAP7_75t_L g528 ( .A(n_308), .B(n_428), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_309), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g488 ( .A(n_309), .B(n_344), .Y(n_488) );
AND2x2_ASAP7_75t_L g504 ( .A(n_309), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g498 ( .A(n_310), .B(n_394), .Y(n_498) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
INVx1_ASAP7_75t_L g380 ( .A(n_312), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_312), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g478 ( .A(n_312), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_312), .B(n_359), .Y(n_503) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_313), .Y(n_350) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_314), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_348), .B1(n_366), .B2(n_369), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_315), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g482 ( .A(n_315), .Y(n_482) );
AND2x4_ASAP7_75t_SL g315 ( .A(n_316), .B(n_328), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g359 ( .A(n_317), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g379 ( .A(n_317), .Y(n_379) );
INVx1_ASAP7_75t_L g406 ( .A(n_317), .Y(n_406) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_323), .Y(n_317) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .C(n_322), .Y(n_319) );
INVxp67_ASAP7_75t_L g565 ( .A(n_321), .Y(n_565) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_328), .Y(n_348) );
AND2x4_ASAP7_75t_L g405 ( .A(n_328), .B(n_406), .Y(n_405) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_328), .B(n_435), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g430 ( .A(n_330), .B(n_373), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_330), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g388 ( .A(n_331), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_332), .A2(n_442), .B1(n_446), .B2(n_449), .Y(n_441) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
AND2x2_ASAP7_75t_L g409 ( .A(n_333), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g448 ( .A(n_333), .Y(n_448) );
NAND2x1_ASAP7_75t_SL g473 ( .A(n_333), .B(n_342), .Y(n_473) );
AND2x2_ASAP7_75t_L g369 ( .A(n_335), .B(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_337), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g342 ( .A(n_338), .Y(n_342) );
INVx2_ASAP7_75t_L g354 ( .A(n_338), .Y(n_354) );
AOI21xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_347), .B(n_351), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_342), .B(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_343), .A2(n_432), .B1(n_436), .B2(n_439), .Y(n_431) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
BUFx2_ASAP7_75t_L g536 ( .A(n_344), .Y(n_536) );
INVx1_ASAP7_75t_SL g543 ( .A(n_344), .Y(n_543) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_345), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B(n_358), .Y(n_351) );
AND2x2_ASAP7_75t_L g355 ( .A(n_353), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g397 ( .A(n_353), .B(n_393), .Y(n_397) );
AND2x2_ASAP7_75t_L g512 ( .A(n_353), .B(n_410), .Y(n_512) );
AND2x2_ASAP7_75t_L g515 ( .A(n_353), .B(n_421), .Y(n_515) );
AND2x4_ASAP7_75t_L g523 ( .A(n_353), .B(n_524), .Y(n_523) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_355), .A2(n_478), .B(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g505 ( .A(n_357), .Y(n_505) );
AND2x2_ASAP7_75t_L g521 ( .A(n_357), .B(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g435 ( .A(n_359), .Y(n_435) );
INVx1_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
AND2x2_ASAP7_75t_L g426 ( .A(n_360), .B(n_379), .Y(n_426) );
NOR2x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_385), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_371), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g372 ( .A(n_364), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_SL g525 ( .A(n_364), .B(n_377), .Y(n_525) );
AND2x2_ASAP7_75t_L g546 ( .A(n_364), .B(n_462), .Y(n_546) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g472 ( .A(n_369), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_374), .B(n_381), .Y(n_371) );
OR2x6_ASAP7_75t_L g424 ( .A(n_373), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g447 ( .A(n_382), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g544 ( .A(n_382), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_383), .B(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_395), .B2(n_397), .Y(n_386) );
OR2x2_ASAP7_75t_L g458 ( .A(n_388), .B(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g464 ( .A(n_393), .Y(n_464) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_407), .B2(n_409), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
AND2x4_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_405), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g468 ( .A(n_408), .B(n_462), .Y(n_468) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_453), .Y(n_412) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_414), .B(n_427), .Y(n_413) );
AOI21xp33_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_422), .Y(n_414) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp33_ASAP7_75t_SL g492 ( .A1(n_424), .A2(n_493), .B1(n_495), .B2(n_498), .Y(n_492) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_425), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g475 ( .A(n_426), .B(n_476), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_431), .C(n_441), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVxp33_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g444 ( .A(n_435), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_436), .A2(n_456), .B1(n_457), .B2(n_460), .C(n_463), .Y(n_455) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
INVx2_ASAP7_75t_SL g494 ( .A(n_440), .Y(n_494) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2x1_ASAP7_75t_L g493 ( .A(n_444), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g490 ( .A(n_450), .Y(n_490) );
INVx1_ASAP7_75t_L g519 ( .A(n_451), .Y(n_519) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR2x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_469), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_467), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g529 ( .A(n_462), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g534 ( .A(n_462), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVxp33_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g487 ( .A(n_466), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_474), .B(n_477), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g530 ( .A(n_476), .Y(n_530) );
AND2x2_ASAP7_75t_L g518 ( .A(n_479), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_R g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_499), .C(n_526), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_486), .B(n_489), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_501), .B(n_510), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_504), .B1(n_506), .B2(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_509), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_520), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_523), .B(n_525), .Y(n_520) );
INVx1_ASAP7_75t_L g539 ( .A(n_523), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B(n_531), .C(n_540), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_535), .B1(n_537), .B2(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
endmodule