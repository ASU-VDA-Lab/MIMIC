module fake_netlist_1_9006_n_697 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_16), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_43), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_74), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_52), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_29), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_7), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_57), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_77), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_64), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_78), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_75), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_65), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_22), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_14), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_53), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_5), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_39), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_21), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_44), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_13), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_55), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_27), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_31), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_25), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_16), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_60), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_116), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_80), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_97), .B(n_0), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_88), .B(n_0), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_93), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_122), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_85), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_84), .B(n_1), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_104), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_84), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_104), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_88), .B(n_1), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_103), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_89), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_101), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_90), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_95), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_99), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_92), .B(n_2), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_92), .B(n_3), .Y(n_166) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_118), .B(n_3), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_114), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_98), .Y(n_170) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_166), .B(n_127), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_130), .B(n_123), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_130), .B(n_109), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_155), .B(n_170), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_142), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_158), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_166), .B(n_127), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_170), .B(n_112), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_128), .B(n_113), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_128), .B(n_105), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
NOR2x1_ASAP7_75t_L g198 ( .A(n_131), .B(n_102), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_168), .B(n_117), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_131), .B(n_119), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_135), .B(n_120), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_135), .B(n_120), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_161), .B(n_98), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_169), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_161), .B(n_100), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_169), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_140), .B(n_121), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_140), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_143), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_152), .B(n_100), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_166), .B(n_123), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_152), .B(n_79), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_153), .B(n_106), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_153), .B(n_111), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_156), .B(n_125), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_156), .B(n_115), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_157), .B(n_160), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_154), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_157), .B(n_108), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_159), .B(n_124), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_205), .B(n_160), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_172), .B(n_159), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_192), .Y(n_244) );
NOR2xp67_ASAP7_75t_L g245 ( .A(n_186), .B(n_163), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_231), .A2(n_137), .B(n_165), .C(n_148), .Y(n_246) );
NOR3xp33_ASAP7_75t_SL g247 ( .A(n_186), .B(n_138), .C(n_141), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_205), .B(n_167), .Y(n_249) );
NAND3xp33_ASAP7_75t_SL g250 ( .A(n_189), .B(n_132), .C(n_129), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
NOR3xp33_ASAP7_75t_SL g252 ( .A(n_199), .B(n_136), .C(n_144), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_176), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_215), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
NOR2xp33_ASAP7_75t_R g256 ( .A(n_183), .B(n_136), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_205), .B(n_164), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_210), .B(n_167), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_210), .B(n_165), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_190), .B(n_162), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_210), .B(n_164), .Y(n_263) );
NOR2xp33_ASAP7_75t_R g264 ( .A(n_178), .B(n_163), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_218), .B(n_162), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
NOR3xp33_ASAP7_75t_SL g267 ( .A(n_179), .B(n_144), .C(n_148), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_216), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_218), .B(n_162), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_228), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_184), .B(n_137), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_221), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_171), .B(n_154), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_172), .B(n_124), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_216), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_192), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_192), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_172), .B(n_91), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_219), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_202), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_172), .B(n_121), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_201), .B(n_94), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_171), .B(n_110), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_233), .A2(n_4), .B(n_5), .C(n_6), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_171), .B(n_4), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_222), .B(n_36), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_222), .B(n_6), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_192), .B(n_8), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_220), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_192), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_223), .B(n_8), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_221), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_223), .B(n_9), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_220), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_194), .B(n_9), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_180), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_226), .B(n_10), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_266), .B(n_244), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_272), .B(n_223), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_267), .B(n_252), .C(n_246), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_242), .B(n_232), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_269), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_259), .A2(n_209), .B(n_191), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_300), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_261), .Y(n_317) );
INVx3_ASAP7_75t_SL g318 ( .A(n_266), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_300), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_242), .B(n_232), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_237), .B(n_232), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
OAI21x1_ASAP7_75t_SL g324 ( .A1(n_266), .A2(n_203), .B(n_204), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_279), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_235), .B1(n_226), .B2(n_231), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_264), .B(n_180), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_300), .A2(n_226), .B1(n_235), .B2(n_198), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_261), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_261), .Y(n_330) );
NAND2xp33_ASAP7_75t_L g331 ( .A(n_262), .B(n_188), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_285), .A2(n_206), .B(n_188), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_262), .A2(n_198), .B(n_217), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_257), .B(n_235), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_285), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_292), .B(n_227), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_244), .B(n_226), .Y(n_337) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_291), .A2(n_293), .A3(n_303), .B(n_288), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_302), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_261), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_288), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_302), .A2(n_227), .B1(n_196), .B2(n_191), .Y(n_342) );
INVx8_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_298), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_276), .A2(n_195), .B1(n_206), .B2(n_211), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_263), .B(n_178), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_249), .B(n_209), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_280), .B(n_236), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_298), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_280), .B(n_211), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_305), .B(n_234), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_241), .B(n_234), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_281), .A2(n_193), .B1(n_208), .B2(n_212), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_281), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_261), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_253), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_282), .B(n_193), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_273), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_253), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_343), .B(n_282), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_294), .B(n_274), .C(n_301), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_359), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_343), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_343), .A2(n_306), .B1(n_284), .B2(n_299), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_308), .A2(n_265), .B(n_270), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_353), .B(n_250), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_336), .A2(n_275), .B1(n_278), .B2(n_249), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_339), .B(n_299), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_343), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_353), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_351), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_339), .B(n_245), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_339), .A2(n_256), .B1(n_178), .B2(n_258), .Y(n_377) );
INVx5_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_327), .Y(n_379) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_324), .B(n_253), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_325), .Y(n_381) );
OAI22xp5_ASAP7_75t_SL g382 ( .A1(n_326), .A2(n_284), .B1(n_290), .B2(n_258), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_346), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_318), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_316), .A2(n_251), .B(n_277), .Y(n_385) );
AOI21xp5_ASAP7_75t_SL g386 ( .A1(n_316), .A2(n_295), .B(n_286), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_337), .B(n_268), .Y(n_387) );
BUFx2_ASAP7_75t_SL g388 ( .A(n_337), .Y(n_388) );
NAND2xp33_ASAP7_75t_R g389 ( .A(n_350), .B(n_247), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_346), .B(n_249), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_336), .B(n_258), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_310), .A2(n_289), .B(n_304), .C(n_287), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_311), .B(n_262), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_362), .A2(n_331), .B(n_324), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_382), .A2(n_321), .B1(n_334), .B2(n_322), .C(n_342), .Y(n_395) );
BUFx4f_ASAP7_75t_SL g396 ( .A(n_371), .Y(n_396) );
INVx6_ASAP7_75t_SL g397 ( .A(n_361), .Y(n_397) );
BUFx4f_ASAP7_75t_SL g398 ( .A(n_371), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_332), .B(n_333), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_390), .A2(n_319), .B1(n_337), .B2(n_328), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_378), .A2(n_328), .B1(n_319), .B2(n_358), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_390), .A2(n_337), .B1(n_348), .B2(n_344), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_383), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_320), .B1(n_335), .B2(n_314), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_376), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_391), .A2(n_345), .B1(n_349), .B2(n_344), .C(n_352), .Y(n_408) );
AOI21x1_ASAP7_75t_L g409 ( .A1(n_380), .A2(n_349), .B(n_352), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_366), .A2(n_320), .B1(n_314), .B2(n_309), .Y(n_410) );
AO31x2_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_309), .A3(n_335), .B(n_341), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_368), .A2(n_348), .B1(n_355), .B2(n_341), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_392), .B(n_331), .C(n_197), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_378), .Y(n_414) );
AO221x2_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_10), .B1(n_11), .B2(n_12), .C(n_15), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_367), .A2(n_333), .B(n_315), .C(n_347), .Y(n_416) );
OR2x6_ASAP7_75t_L g417 ( .A(n_388), .B(n_350), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_393), .B(n_359), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_372), .B(n_338), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_338), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_373), .B(n_338), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_378), .A2(n_358), .B1(n_350), .B2(n_355), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_407), .B(n_369), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_395), .A2(n_369), .B1(n_421), .B2(n_407), .C(n_420), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_419), .B(n_338), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_396), .A2(n_378), .B1(n_389), .B2(n_375), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_394), .A2(n_385), .B(n_174), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_413), .A2(n_386), .B(n_230), .Y(n_428) );
AOI21xp33_ASAP7_75t_SL g429 ( .A1(n_414), .A2(n_389), .B(n_379), .Y(n_429) );
NOR4xp25_ASAP7_75t_SL g430 ( .A(n_415), .B(n_377), .C(n_229), .D(n_230), .Y(n_430) );
NOR2xp67_ASAP7_75t_SL g431 ( .A(n_414), .B(n_384), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_405), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_409), .A2(n_229), .B(n_271), .Y(n_433) );
AOI31xp33_ASAP7_75t_L g434 ( .A1(n_422), .A2(n_365), .A3(n_387), .B(n_307), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_417), .A2(n_361), .B1(n_364), .B2(n_375), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_415), .A2(n_375), .B1(n_364), .B2(n_361), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_419), .B(n_338), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_415), .A2(n_384), .B1(n_370), .B2(n_348), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_420), .B(n_387), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_234), .B(n_200), .C(n_187), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_415), .A2(n_370), .B1(n_330), .B2(n_329), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_418), .B(n_348), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_354), .B(n_251), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_358), .Y(n_445) );
AND2x6_ASAP7_75t_SL g446 ( .A(n_405), .B(n_358), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_417), .A2(n_307), .B1(n_318), .B2(n_268), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_400), .A2(n_360), .B1(n_357), .B2(n_312), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
NAND4xp75_ASAP7_75t_L g450 ( .A(n_418), .B(n_187), .C(n_200), .D(n_207), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
NOR2xp33_ASAP7_75t_R g452 ( .A(n_398), .B(n_318), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_402), .A2(n_238), .B1(n_357), .B2(n_323), .C(n_313), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_404), .B(n_273), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_410), .A2(n_197), .B1(n_208), .B2(n_212), .C(n_225), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_417), .A2(n_307), .B1(n_268), .B2(n_356), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_411), .B(n_213), .Y(n_457) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_408), .A2(n_207), .B1(n_213), .B2(n_225), .C1(n_296), .C2(n_283), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_404), .B(n_297), .Y(n_459) );
INVx4_ASAP7_75t_L g460 ( .A(n_446), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_439), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_439), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_445), .B(n_411), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_423), .B(n_411), .Y(n_464) );
AOI21xp5_ASAP7_75t_SL g465 ( .A1(n_434), .A2(n_417), .B(n_401), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_426), .A2(n_416), .A3(n_397), .B(n_283), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_449), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_425), .B(n_399), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_427), .Y(n_470) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_424), .A2(n_409), .B(n_399), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_399), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_437), .B(n_399), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_437), .B(n_317), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_440), .B(n_197), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_440), .B(n_197), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_457), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_457), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_435), .A2(n_397), .B1(n_317), .B2(n_329), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_443), .B(n_197), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_449), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_451), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_438), .B(n_11), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_433), .B(n_317), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_429), .B(n_17), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_433), .B(n_317), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_442), .B(n_173), .C(n_177), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_454), .B(n_18), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_454), .B(n_19), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_428), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_428), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_430), .B(n_173), .C(n_177), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_436), .B(n_19), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_428), .B(n_21), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_432), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_431), .Y(n_503) );
AOI21xp33_ASAP7_75t_SL g504 ( .A1(n_456), .A2(n_22), .B(n_23), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_441), .B(n_23), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_431), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_452), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_448), .A2(n_174), .B1(n_175), .B2(n_181), .C(n_182), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_493), .B(n_24), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_479), .B(n_455), .Y(n_513) );
OR2x6_ASAP7_75t_L g514 ( .A(n_465), .B(n_397), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_469), .B(n_24), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_469), .B(n_26), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_495), .B(n_458), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_465), .A2(n_453), .B(n_330), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_462), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_503), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_481), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_495), .B(n_296), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_473), .B(n_28), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_477), .B(n_297), .Y(n_528) );
OAI211xp5_ASAP7_75t_L g529 ( .A1(n_460), .A2(n_175), .B(n_182), .C(n_181), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_473), .B(n_34), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_482), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_478), .B(n_356), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_460), .A2(n_317), .B1(n_329), .B2(n_356), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_478), .B(n_356), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_463), .B(n_472), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_502), .B(n_35), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_463), .B(n_37), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_463), .B(n_40), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_468), .B(n_356), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_491), .B(n_329), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_500), .A2(n_360), .B1(n_357), .B2(n_312), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_492), .B(n_340), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_472), .B(n_42), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_508), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_492), .B(n_340), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_474), .B(n_45), .Y(n_549) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_503), .A2(n_329), .B(n_340), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_484), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_508), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_511), .B(n_500), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_474), .B(n_48), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_474), .B(n_49), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_460), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_506), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_511), .B(n_340), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_464), .B(n_340), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_475), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_466), .B(n_330), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_506), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_476), .B(n_330), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_476), .B(n_330), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_485), .B(n_173), .Y(n_566) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_507), .B(n_360), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_557), .B(n_488), .C(n_501), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_556), .A2(n_483), .B1(n_505), .B2(n_510), .C1(n_507), .C2(n_496), .Y(n_572) );
XNOR2xp5_ASAP7_75t_L g573 ( .A(n_547), .B(n_475), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_552), .B(n_510), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_535), .B(n_510), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_567), .B(n_490), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_514), .A2(n_471), .B1(n_480), .B2(n_487), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_567), .A2(n_504), .B(n_499), .C(n_487), .Y(n_578) );
OAI32xp33_ASAP7_75t_L g579 ( .A1(n_538), .A2(n_498), .A3(n_494), .B1(n_486), .B2(n_471), .Y(n_579) );
NOR2xp33_ASAP7_75t_R g580 ( .A(n_515), .B(n_50), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_513), .A2(n_487), .B(n_489), .Y(n_581) );
OAI31xp33_ASAP7_75t_SL g582 ( .A1(n_539), .A2(n_489), .A3(n_494), .B(n_498), .Y(n_582) );
OAI32xp33_ASAP7_75t_L g583 ( .A1(n_512), .A2(n_471), .A3(n_497), .B1(n_489), .B2(n_470), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_514), .A2(n_471), .B1(n_470), .B2(n_497), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_535), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_560), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_514), .A2(n_470), .B1(n_312), .B2(n_323), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_515), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_569), .B(n_470), .Y(n_589) );
NOR4xp25_ASAP7_75t_L g590 ( .A(n_563), .B(n_509), .C(n_470), .D(n_323), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_553), .B(n_54), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_514), .A2(n_313), .B1(n_255), .B2(n_254), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_519), .A2(n_313), .B1(n_173), .B2(n_177), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_539), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_517), .B(n_58), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_516), .B(n_59), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_544), .A2(n_173), .B1(n_177), .B2(n_254), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_561), .A2(n_255), .B(n_254), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_561), .B(n_177), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_523), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_61), .Y(n_601) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_533), .A2(n_248), .B(n_239), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_540), .B(n_62), .Y(n_603) );
OR4x1_ASAP7_75t_L g604 ( .A(n_524), .B(n_63), .C(n_67), .D(n_68), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_518), .B(n_70), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_531), .B(n_73), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
AOI32xp33_ASAP7_75t_SL g609 ( .A1(n_536), .A2(n_76), .A3(n_185), .B1(n_255), .B2(n_243), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_524), .A2(n_185), .B1(n_239), .B2(n_248), .C(n_243), .Y(n_611) );
OAI33xp33_ASAP7_75t_L g612 ( .A1(n_513), .A2(n_185), .A3(n_243), .B1(n_254), .B2(n_255), .B3(n_260), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_522), .A2(n_243), .B(n_254), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_529), .A2(n_243), .B1(n_255), .B2(n_260), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_516), .B(n_260), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_521), .B(n_537), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_542), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g618 ( .A1(n_549), .A2(n_555), .B(n_554), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_570), .B(n_568), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_594), .B(n_521), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_573), .B(n_530), .Y(n_621) );
XNOR2xp5_ASAP7_75t_L g622 ( .A(n_585), .B(n_530), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_586), .B(n_527), .Y(n_623) );
OAI321xp33_ASAP7_75t_L g624 ( .A1(n_581), .A2(n_546), .A3(n_527), .B1(n_549), .B2(n_555), .C(n_554), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_588), .B(n_551), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_575), .B(n_546), .Y(n_626) );
NOR3xp33_ASAP7_75t_SL g627 ( .A(n_618), .B(n_548), .C(n_545), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_600), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_617), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_616), .B(n_566), .Y(n_630) );
CKINVDCx20_ASAP7_75t_L g631 ( .A(n_580), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_582), .A2(n_559), .B(n_543), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_574), .B(n_562), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_618), .B(n_528), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_572), .B(n_566), .C(n_562), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_612), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_572), .A2(n_571), .B1(n_610), .B2(n_581), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_589), .B(n_541), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_606), .B(n_532), .Y(n_639) );
INVx3_ASAP7_75t_SL g640 ( .A(n_599), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_591), .B(n_528), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_605), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_582), .B(n_532), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_576), .B(n_526), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_608), .Y(n_645) );
NOR4xp25_ASAP7_75t_SL g646 ( .A(n_578), .B(n_550), .C(n_541), .D(n_534), .Y(n_646) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_598), .B(n_534), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_601), .A2(n_565), .B1(n_564), .B2(n_558), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_577), .B(n_590), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_590), .B(n_593), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_607), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_619), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_634), .A2(n_584), .B1(n_603), .B2(n_587), .Y(n_653) );
AOI211xp5_ASAP7_75t_SL g654 ( .A1(n_624), .A2(n_584), .B(n_613), .C(n_614), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_622), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_630), .Y(n_656) );
NAND2x1_ASAP7_75t_L g657 ( .A(n_627), .B(n_592), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_637), .B(n_579), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_627), .A2(n_595), .B1(n_596), .B2(n_597), .C(n_609), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_640), .B(n_615), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_628), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_629), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_636), .B(n_604), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_620), .A2(n_583), .B(n_611), .C(n_602), .Y(n_664) );
NOR3xp33_ASAP7_75t_SL g665 ( .A(n_631), .B(n_615), .C(n_620), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_625), .B(n_633), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_621), .B(n_642), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_643), .B(n_626), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_639), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_655), .A2(n_634), .B1(n_649), .B2(n_635), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_665), .A2(n_636), .B(n_632), .C(n_644), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_658), .A2(n_644), .B1(n_650), .B2(n_640), .C(n_651), .Y(n_672) );
NOR2xp33_ASAP7_75t_R g673 ( .A(n_655), .B(n_641), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_656), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_653), .A2(n_623), .B1(n_641), .B2(n_648), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_663), .A2(n_647), .B1(n_638), .B2(n_645), .Y(n_676) );
AOI211xp5_ASAP7_75t_SL g677 ( .A1(n_664), .A2(n_646), .B(n_659), .C(n_654), .Y(n_677) );
AOI21xp33_ASAP7_75t_SL g678 ( .A1(n_667), .A2(n_660), .B(n_668), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_657), .B(n_660), .C(n_667), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_652), .A2(n_669), .B(n_666), .C(n_662), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_661), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_668), .A2(n_665), .B(n_654), .C(n_663), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_660), .A2(n_620), .B(n_663), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_663), .B1(n_637), .B2(n_634), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_673), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_677), .A2(n_670), .B1(n_679), .B2(n_682), .C(n_684), .Y(n_686) );
NOR3xp33_ASAP7_75t_SL g687 ( .A(n_671), .B(n_672), .C(n_683), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_678), .Y(n_688) );
INVxp33_ASAP7_75t_SL g689 ( .A(n_673), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_685), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_689), .A2(n_686), .B1(n_688), .B2(n_687), .Y(n_691) );
NOR3xp33_ASAP7_75t_SL g692 ( .A(n_689), .B(n_671), .C(n_680), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_690), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_691), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_693), .Y(n_695) );
OAI321xp33_ASAP7_75t_L g696 ( .A1(n_695), .A2(n_694), .A3(n_692), .B1(n_676), .B2(n_675), .C(n_674), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_694), .B(n_681), .Y(n_697) );
endmodule