module real_aes_2519_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_831, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_831;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_782;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g235 ( .A(n_0), .B(n_157), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_1), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g150 ( .A(n_2), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_3), .B(n_163), .Y(n_176) );
NAND2xp33_ASAP7_75t_SL g227 ( .A(n_4), .B(n_161), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_5), .Y(n_829) );
INVx1_ASAP7_75t_L g208 ( .A(n_6), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_7), .B(n_181), .Y(n_554) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_8), .A2(n_125), .B1(n_126), .B2(n_128), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_8), .Y(n_125) );
INVx1_ASAP7_75t_L g534 ( .A(n_9), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_10), .Y(n_119) );
AND2x2_ASAP7_75t_L g174 ( .A(n_11), .B(n_167), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_12), .Y(n_501) );
INVx2_ASAP7_75t_L g168 ( .A(n_13), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_14), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_15), .B(n_28), .Y(n_730) );
INVx1_ASAP7_75t_L g562 ( .A(n_16), .Y(n_562) );
OAI22xp5_ASAP7_75t_SL g816 ( .A1(n_17), .A2(n_28), .B1(n_784), .B2(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_17), .Y(n_817) );
AOI221x1_ASAP7_75t_L g221 ( .A1(n_18), .A2(n_145), .B1(n_222), .B2(n_224), .C(n_226), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_19), .B(n_163), .Y(n_196) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g560 ( .A(n_21), .Y(n_560) );
INVx1_ASAP7_75t_SL g483 ( .A(n_22), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_23), .B(n_164), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_24), .A2(n_145), .B(n_178), .Y(n_177) );
AOI221xp5_ASAP7_75t_SL g188 ( .A1(n_25), .A2(n_41), .B1(n_145), .B2(n_163), .C(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_26), .B(n_157), .Y(n_179) );
AOI33xp33_ASAP7_75t_L g520 ( .A1(n_27), .A2(n_54), .A3(n_211), .B1(n_217), .B2(n_521), .B3(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g784 ( .A(n_28), .Y(n_784) );
INVx1_ASAP7_75t_L g494 ( .A(n_29), .Y(n_494) );
OR2x2_ASAP7_75t_L g169 ( .A(n_30), .B(n_94), .Y(n_169) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_30), .A2(n_94), .B(n_168), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_31), .B(n_153), .Y(n_200) );
INVxp67_ASAP7_75t_L g220 ( .A(n_32), .Y(n_220) );
AND2x2_ASAP7_75t_L g251 ( .A(n_33), .B(n_166), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_34), .B(n_209), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_35), .A2(n_145), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_36), .B(n_153), .Y(n_190) );
AND2x2_ASAP7_75t_L g146 ( .A(n_37), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g161 ( .A(n_37), .B(n_150), .Y(n_161) );
INVx1_ASAP7_75t_L g216 ( .A(n_37), .Y(n_216) );
OR2x6_ASAP7_75t_L g113 ( .A(n_38), .B(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_39), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_40), .B(n_209), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_42), .A2(n_181), .B1(n_225), .B2(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_43), .B(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_44), .A2(n_84), .B1(n_145), .B2(n_214), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_45), .B(n_164), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_46), .B(n_157), .Y(n_249) );
INVx1_ASAP7_75t_L g792 ( .A(n_47), .Y(n_792) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_48), .B(n_88), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_49), .B(n_201), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_50), .B(n_164), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_51), .Y(n_547) );
AND2x2_ASAP7_75t_L g238 ( .A(n_52), .B(n_166), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_53), .B(n_166), .Y(n_192) );
XOR2xp5_ASAP7_75t_L g811 ( .A(n_53), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_55), .B(n_164), .Y(n_512) );
INVx1_ASAP7_75t_L g149 ( .A(n_56), .Y(n_149) );
INVx1_ASAP7_75t_L g159 ( .A(n_56), .Y(n_159) );
AND2x2_ASAP7_75t_L g513 ( .A(n_57), .B(n_166), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_58), .A2(n_77), .B1(n_209), .B2(n_214), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_59), .B(n_209), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_60), .B(n_163), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_61), .A2(n_124), .B1(n_129), .B2(n_130), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_61), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_62), .B(n_225), .Y(n_503) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_63), .A2(n_214), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g170 ( .A(n_64), .B(n_166), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_65), .B(n_153), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_66), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_SL g203 ( .A(n_67), .B(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g557 ( .A(n_68), .Y(n_557) );
XNOR2xp5_ASAP7_75t_L g126 ( .A(n_69), .B(n_127), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_70), .A2(n_145), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g511 ( .A(n_71), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_72), .B(n_153), .Y(n_180) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_73), .B(n_201), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_74), .A2(n_214), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g147 ( .A(n_75), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_75), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_76), .B(n_209), .Y(n_523) );
AND2x2_ASAP7_75t_L g485 ( .A(n_78), .B(n_224), .Y(n_485) );
INVx1_ASAP7_75t_L g558 ( .A(n_79), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_80), .A2(n_214), .B(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_81), .A2(n_214), .B(n_284), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_82), .B(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_83), .A2(n_87), .B1(n_163), .B2(n_209), .Y(n_286) );
INVx1_ASAP7_75t_L g116 ( .A(n_85), .Y(n_116) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_86), .B(n_224), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_89), .A2(n_214), .B1(n_518), .B2(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_90), .B(n_157), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_91), .B(n_157), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_92), .B(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_93), .A2(n_145), .B(n_151), .Y(n_144) );
INVx1_ASAP7_75t_L g474 ( .A(n_95), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_96), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g524 ( .A(n_97), .B(n_224), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_98), .A2(n_492), .B(n_493), .C(n_495), .Y(n_491) );
INVxp67_ASAP7_75t_L g223 ( .A(n_99), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_100), .B(n_163), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_101), .B(n_153), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_102), .A2(n_145), .B(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_SL g790 ( .A(n_103), .Y(n_790) );
BUFx2_ASAP7_75t_L g803 ( .A(n_103), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_104), .B(n_164), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_120), .B(n_828), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_108), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_117), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_111), .B(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g785 ( .A(n_112), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_112), .B(n_797), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_113), .Y(n_797) );
OAI32xp33_ASAP7_75t_L g798 ( .A1(n_113), .A2(n_799), .A3(n_800), .B1(n_801), .B2(n_832), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_804), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_786), .B(n_798), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_131), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_123), .Y(n_827) );
INVxp33_ASAP7_75t_L g130 ( .A(n_124), .Y(n_130) );
INVx1_ASAP7_75t_L g128 ( .A(n_126), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_132), .Y(n_826) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_460), .Y(n_132) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_399), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_292), .C(n_343), .Y(n_135) );
OAI211xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_182), .B(n_239), .C(n_270), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_141), .B(n_244), .Y(n_407) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g252 ( .A(n_142), .B(n_173), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_142), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g269 ( .A(n_142), .B(n_259), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_142), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g306 ( .A(n_142), .B(n_282), .Y(n_306) );
INVx2_ASAP7_75t_L g332 ( .A(n_142), .Y(n_332) );
AND2x4_ASAP7_75t_L g341 ( .A(n_142), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g446 ( .A(n_142), .B(n_313), .Y(n_446) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_165), .B(n_170), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_162), .Y(n_143) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
BUFx3_ASAP7_75t_L g213 ( .A(n_146), .Y(n_213) );
AND2x6_ASAP7_75t_L g157 ( .A(n_147), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g218 ( .A(n_147), .Y(n_218) );
AND2x4_ASAP7_75t_L g214 ( .A(n_148), .B(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x4_ASAP7_75t_L g153 ( .A(n_149), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B(n_160), .Y(n_151) );
INVxp67_ASAP7_75t_L g563 ( .A(n_153), .Y(n_563) );
AND2x4_ASAP7_75t_L g164 ( .A(n_154), .B(n_158), .Y(n_164) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVxp67_ASAP7_75t_L g561 ( .A(n_157), .Y(n_561) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_160), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_160), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_160), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_160), .A2(n_248), .B(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_160), .A2(n_474), .B(n_475), .C(n_476), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_160), .A2(n_475), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_160), .A2(n_475), .B(n_511), .C(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g518 ( .A(n_160), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_160), .A2(n_475), .B(n_534), .C(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_160), .A2(n_550), .B(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_160), .B(n_181), .Y(n_564) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g163 ( .A(n_161), .B(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_161), .Y(n_495) );
INVx1_ASAP7_75t_L g228 ( .A(n_164), .Y(n_228) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_165), .A2(n_245), .B(n_251), .Y(n_244) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_165), .A2(n_245), .B(n_251), .Y(n_259) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_165), .A2(n_479), .B(n_485), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_166), .A2(n_188), .B(n_192), .Y(n_187) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x4_ASAP7_75t_L g181 ( .A(n_168), .B(n_169), .Y(n_181) );
AND2x2_ASAP7_75t_L g330 ( .A(n_171), .B(n_331), .Y(n_330) );
OAI32xp33_ASAP7_75t_L g413 ( .A1(n_171), .A2(n_335), .A3(n_339), .B1(n_346), .B2(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_171), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g267 ( .A(n_172), .B(n_268), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_172), .B(n_262), .C(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g366 ( .A(n_172), .B(n_269), .Y(n_366) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
INVx5_ASAP7_75t_L g291 ( .A(n_173), .Y(n_291) );
AND2x4_ASAP7_75t_L g347 ( .A(n_173), .B(n_259), .Y(n_347) );
OR2x2_ASAP7_75t_L g362 ( .A(n_173), .B(n_282), .Y(n_362) );
OR2x2_ASAP7_75t_L g388 ( .A(n_173), .B(n_244), .Y(n_388) );
AND2x2_ASAP7_75t_L g396 ( .A(n_173), .B(n_342), .Y(n_396) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_173), .B(n_341), .Y(n_421) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_181), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_181), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_181), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_181), .B(n_223), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g226 ( .A(n_181), .B(n_227), .C(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_181), .A2(n_472), .B(n_477), .Y(n_471) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_183), .B(n_341), .Y(n_417) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_184), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x6_ASAP7_75t_SL g241 ( .A(n_185), .B(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g266 ( .A(n_186), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_186), .B(n_301), .Y(n_319) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_186), .Y(n_457) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g274 ( .A(n_187), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_187), .B(n_230), .Y(n_299) );
INVx2_ASAP7_75t_L g327 ( .A(n_187), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_187), .B(n_194), .Y(n_368) );
BUFx3_ASAP7_75t_L g392 ( .A(n_187), .Y(n_392) );
OR2x2_ASAP7_75t_L g404 ( .A(n_187), .B(n_194), .Y(n_404) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_187), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_193), .A2(n_435), .B1(n_438), .B2(n_439), .Y(n_434) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_204), .Y(n_193) );
INVx1_ASAP7_75t_L g262 ( .A(n_194), .Y(n_262) );
OR2x2_ASAP7_75t_L g273 ( .A(n_194), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g280 ( .A(n_194), .Y(n_280) );
AND2x4_ASAP7_75t_SL g297 ( .A(n_194), .B(n_205), .Y(n_297) );
AND2x4_ASAP7_75t_L g302 ( .A(n_194), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g311 ( .A(n_194), .Y(n_311) );
OR2x2_ASAP7_75t_L g317 ( .A(n_194), .B(n_205), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_194), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_194), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_194), .B(n_299), .Y(n_433) );
OR2x2_ASAP7_75t_L g449 ( .A(n_194), .B(n_352), .Y(n_449) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_203), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_201), .Y(n_195) );
INVx2_ASAP7_75t_SL g284 ( .A(n_201), .Y(n_284) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_201), .A2(n_532), .B(n_536), .Y(n_531) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g225 ( .A(n_202), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_204), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_204), .B(n_266), .Y(n_382) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_229), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_205), .B(n_230), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_205), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_205), .B(n_274), .Y(n_278) );
INVx3_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
INVx1_ASAP7_75t_L g336 ( .A(n_205), .Y(n_336) );
AND2x2_ASAP7_75t_L g416 ( .A(n_205), .B(n_280), .Y(n_416) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_221), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B1(n_214), .B2(n_219), .Y(n_206) );
INVx1_ASAP7_75t_L g504 ( .A(n_209), .Y(n_504) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g545 ( .A(n_210), .Y(n_545) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
OR2x6_ASAP7_75t_L g475 ( .A(n_211), .B(n_218), .Y(n_475) );
INVxp33_ASAP7_75t_L g521 ( .A(n_211), .Y(n_521) );
INVx1_ASAP7_75t_L g546 ( .A(n_213), .Y(n_546) );
INVxp67_ASAP7_75t_L g502 ( .A(n_214), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx1_ASAP7_75t_L g522 ( .A(n_217), .Y(n_522) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_224), .A2(n_491), .B1(n_496), .B2(n_497), .Y(n_490) );
INVx3_ASAP7_75t_L g497 ( .A(n_224), .Y(n_497) );
INVx4_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_225), .A2(n_232), .B(n_238), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_225), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_228), .B(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_228), .A2(n_475), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_230), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_230), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g352 ( .A(n_230), .B(n_274), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_230), .B(n_303), .Y(n_369) );
INVx1_ASAP7_75t_L g375 ( .A(n_230), .Y(n_375) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_237), .Y(n_232) );
AOI222xp33_ASAP7_75t_SL g239 ( .A1(n_240), .A2(n_243), .B1(n_253), .B2(n_260), .C1(n_263), .C2(n_267), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_252), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_244), .B(n_313), .Y(n_364) );
AND2x4_ASAP7_75t_L g380 ( .A(n_244), .B(n_291), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g305 ( .A(n_256), .B(n_306), .Y(n_305) );
AOI222xp33_ASAP7_75t_L g270 ( .A1(n_257), .A2(n_271), .B1(n_276), .B2(n_281), .C1(n_289), .C2(n_831), .Y(n_270) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g409 ( .A(n_258), .B(n_313), .Y(n_409) );
OR2x2_ASAP7_75t_L g452 ( .A(n_258), .B(n_358), .Y(n_452) );
AND2x2_ASAP7_75t_L g281 ( .A(n_259), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_259), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_260), .A2(n_371), .B(n_376), .C(n_377), .Y(n_370) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g398 ( .A(n_262), .Y(n_398) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g328 ( .A(n_267), .Y(n_328) );
AND2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI31xp33_ASAP7_75t_L g363 ( .A1(n_271), .A2(n_289), .A3(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_272), .A2(n_322), .B(n_366), .C(n_367), .Y(n_365) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
OR2x2_ASAP7_75t_L g354 ( .A(n_273), .B(n_303), .Y(n_354) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
BUFx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
AND2x2_ASAP7_75t_L g331 ( .A(n_282), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_288), .Y(n_283) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_284), .A2(n_516), .B(n_524), .Y(n_515) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_284), .A2(n_516), .B(n_524), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_291), .B(n_348), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_304), .B(n_307), .C(n_329), .Y(n_292) );
INVxp33_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_295), .B(n_300), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g333 ( .A(n_297), .B(n_326), .Y(n_333) );
OR2x2_ASAP7_75t_L g309 ( .A(n_298), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g339 ( .A(n_298), .B(n_313), .Y(n_339) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g415 ( .A(n_299), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_302), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_302), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g450 ( .A(n_302), .B(n_326), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_302), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g393 ( .A(n_303), .B(n_375), .Y(n_393) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AOI322xp5_ASAP7_75t_L g447 ( .A1(n_306), .A2(n_326), .A3(n_380), .B1(n_405), .B2(n_448), .C1(n_450), .C2(n_451), .Y(n_447) );
AOI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_312), .B(n_314), .C(n_323), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_310), .B(n_338), .Y(n_360) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g325 ( .A(n_311), .B(n_326), .Y(n_325) );
NOR2x1p5_ASAP7_75t_L g391 ( .A(n_311), .B(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_311), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_312), .A2(n_330), .B(n_333), .C(n_334), .Y(n_329) );
AND2x4_ASAP7_75t_L g348 ( .A(n_313), .B(n_332), .Y(n_348) );
INVx2_ASAP7_75t_L g358 ( .A(n_313), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_313), .B(n_347), .Y(n_378) );
AND2x2_ASAP7_75t_L g420 ( .A(n_313), .B(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_313), .B(n_437), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_313), .B(n_341), .Y(n_459) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_320), .Y(n_314) );
AND2x2_ASAP7_75t_L g410 ( .A(n_316), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g338 ( .A(n_319), .Y(n_338) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_331), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B(n_339), .C(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_338), .Y(n_422) );
INVx3_ASAP7_75t_SL g437 ( .A(n_341), .Y(n_437) );
NAND5xp2_ASAP7_75t_L g343 ( .A(n_344), .B(n_363), .C(n_370), .D(n_383), .E(n_394), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B1(n_353), .B2(n_355), .C1(n_359), .C2(n_361), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_346), .A2(n_427), .B1(n_431), .B2(n_432), .Y(n_426) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g376 ( .A(n_347), .B(n_348), .Y(n_376) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_357), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_358), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_358), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g406 ( .A(n_358), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g436 ( .A(n_362), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_369), .Y(n_384) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_380), .A2(n_384), .B1(n_385), .B2(n_389), .Y(n_383) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g397 ( .A(n_382), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g402 ( .A(n_384), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_SL g430 ( .A(n_393), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_418), .C(n_441), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_417), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_408), .B2(n_410), .C(n_413), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g442 ( .A(n_404), .B(n_430), .Y(n_442) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
OAI321xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .A3(n_423), .B1(n_425), .B2(n_426), .C(n_434), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_432), .A2(n_454), .B1(n_458), .B2(n_459), .Y(n_453) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .B(n_447), .C(n_453), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_781), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_731), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_671), .B(n_730), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_463), .B(n_732), .C(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g822 ( .A(n_463), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_635), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_576), .C(n_605), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_565), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_486), .B1(n_525), .B2(n_537), .Y(n_466) );
NAND2x1_ASAP7_75t_L g767 ( .A(n_467), .B(n_566), .Y(n_767) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx2_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
INVx4_ASAP7_75t_L g581 ( .A(n_469), .Y(n_581) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_469), .Y(n_601) );
AND2x4_ASAP7_75t_L g612 ( .A(n_469), .B(n_580), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_469), .B(n_542), .Y(n_618) );
NOR2x1_ASAP7_75t_SL g691 ( .A(n_469), .B(n_553), .Y(n_691) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_L g492 ( .A(n_475), .Y(n_492) );
INVx2_ASAP7_75t_L g552 ( .A(n_475), .Y(n_552) );
INVx2_ASAP7_75t_L g584 ( .A(n_478), .Y(n_584) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_478), .Y(n_598) );
INVx1_ASAP7_75t_L g609 ( .A(n_478), .Y(n_609) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_478), .Y(n_621) );
AND2x2_ASAP7_75t_L g653 ( .A(n_478), .B(n_553), .Y(n_653) );
INVx1_ASAP7_75t_L g679 ( .A(n_478), .Y(n_679) );
AND2x2_ASAP7_75t_L g741 ( .A(n_478), .B(n_569), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_505), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g634 ( .A(n_488), .B(n_573), .Y(n_634) );
INVx2_ASAP7_75t_L g676 ( .A(n_488), .Y(n_676) );
AND2x2_ASAP7_75t_L g778 ( .A(n_488), .B(n_505), .Y(n_778) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_489), .B(n_528), .Y(n_572) );
INVx2_ASAP7_75t_L g593 ( .A(n_489), .Y(n_593) );
AND2x4_ASAP7_75t_L g615 ( .A(n_489), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g650 ( .A(n_489), .Y(n_650) );
AND2x2_ASAP7_75t_L g774 ( .A(n_489), .B(n_531), .Y(n_774) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_497), .A2(n_507), .B(n_513), .Y(n_506) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_497), .A2(n_507), .B(n_513), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g748 ( .A(n_505), .Y(n_748) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g623 ( .A(n_506), .B(n_593), .Y(n_623) );
AND2x2_ASAP7_75t_L g628 ( .A(n_506), .B(n_593), .Y(n_628) );
INVx2_ASAP7_75t_L g641 ( .A(n_506), .Y(n_641) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_506), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x4_ASAP7_75t_L g614 ( .A(n_514), .B(n_527), .Y(n_614) );
AND2x2_ASAP7_75t_L g629 ( .A(n_514), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g684 ( .A(n_514), .Y(n_684) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_515), .B(n_531), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_515), .B(n_528), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVxp33_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
INVx3_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_528), .Y(n_588) );
AND2x2_ASAP7_75t_L g702 ( .A(n_528), .B(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g645 ( .A(n_529), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_529), .B(n_684), .Y(n_725) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g592 ( .A(n_530), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g573 ( .A(n_531), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g616 ( .A(n_531), .Y(n_616) );
INVxp67_ASAP7_75t_L g630 ( .A(n_531), .Y(n_630) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_531), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_531), .Y(n_707) );
INVx1_ASAP7_75t_L g685 ( .A(n_537), .Y(n_685) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_538), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g727 ( .A(n_539), .B(n_568), .Y(n_727) );
OR2x2_ASAP7_75t_L g779 ( .A(n_540), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g678 ( .A(n_541), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g714 ( .A(n_541), .B(n_601), .Y(n_714) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_553), .Y(n_541) );
AND2x4_ASAP7_75t_L g568 ( .A(n_542), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g580 ( .A(n_542), .Y(n_580) );
INVx2_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_542), .Y(n_723) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .C(n_547), .Y(n_544) );
INVx3_ASAP7_75t_L g569 ( .A(n_553), .Y(n_569) );
INVx2_ASAP7_75t_L g663 ( .A(n_553), .Y(n_663) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B(n_564), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_567), .B(n_643), .Y(n_660) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_567), .B(n_581), .Y(n_752) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_568), .B(n_643), .Y(n_729) );
AND2x2_ASAP7_75t_L g596 ( .A(n_569), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g610 ( .A(n_569), .Y(n_610) );
AOI22xp5_ASAP7_75t_SL g658 ( .A1(n_570), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_658) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_571), .B(n_629), .Y(n_655) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g763 ( .A(n_572), .B(n_604), .Y(n_763) );
AND2x2_ASAP7_75t_L g586 ( .A(n_573), .B(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g622 ( .A(n_573), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g765 ( .A(n_573), .B(n_676), .Y(n_765) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g640 ( .A(n_575), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g666 ( .A(n_575), .Y(n_666) );
AND2x2_ASAP7_75t_L g701 ( .A(n_575), .B(n_593), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_585), .B1(n_589), .B2(n_594), .C(n_599), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g657 ( .A(n_579), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_579), .B(n_653), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_579), .B(n_741), .Y(n_740) );
AND2x4_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NOR2xp67_ASAP7_75t_SL g625 ( .A(n_581), .B(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
AND2x4_ASAP7_75t_SL g722 ( .A(n_581), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g769 ( .A(n_581), .B(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_584), .Y(n_780) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221x1_ASAP7_75t_L g733 ( .A1(n_586), .A2(n_734), .B1(n_736), .B2(n_737), .C(n_739), .Y(n_733) );
AND2x2_ASAP7_75t_L g659 ( .A(n_587), .B(n_615), .Y(n_659) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g602 ( .A(n_590), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_590), .B(n_592), .Y(n_776) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_596), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_596), .B(n_609), .Y(n_626) );
INVx2_ASAP7_75t_L g633 ( .A(n_596), .Y(n_633) );
INVx1_ASAP7_75t_L g695 ( .A(n_597), .Y(n_695) );
BUFx2_ASAP7_75t_L g715 ( .A(n_598), .Y(n_715) );
NAND2xp33_ASAP7_75t_SL g599 ( .A(n_600), .B(n_602), .Y(n_599) );
OR2x6_ASAP7_75t_L g632 ( .A(n_601), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g761 ( .A(n_601), .B(n_653), .Y(n_761) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_624), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_613), .B1(n_617), .B2(n_622), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_608), .B(n_612), .Y(n_670) );
AND2x4_ASAP7_75t_L g736 ( .A(n_608), .B(n_694), .Y(n_736) );
AND2x4_ASAP7_75t_SL g608 ( .A(n_609), .B(n_610), .Y(n_608) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_609), .Y(n_751) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_612), .B(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_612), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_612), .B(n_643), .Y(n_735) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g756 ( .A(n_614), .B(n_675), .Y(n_756) );
INVx3_ASAP7_75t_L g667 ( .A(n_615), .Y(n_667) );
AND2x2_ASAP7_75t_L g688 ( .A(n_615), .B(n_640), .Y(n_688) );
NAND2x1_ASAP7_75t_SL g759 ( .A(n_615), .B(n_666), .Y(n_759) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_631), .B2(n_634), .Y(n_624) );
BUFx2_ASAP7_75t_L g680 ( .A(n_626), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_627), .A2(n_718), .B1(n_727), .B2(n_728), .Y(n_726) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_628), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g648 ( .A(n_629), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_633), .B(n_713), .C(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g668 ( .A(n_634), .Y(n_668) );
AOI211x1_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_644), .B(n_646), .C(n_664), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_639), .B(n_727), .Y(n_746) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_640), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g718 ( .A(n_640), .B(n_676), .Y(n_718) );
AND2x2_ASAP7_75t_L g773 ( .A(n_640), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g696 ( .A(n_643), .Y(n_696) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g738 ( .A(n_645), .B(n_683), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_658), .Y(n_646) );
AOI22xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_651), .B1(n_654), .B2(n_656), .Y(n_647) );
BUFx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g711 ( .A(n_650), .B(n_706), .Y(n_711) );
INVx1_ASAP7_75t_SL g753 ( .A(n_650), .Y(n_753) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_653), .B(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g757 ( .A(n_662), .B(n_679), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_669), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_666), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g681 ( .A(n_667), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_671), .Y(n_824) );
NAND3x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_708), .C(n_716), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g782 ( .A(n_672), .B(n_708), .C(n_716), .D(n_783), .Y(n_782) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_686), .Y(n_672) );
OAI222xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B1(n_680), .B2(n_681), .C1(n_683), .C2(n_685), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g760 ( .A1(n_678), .A2(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_679), .B(n_694), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_682), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_697), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_690), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_694), .B(n_696), .Y(n_699) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_704), .B2(n_705), .Y(n_697) );
AND2x4_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g705 ( .A(n_701), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_709), .B(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g742 ( .A(n_711), .Y(n_742) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_726), .Y(n_716) );
AOI22xp5_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp33_ASAP7_75t_L g731 ( .A(n_730), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g823 ( .A(n_732), .Y(n_823) );
NAND3x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_744), .C(n_764), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_736), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g770 ( .A(n_741), .Y(n_770) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_745), .B(n_754), .Y(n_744) );
AOI21xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_747), .B(n_753), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_760), .Y(n_754) );
INVx2_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_759), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_768), .B2(n_771), .C(n_775), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g825 ( .A(n_787), .B(n_826), .C(n_827), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_793), .Y(n_787) );
INVxp33_ASAP7_75t_L g800 ( .A(n_788), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_793), .Y(n_799) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR2x1_ASAP7_75t_R g802 ( .A(n_796), .B(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_799), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_803), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_811), .B(n_825), .Y(n_804) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
BUFx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_813), .A2(n_814), .B1(n_820), .B2(n_821), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_818), .B2(n_819), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AND3x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .C(n_824), .Y(n_821) );
endmodule