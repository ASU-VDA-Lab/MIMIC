module fake_jpeg_9443_n_311 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_20),
.B(n_18),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_59),
.B1(n_27),
.B2(n_34),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_23),
.B1(n_26),
.B2(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_44),
.B1(n_40),
.B2(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_17),
.B1(n_34),
.B2(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_28),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_76),
.B1(n_81),
.B2(n_38),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_84),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_75),
.B1(n_85),
.B2(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_44),
.B1(n_36),
.B2(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_44),
.B1(n_41),
.B2(n_37),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_36),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_90),
.B(n_1),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_44),
.B1(n_41),
.B2(n_36),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_43),
.B(n_32),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_43),
.B(n_38),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_17),
.B1(n_18),
.B2(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_89),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_35),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_43),
.C(n_38),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_12),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_12),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_33),
.B(n_22),
.C(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_125),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_112),
.B(n_121),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_43),
.B1(n_30),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_124),
.B1(n_68),
.B2(n_72),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_127),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_32),
.B(n_33),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_10),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_73),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_1),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_122),
.B(n_119),
.Y(n_147)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_143),
.B1(n_157),
.B2(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_74),
.B1(n_78),
.B2(n_71),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_117),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_157),
.C(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_150),
.B(n_98),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_104),
.B(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_104),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_103),
.B1(n_68),
.B2(n_100),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_67),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_67),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_96),
.B1(n_90),
.B2(n_95),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_173),
.B(n_184),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_168),
.C(n_171),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_105),
.B1(n_123),
.B2(n_112),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_193),
.B1(n_97),
.B2(n_162),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_142),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_183),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_110),
.B(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_123),
.B1(n_112),
.B2(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_189),
.B1(n_150),
.B2(n_146),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_73),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_125),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_75),
.B(n_91),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_149),
.B(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_148),
.B1(n_159),
.B2(n_140),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_94),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_92),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_152),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_133),
.A2(n_135),
.B1(n_151),
.B2(n_141),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_184),
.B1(n_173),
.B2(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_192),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_129),
.B1(n_181),
.B2(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_213),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_169),
.C(n_166),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_215),
.B1(n_217),
.B2(n_182),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_214),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_165),
.A2(n_80),
.B(n_79),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_80),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_93),
.B1(n_70),
.B2(n_129),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_113),
.B(n_32),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_129),
.B1(n_120),
.B2(n_99),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_166),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_239),
.C(n_204),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_172),
.B1(n_175),
.B2(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_167),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_241),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_200),
.B1(n_216),
.B2(n_189),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_242),
.B(n_198),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_171),
.B1(n_194),
.B2(n_168),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_195),
.A2(n_183),
.B1(n_190),
.B2(n_118),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_208),
.B1(n_218),
.B2(n_217),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_106),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_201),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_118),
.C(n_83),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_88),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_255),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_254),
.C(n_257),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_248),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_201),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_204),
.B(n_213),
.C(n_214),
.D(n_195),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_205),
.C(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_221),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_224),
.B1(n_234),
.B2(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_266),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_229),
.B1(n_237),
.B2(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_214),
.B1(n_235),
.B2(n_226),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_270),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_255),
.B1(n_257),
.B2(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_273),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_251),
.B(n_250),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_283),
.B(n_9),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_233),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_284),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_231),
.B(n_269),
.Y(n_283)
);

NAND4xp25_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_219),
.C(n_220),
.D(n_199),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_254),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_263),
.C(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_270),
.C(n_245),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_294),
.C(n_11),
.Y(n_302)
);

AOI31xp33_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_261),
.A3(n_266),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_242),
.C(n_220),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_10),
.B(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_301),
.A3(n_11),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_5),
.B1(n_8),
.B2(n_13),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_22),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_281),
.B1(n_277),
.B2(n_6),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_13),
.C(n_15),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_304),
.A3(n_305),
.B1(n_306),
.B2(n_16),
.C1(n_4),
.C2(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_299),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_308),
.B(n_296),
.C(n_16),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_16),
.Y(n_311)
);


endmodule