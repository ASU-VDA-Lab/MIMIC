module fake_jpeg_23723_n_244 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_58),
.B1(n_24),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_14),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_20),
.B1(n_32),
.B2(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_51),
.B1(n_55),
.B2(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_29),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_13),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_57),
.B1(n_45),
.B2(n_41),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_75),
.B1(n_59),
.B2(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_14),
.B1(n_26),
.B2(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_98),
.B(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_71),
.B1(n_65),
.B2(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_77),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_90),
.B1(n_98),
.B2(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_94),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_45),
.A3(n_35),
.B1(n_38),
.B2(n_47),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_40),
.A3(n_16),
.B1(n_43),
.B2(n_50),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_51),
.B1(n_42),
.B2(n_21),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_62),
.B1(n_28),
.B2(n_27),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_39),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_14),
.B1(n_28),
.B2(n_27),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_74),
.B1(n_73),
.B2(n_71),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_34),
.CI(n_31),
.CON(n_96),
.SN(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_23),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_99),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_108),
.B1(n_116),
.B2(n_119),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_1),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_111),
.B(n_115),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_23),
.B(n_31),
.C(n_34),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_65),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_84),
.B1(n_99),
.B2(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_81),
.B1(n_90),
.B2(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_31),
.B1(n_40),
.B2(n_34),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_121),
.Y(n_157)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_18),
.B(n_23),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_127),
.B(n_139),
.Y(n_147)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_R g127 ( 
.A(n_115),
.B(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_140),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_21),
.B(n_23),
.Y(n_161)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_23),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_101),
.B1(n_91),
.B2(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_152),
.B1(n_158),
.B2(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_117),
.C(n_103),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_162),
.C(n_123),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_105),
.B1(n_118),
.B2(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_120),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_129),
.B(n_122),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_18),
.B1(n_16),
.B2(n_21),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_60),
.B(n_93),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_155),
.B(n_131),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_21),
.B1(n_23),
.B2(n_16),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_50),
.B1(n_43),
.B2(n_93),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_50),
.B1(n_43),
.B2(n_93),
.Y(n_159)
);

XNOR2x2_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_139),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_23),
.C(n_2),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_123),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_171),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_157),
.B1(n_8),
.B2(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_174),
.C(n_180),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_156),
.B1(n_151),
.B2(n_143),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_135),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_132),
.B(n_135),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_173),
.B(n_154),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_128),
.B(n_125),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_129),
.C(n_133),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_124),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_7),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_7),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_1),
.C(n_3),
.Y(n_180)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_155),
.A3(n_148),
.B1(n_145),
.B2(n_154),
.C1(n_153),
.C2(n_143),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_184),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_151),
.B1(n_148),
.B2(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_190),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_159),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_168),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_176),
.C(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_208),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_166),
.B(n_178),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_205),
.A2(n_181),
.B(n_179),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_175),
.C(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_216),
.B(n_217),
.C(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_12),
.C(n_6),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_193),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_215),
.B1(n_218),
.B2(n_9),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_205),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_6),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_200),
.B(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_227),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_206),
.C(n_204),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_225),
.B(n_217),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_9),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_10),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_231),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_209),
.Y(n_231)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_226),
.B(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_5),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_12),
.B1(n_5),
.B2(n_10),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_5),
.B(n_11),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_223),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.C(n_230),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_236),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_240),
.B(n_1),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_4),
.Y(n_244)
);


endmodule