module fake_jpeg_19201_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_82),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_64),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_59),
.B(n_62),
.C(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_60),
.B1(n_73),
.B2(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_55),
.B1(n_64),
.B2(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_73),
.B1(n_68),
.B2(n_74),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_69),
.B1(n_64),
.B2(n_55),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_107),
.B1(n_90),
.B2(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_103),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_71),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_57),
.A3(n_66),
.B1(n_65),
.B2(n_3),
.Y(n_121)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_57),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_52),
.B1(n_53),
.B2(n_72),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_50),
.B1(n_75),
.B2(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_114),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_58),
.C(n_63),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_90),
.B(n_76),
.C(n_54),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_111),
.B(n_110),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_14),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_16),
.A3(n_47),
.B1(n_45),
.B2(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_17),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_96),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_136),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_109),
.C(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_143),
.C(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_134),
.B1(n_4),
.B2(n_5),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_13),
.C(n_33),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_48),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_131),
.B1(n_125),
.B2(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_144),
.B1(n_145),
.B2(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_150),
.C(n_152),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_151),
.B1(n_147),
.B2(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_29),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_27),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_141),
.B(n_26),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_24),
.C(n_18),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_3),
.B(n_4),
.C(n_6),
.D(n_8),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_9),
.B(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_9),
.Y(n_163)
);


endmodule