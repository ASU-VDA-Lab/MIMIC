module fake_netlist_5_2351_n_1994 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1994);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1994;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_44),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_15),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_79),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_107),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_39),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_19),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_94),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_71),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_67),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_65),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_30),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_125),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_178),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_65),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_95),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_143),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_26),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_180),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_38),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_171),
.Y(n_256)
);

BUFx8_ASAP7_75t_SL g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_25),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_62),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_86),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_105),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_80),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_32),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_159),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_147),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_44),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_0),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_87),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_56),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_185),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_191),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_43),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_121),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_113),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_0),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_112),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_99),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_177),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_78),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_173),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_38),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_83),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_104),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_97),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_118),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_96),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_11),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_114),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_151),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_186),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_42),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_35),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_45),
.Y(n_312)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_163),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_63),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_103),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_14),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_14),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_72),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_47),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_134),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_199),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_156),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_111),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_135),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_47),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_162),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_70),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_92),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_33),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_193),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_49),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_12),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_74),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_164),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_144),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_57),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_21),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_133),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_12),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_51),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_183),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_48),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_41),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_174),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_60),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_13),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_7),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_18),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_36),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_52),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_37),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_84),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_194),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_139),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_35),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_197),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_68),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_19),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_149),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_120),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_158),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_117),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_106),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_188),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_11),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_7),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_49),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_37),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_175),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_66),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_8),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_81),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_140),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_45),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_85),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_145),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_4),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_59),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_165),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_91),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_122),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_154),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_33),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_57),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_1),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_179),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_93),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_28),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_137),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_8),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_182),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_27),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_176),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_397),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_228),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_255),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_255),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_216),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_216),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_230),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_255),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_255),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_313),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_204),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_215),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_246),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_204),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_294),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_211),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_315),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_211),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_287),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_203),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_203),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_253),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_217),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_315),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_380),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_221),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_328),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_221),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_287),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_239),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_233),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_232),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_232),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_251),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_251),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_259),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_259),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_282),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_282),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_206),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_212),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_231),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_235),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_233),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_336),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_280),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_260),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_205),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_336),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_243),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_248),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_254),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_287),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_261),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_280),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_263),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_313),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_202),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_239),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_209),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_220),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_202),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_392),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_368),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_316),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_274),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_274),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_348),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_267),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_268),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_271),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_322),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_324),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_272),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_339),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_222),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_368),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_223),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_347),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_352),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_375),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_310),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_310),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_236),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_278),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_236),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_241),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_310),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_225),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_226),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_279),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_285),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_503),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_438),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

CKINVDCx11_ASAP7_75t_R g516 ( 
.A(n_414),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_416),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_500),
.A2(n_332),
.B(n_279),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_424),
.B(n_332),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_432),
.B(n_244),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_416),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_436),
.B(n_241),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_404),
.B(n_250),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_474),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_413),
.A2(n_265),
.B(n_262),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_474),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_442),
.B(n_348),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_417),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_413),
.A2(n_283),
.B(n_266),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_469),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_418),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_447),
.B(n_348),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_469),
.B(n_202),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_419),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_420),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_408),
.B(n_314),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_406),
.B(n_286),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_409),
.B(n_443),
.C(n_441),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_422),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_417),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_423),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_500),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_457),
.B(n_218),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_433),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_502),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_507),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_459),
.B(n_202),
.Y(n_566)
);

CKINVDCx11_ASAP7_75t_R g567 ( 
.A(n_425),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_486),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_421),
.B(n_213),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_430),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_430),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_444),
.B(n_237),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_435),
.Y(n_574)
);

BUFx8_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_407),
.B(n_290),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_445),
.B(n_306),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_427),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_218),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_489),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_448),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_433),
.B(n_224),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_429),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_489),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_429),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_439),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_472),
.A2(n_295),
.B(n_292),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_473),
.B(n_297),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_454),
.B(n_224),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_490),
.B(n_308),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_439),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_591),
.A2(n_329),
.B(n_309),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_550),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_592),
.A2(n_492),
.B1(n_506),
.B2(n_505),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_566),
.Y(n_599)
);

INVx8_ASAP7_75t_L g600 ( 
.A(n_586),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_517),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

NAND3xp33_ASAP7_75t_L g604 ( 
.A(n_523),
.B(n_528),
.C(n_592),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_566),
.B(n_570),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_545),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_434),
.C(n_410),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_224),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_561),
.B(n_428),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_561),
.B(n_431),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_566),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_524),
.A2(n_401),
.B1(n_482),
.B2(n_456),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_591),
.A2(n_341),
.B(n_337),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_537),
.A2(n_401),
.B1(n_482),
.B2(n_456),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_580),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_562),
.B(n_475),
.Y(n_621)
);

OAI21xp33_ASAP7_75t_SL g622 ( 
.A1(n_548),
.A2(n_494),
.B(n_493),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_580),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_516),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_580),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_580),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_594),
.B(n_483),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_562),
.B(n_483),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_510),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_519),
.B(n_402),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_548),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_575),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_514),
.B(n_496),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_594),
.B(n_485),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_510),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_567),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_532),
.B(n_471),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_532),
.B(n_471),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_587),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_585),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_513),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_577),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_478),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_517),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_594),
.B(n_224),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_537),
.B(n_440),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_514),
.B(n_485),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_547),
.B(n_488),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_547),
.B(n_488),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_594),
.B(n_498),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_548),
.A2(n_450),
.B1(n_451),
.B2(n_449),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_532),
.B(n_460),
.C(n_452),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_582),
.B(n_498),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_555),
.B(n_466),
.C(n_464),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_582),
.B(n_501),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_585),
.B(n_351),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_554),
.B(n_478),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_513),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_575),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_573),
.A2(n_242),
.B1(n_258),
.B2(n_207),
.Y(n_668)
);

AOI21x1_ASAP7_75t_L g669 ( 
.A1(n_522),
.A2(n_371),
.B(n_363),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_573),
.B(n_501),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_517),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_520),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_590),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_590),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_590),
.Y(n_678)
);

AO21x1_ASAP7_75t_L g679 ( 
.A1(n_554),
.A2(n_394),
.B(n_389),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_556),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_520),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_554),
.A2(n_576),
.B1(n_552),
.B2(n_578),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_526),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_538),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_518),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_526),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_518),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_590),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_574),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_535),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_578),
.B(n_508),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_590),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_527),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_518),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_527),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_518),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_554),
.B(n_479),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_557),
.B(n_508),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_575),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_586),
.B(n_454),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_575),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_533),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_533),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_522),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_539),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_595),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_586),
.B(n_458),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_595),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_539),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_552),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_540),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_571),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_595),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_586),
.B(n_227),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_595),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_576),
.B(n_463),
.C(n_461),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_540),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_542),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_542),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_595),
.Y(n_723)
);

INVx4_ASAP7_75t_SL g724 ( 
.A(n_586),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_531),
.B(n_458),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_576),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_551),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_518),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_518),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_R g731 ( 
.A(n_512),
.B(n_522),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_546),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_551),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_586),
.B(n_481),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_586),
.B(n_227),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_586),
.B(n_481),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_530),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_546),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_555),
.B(n_396),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_558),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_558),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_551),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_559),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_641),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_661),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_712),
.B(n_426),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_690),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_641),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_649),
.B(n_499),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_605),
.B(n_531),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_643),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_653),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_599),
.A2(n_593),
.B1(n_453),
.B2(n_455),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_606),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_229),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_599),
.B(n_563),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_606),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_632),
.A2(n_522),
.B1(n_541),
.B2(n_535),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_611),
.B(n_307),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_671),
.B(n_317),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_615),
.B(n_563),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_712),
.B(n_219),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_632),
.B(n_227),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_R g766 ( 
.A(n_631),
.B(n_437),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_653),
.B(n_504),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_632),
.B(n_227),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_680),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_SL g770 ( 
.A(n_615),
.B(n_207),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_628),
.B(n_219),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_604),
.B(n_563),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_706),
.B(n_298),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_706),
.A2(n_530),
.B(n_515),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_563),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_622),
.A2(n_541),
.B1(n_258),
.B2(n_281),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_607),
.A2(n_398),
.B1(n_494),
.B2(n_493),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_663),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_650),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_658),
.B(n_564),
.Y(n_780)
);

NAND2x1_ASAP7_75t_L g781 ( 
.A(n_673),
.B(n_511),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_733),
.B(n_564),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_740),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_682),
.B(n_613),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_613),
.B(n_564),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_625),
.B(n_564),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_706),
.B(n_298),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_665),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_622),
.A2(n_242),
.B1(n_372),
.B2(n_349),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_644),
.B(n_568),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_379),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_629),
.B(n_379),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_621),
.B(n_382),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_690),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_625),
.B(n_593),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_731),
.A2(n_593),
.B1(n_476),
.B2(n_491),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_630),
.B(n_593),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_691),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_665),
.Y(n_799)
);

INVx8_ASAP7_75t_L g800 ( 
.A(n_664),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_638),
.B(n_593),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_607),
.B(n_382),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_655),
.A2(n_593),
.B1(n_302),
.B2(n_303),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_664),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_638),
.B(n_593),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_690),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_648),
.B(n_583),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_648),
.B(n_583),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_597),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_603),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_714),
.B(n_569),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_666),
.B(n_583),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_659),
.B(n_298),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_666),
.B(n_583),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_674),
.B(n_559),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_714),
.B(n_636),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_598),
.B(n_383),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_644),
.B(n_647),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_674),
.B(n_559),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_689),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_647),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_656),
.A2(n_330),
.B1(n_264),
.B2(n_270),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_619),
.B(n_383),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_697),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_681),
.B(n_559),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_636),
.B(n_569),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_681),
.A2(n_588),
.B(n_584),
.C(n_581),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_683),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_633),
.B(n_477),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_683),
.B(n_559),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_686),
.B(n_559),
.Y(n_831)
);

AO221x1_ASAP7_75t_L g832 ( 
.A1(n_616),
.A2(n_298),
.B1(n_369),
.B2(n_319),
.C(n_301),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_647),
.B(n_301),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_686),
.B(n_544),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_725),
.B(n_387),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_693),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_693),
.B(n_387),
.Y(n_837)
);

O2A1O1Ixp5_ASAP7_75t_L g838 ( 
.A1(n_669),
.A2(n_515),
.B(n_534),
.C(n_536),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_695),
.B(n_544),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_679),
.A2(n_372),
.B1(n_281),
.B2(n_300),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_660),
.B(n_719),
.C(n_662),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_727),
.B(n_301),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_695),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_702),
.A2(n_588),
.B(n_584),
.C(n_581),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_702),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_679),
.A2(n_300),
.B1(n_349),
.B2(n_579),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_727),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_636),
.B(n_579),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_705),
.B(n_388),
.Y(n_849)
);

BUFx5_ASAP7_75t_L g850 ( 
.A(n_608),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_664),
.A2(n_289),
.B1(n_208),
.B2(n_210),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_707),
.B(n_544),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_707),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_636),
.B(n_388),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_711),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_728),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_664),
.A2(n_291),
.B1(n_214),
.B2(n_234),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_684),
.B(n_393),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_728),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_SL g860 ( 
.A(n_633),
.B(n_257),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_734),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_711),
.B(n_553),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_684),
.B(n_393),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_734),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_713),
.B(n_293),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_713),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_660),
.B(n_560),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_720),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_720),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_667),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_684),
.B(n_238),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_721),
.B(n_553),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_721),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_722),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_743),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_684),
.B(n_717),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_717),
.B(n_240),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_743),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_732),
.B(n_739),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_609),
.B(n_301),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_739),
.B(n_553),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_596),
.A2(n_313),
.B1(n_386),
.B2(n_369),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_609),
.B(n_319),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_612),
.B(n_319),
.Y(n_884)
);

AO22x2_ASAP7_75t_L g885 ( 
.A1(n_668),
.A2(n_495),
.B1(n_497),
.B2(n_565),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_741),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_741),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_742),
.B(n_553),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_742),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_608),
.B(n_553),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_608),
.B(n_553),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_698),
.B(n_296),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_612),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_620),
.B(n_319),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_596),
.A2(n_386),
.B1(n_313),
.B2(n_369),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_596),
.A2(n_617),
.B1(n_652),
.B2(n_608),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_756),
.B(n_717),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

BUFx12f_ASAP7_75t_L g899 ( 
.A(n_870),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_886),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_811),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_887),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_821),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_746),
.B(n_667),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_889),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_847),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_756),
.B(n_608),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_778),
.B(n_699),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_828),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_836),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_747),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_820),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_826),
.B(n_699),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_760),
.B(n_668),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_753),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_879),
.B(n_652),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_821),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_821),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_843),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_879),
.B(n_652),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_845),
.Y(n_922)
);

NOR2x2_ASAP7_75t_L g923 ( 
.A(n_829),
.B(n_740),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_864),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_761),
.B(n_652),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_748),
.B(n_724),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_853),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_855),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_866),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_654),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_798),
.B(n_635),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_767),
.B(n_701),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_848),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_748),
.B(n_794),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_868),
.B(n_869),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_873),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_796),
.B(n_689),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_802),
.A2(n_700),
.B(n_735),
.C(n_709),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_874),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_809),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_745),
.B(n_740),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_783),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_766),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_748),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_821),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_766),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_856),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_790),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_780),
.B(n_652),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_751),
.B(n_740),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_790),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_859),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_771),
.B(n_673),
.Y(n_954)
);

BUFx12f_ASAP7_75t_SL g955 ( 
.A(n_829),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_771),
.B(n_791),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_816),
.B(n_624),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_783),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_751),
.B(n_737),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_791),
.B(n_724),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_861),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_749),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_875),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_748),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_892),
.B(n_724),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_896),
.A2(n_744),
.B(n_646),
.C(n_645),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_770),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_752),
.B(n_673),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_SL g969 ( 
.A(n_823),
.B(n_395),
.C(n_392),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_892),
.B(n_724),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_878),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_754),
.B(n_726),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_755),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_758),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_870),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_762),
.B(n_673),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_802),
.B(n_600),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_773),
.A2(n_669),
.B(n_623),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_794),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_750),
.B(n_600),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_794),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_794),
.B(n_620),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_773),
.A2(n_600),
.B(n_617),
.Y(n_983)
);

NOR2x2_ASAP7_75t_L g984 ( 
.A(n_829),
.B(n_624),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_806),
.B(n_850),
.Y(n_985)
);

OAI22xp33_ASAP7_75t_L g986 ( 
.A1(n_784),
.A2(n_395),
.B1(n_399),
.B2(n_362),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_787),
.A2(n_626),
.B(n_623),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_779),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_885),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_806),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_788),
.B(n_639),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_764),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_799),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_806),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_787),
.A2(n_600),
.B(n_626),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_806),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_824),
.B(n_257),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_817),
.B(n_639),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_789),
.B(n_365),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_772),
.B(n_627),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_782),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_800),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_837),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_835),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_800),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_841),
.B(n_495),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_793),
.B(n_304),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_837),
.B(n_651),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_800),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_775),
.A2(n_763),
.B(n_757),
.Y(n_1010)
);

CKINVDCx6p67_ASAP7_75t_R g1011 ( 
.A(n_876),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_867),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_849),
.B(n_651),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_765),
.A2(n_768),
.B(n_896),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_849),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_850),
.B(n_627),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_865),
.B(n_672),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_776),
.A2(n_313),
.B1(n_386),
.B2(n_369),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_SL g1019 ( 
.A(n_835),
.B(n_399),
.C(n_312),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_841),
.B(n_497),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_850),
.B(n_640),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_804),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_885),
.Y(n_1023)
);

BUFx5_ASAP7_75t_L g1024 ( 
.A(n_850),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_865),
.B(n_672),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_818),
.A2(n_646),
.B1(n_640),
.B2(n_657),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_789),
.B(n_792),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_871),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_818),
.A2(n_692),
.B1(n_645),
.B2(n_657),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_804),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_877),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_885),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_776),
.B(n_672),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_777),
.B(n_685),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_854),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_882),
.A2(n_313),
.B1(n_386),
.B2(n_400),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_777),
.B(n_685),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_858),
.B(n_305),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_765),
.A2(n_642),
.B1(n_670),
.B2(n_676),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_785),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_768),
.A2(n_642),
.B1(n_670),
.B2(n_676),
.Y(n_1042)
);

AND2x6_ASAP7_75t_L g1043 ( 
.A(n_795),
.B(n_677),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_863),
.B(n_840),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_759),
.A2(n_600),
.B(n_678),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_777),
.B(n_685),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_804),
.A2(n_710),
.B1(n_678),
.B2(n_692),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_786),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_774),
.A2(n_703),
.B(n_688),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_807),
.B(n_687),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_808),
.B(n_687),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_812),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_814),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_827),
.B(n_687),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_810),
.B(n_844),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_851),
.A2(n_703),
.B1(n_688),
.B2(n_704),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_822),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_838),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_815),
.B(n_694),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_857),
.B(n_704),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_834),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_840),
.B(n_318),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_852),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_781),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_862),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_819),
.B(n_694),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_872),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_881),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_860),
.B(n_320),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_850),
.B(n_708),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1018),
.A2(n_846),
.B1(n_882),
.B2(n_895),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_897),
.B(n_846),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_912),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_956),
.A2(n_833),
.B(n_813),
.C(n_830),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_973),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_909),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1003),
.B(n_825),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_910),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_914),
.A2(n_842),
.B(n_894),
.C(n_880),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_924),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1049),
.A2(n_759),
.B(n_888),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1002),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_SL g1084 ( 
.A(n_955),
.B(n_365),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1018),
.A2(n_797),
.B1(n_801),
.B2(n_805),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_977),
.A2(n_618),
.B(n_601),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1045),
.A2(n_618),
.B(n_601),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1003),
.B(n_1015),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_831),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1015),
.B(n_832),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_951),
.B(n_708),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_943),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_991),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_943),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1037),
.A2(n_803),
.B1(n_891),
.B2(n_890),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1045),
.A2(n_618),
.B(n_601),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_934),
.B(n_850),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_931),
.B(n_323),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_983),
.A2(n_634),
.B(n_618),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_991),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1031),
.B(n_710),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1053),
.B(n_715),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1037),
.A2(n_331),
.B1(n_335),
.B2(n_338),
.Y(n_1103)
);

BUFx4f_ASAP7_75t_L g1104 ( 
.A(n_899),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1044),
.A2(n_951),
.B1(n_1057),
.B2(n_938),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_983),
.A2(n_634),
.B(n_602),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_L g1107 ( 
.A(n_944),
.B(n_947),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_920),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1053),
.B(n_715),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_959),
.A2(n_884),
.B(n_883),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1006),
.B(n_718),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1010),
.A2(n_634),
.B(n_602),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1031),
.B(n_718),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1010),
.A2(n_884),
.B(n_883),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1041),
.B(n_723),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1014),
.A2(n_377),
.B1(n_343),
.B2(n_344),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_915),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1063),
.A2(n_894),
.B(n_716),
.C(n_736),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1027),
.A2(n_386),
.B1(n_400),
.B2(n_723),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_941),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_975),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_974),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_911),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1004),
.B(n_245),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_995),
.A2(n_634),
.B(n_602),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1007),
.A2(n_738),
.B(n_730),
.C(n_729),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_922),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_L g1129 ( 
.A1(n_960),
.A2(n_738),
.B(n_730),
.C(n_729),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_1007),
.A2(n_738),
.B(n_730),
.C(n_729),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_901),
.B(n_381),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1048),
.B(n_696),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1052),
.B(n_696),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_928),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1033),
.A2(n_373),
.B1(n_353),
.B2(n_354),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_932),
.B(n_247),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1063),
.B(n_350),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_954),
.A2(n_525),
.B(n_521),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_926),
.A2(n_696),
.B(n_589),
.C(n_479),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_957),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_933),
.B(n_355),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_SL g1143 ( 
.A(n_1029),
.B(n_378),
.C(n_356),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_942),
.B(n_480),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_948),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_989),
.A2(n_357),
.B1(n_358),
.B2(n_374),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_936),
.A2(n_930),
.B(n_929),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_979),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_937),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_945),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_953),
.Y(n_1151)
);

NAND2x1_ASAP7_75t_L g1152 ( 
.A(n_945),
.B(n_602),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_933),
.B(n_967),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1062),
.B(n_602),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_942),
.B(n_249),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_999),
.A2(n_480),
.B(n_484),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_992),
.A2(n_360),
.B1(n_256),
.B2(n_269),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_940),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_1039),
.B(n_364),
.C(n_273),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1069),
.B(n_675),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_1039),
.A2(n_589),
.B(n_515),
.C(n_511),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1036),
.B(n_252),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1032),
.A2(n_381),
.B1(n_277),
.B2(n_284),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_995),
.A2(n_675),
.B(n_614),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_907),
.A2(n_525),
.B(n_536),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_939),
.A2(n_511),
.B(n_521),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_945),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1006),
.B(n_275),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_981),
.A2(n_675),
.B(n_614),
.Y(n_1169)
);

BUFx8_ASAP7_75t_L g1170 ( 
.A(n_1023),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_961),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1020),
.B(n_997),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1011),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_963),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1002),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_972),
.A2(n_366),
.B(n_299),
.C(n_321),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_981),
.B(n_288),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1020),
.B(n_325),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_958),
.B(n_326),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1061),
.B(n_327),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_962),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1012),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1017),
.A2(n_525),
.B(n_543),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_913),
.B(n_333),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_994),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_994),
.A2(n_614),
.B(n_530),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1019),
.B(n_370),
.C(n_340),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_998),
.A2(n_376),
.B(n_342),
.C(n_345),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_964),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_984),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_987),
.A2(n_543),
.B(n_534),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_988),
.B(n_334),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_993),
.B(n_359),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1005),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_400),
.B1(n_361),
.B2(n_367),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_949),
.B(n_381),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_L g1198 ( 
.A(n_1070),
.B(n_521),
.C(n_534),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_R g1199 ( 
.A(n_1005),
.B(n_73),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_978),
.A2(n_543),
.B(n_614),
.Y(n_1200)
);

BUFx8_ASAP7_75t_L g1201 ( 
.A(n_1005),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1064),
.B(n_386),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_916),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1066),
.B(n_530),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_964),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_904),
.B(n_2),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_985),
.A2(n_530),
.B(n_198),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1068),
.B(n_4),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1025),
.B(n_900),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_952),
.B(n_195),
.Y(n_1210)
);

INVxp67_ASAP7_75t_SL g1211 ( 
.A(n_964),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_908),
.B(n_9),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_1009),
.B(n_9),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1165),
.A2(n_1046),
.A3(n_1035),
.B(n_1038),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1081),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1126),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1137),
.A2(n_1019),
.B(n_969),
.C(n_1060),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1166),
.A2(n_1013),
.B(n_1008),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1144),
.B(n_1141),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1121),
.Y(n_1220)
);

AO21x1_ASAP7_75t_L g1221 ( 
.A1(n_1072),
.A2(n_970),
.B(n_965),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1098),
.B(n_986),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1148),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1072),
.A2(n_921),
.A3(n_1058),
.B(n_950),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1166),
.A2(n_1054),
.B(n_1055),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1073),
.B(n_902),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1105),
.A2(n_1022),
.B1(n_1009),
.B2(n_1047),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1112),
.A2(n_1125),
.B(n_1096),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1197),
.B(n_905),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_982),
.B(n_1067),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1127),
.A2(n_1051),
.A3(n_1050),
.B(n_1059),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1191),
.A2(n_982),
.B(n_1042),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1106),
.A2(n_1099),
.B(n_1086),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1088),
.B(n_971),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1209),
.A2(n_980),
.B(n_966),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1200),
.A2(n_1040),
.B(n_935),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1209),
.A2(n_935),
.B(n_985),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_996),
.B(n_964),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1164),
.A2(n_1030),
.B(n_1026),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1172),
.B(n_1140),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_SL g1241 ( 
.A1(n_1091),
.A2(n_1207),
.B(n_1089),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1114),
.A2(n_996),
.B(n_1024),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1153),
.B(n_1009),
.Y(n_1243)
);

AND2x6_ASAP7_75t_L g1244 ( 
.A(n_1083),
.B(n_1009),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1083),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1091),
.A2(n_1195),
.A3(n_1085),
.B(n_1095),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1195),
.A2(n_976),
.A3(n_968),
.B(n_898),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1142),
.A2(n_1147),
.B(n_1212),
.C(n_1206),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1148),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1093),
.B(n_1022),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1078),
.B(n_903),
.Y(n_1251)
);

AO22x1_ASAP7_75t_L g1252 ( 
.A1(n_1173),
.A2(n_1022),
.B1(n_1000),
.B2(n_917),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1074),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1077),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1100),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1183),
.A2(n_1071),
.B(n_1016),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1130),
.A2(n_1056),
.B(n_1016),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1144),
.B(n_906),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1116),
.B(n_919),
.C(n_925),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1131),
.B(n_1022),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1089),
.B(n_903),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1079),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1138),
.A2(n_1071),
.B(n_1021),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1120),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1104),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1108),
.B(n_917),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1185),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1201),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1128),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1161),
.A2(n_927),
.B(n_1000),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_SL g1271 ( 
.A1(n_1208),
.A2(n_946),
.B(n_1000),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1134),
.B(n_918),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1149),
.B(n_990),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1090),
.A2(n_946),
.B(n_1000),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1082),
.A2(n_1024),
.B(n_1065),
.Y(n_1275)
);

BUFx4f_ASAP7_75t_L g1276 ( 
.A(n_1175),
.Y(n_1276)
);

NOR2x1_ASAP7_75t_R g1277 ( 
.A(n_1190),
.B(n_923),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1201),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1075),
.A2(n_1000),
.B(n_1043),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1210),
.A2(n_1028),
.B(n_1065),
.C(n_1043),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1080),
.A2(n_1118),
.B(n_1159),
.C(n_1184),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1158),
.B(n_1028),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1168),
.A2(n_1043),
.B(n_1024),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1117),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1182),
.A2(n_1155),
.B1(n_1107),
.B2(n_1092),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1181),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1094),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1178),
.B(n_1043),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1154),
.A2(n_161),
.B(n_160),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1136),
.B(n_10),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1110),
.A2(n_150),
.B(n_142),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1129),
.A2(n_1139),
.B(n_1204),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1163),
.A2(n_13),
.B(n_15),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1076),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1122),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1104),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1204),
.A2(n_141),
.B(n_136),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1115),
.A2(n_132),
.B(n_128),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1141),
.B(n_1123),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1175),
.B(n_127),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1196),
.B(n_16),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_R g1303 ( 
.A(n_1175),
.B(n_126),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1188),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_22),
.B(n_27),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1111),
.A2(n_124),
.B(n_119),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1180),
.B(n_1162),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1170),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1203),
.A2(n_29),
.A3(n_31),
.B(n_32),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1213),
.B(n_29),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1179),
.B(n_31),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1211),
.A2(n_110),
.B(n_102),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1116),
.A2(n_34),
.B(n_40),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1115),
.A2(n_101),
.B(n_90),
.Y(n_1314)
);

AO22x2_ASAP7_75t_L g1315 ( 
.A1(n_1135),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1124),
.B(n_42),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1146),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.C(n_55),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1202),
.A2(n_46),
.A3(n_53),
.B(n_55),
.Y(n_1318)
);

NAND3x1_ASAP7_75t_L g1319 ( 
.A(n_1157),
.B(n_58),
.C(n_59),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1180),
.B(n_60),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1192),
.B(n_61),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1170),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1154),
.A2(n_76),
.B(n_88),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1193),
.B(n_61),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1132),
.A2(n_75),
.B(n_77),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1176),
.A2(n_89),
.B(n_63),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1202),
.A2(n_1160),
.B(n_1119),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1102),
.B(n_1109),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1132),
.A2(n_1133),
.B(n_1186),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1160),
.A2(n_1101),
.B(n_1113),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1194),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1097),
.A2(n_1152),
.B(n_1177),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1194),
.B(n_1113),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1198),
.A2(n_1169),
.B(n_1151),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1145),
.A2(n_1171),
.B(n_1174),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1205),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1135),
.A2(n_1103),
.B(n_1187),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1150),
.B(n_1167),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1150),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_R g1340 ( 
.A(n_1084),
.B(n_1205),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1167),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1146),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1189),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1189),
.A2(n_1103),
.B(n_1199),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1143),
.A2(n_931),
.B(n_1137),
.C(n_914),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1137),
.B(n_760),
.C(n_756),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1137),
.A2(n_760),
.B(n_756),
.C(n_914),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1112),
.A2(n_632),
.B(n_977),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1137),
.A2(n_931),
.B(n_914),
.C(n_956),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1140),
.B(n_689),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1098),
.A2(n_914),
.B(n_760),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1137),
.A2(n_931),
.B(n_914),
.C(n_956),
.Y(n_1352)
);

AO32x2_ASAP7_75t_L g1353 ( 
.A1(n_1072),
.A2(n_1033),
.A3(n_1203),
.B1(n_1195),
.B2(n_1116),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1183),
.A2(n_1138),
.B(n_1091),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1077),
.Y(n_1355)
);

AO32x2_ASAP7_75t_L g1356 ( 
.A1(n_1072),
.A2(n_1033),
.A3(n_1203),
.B1(n_1195),
.B2(n_1116),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1098),
.B(n_1003),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1148),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1137),
.A2(n_931),
.B(n_914),
.C(n_956),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1072),
.A2(n_956),
.B1(n_615),
.B2(n_599),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1092),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1262),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1269),
.Y(n_1363)
);

AOI22x1_ASAP7_75t_L g1364 ( 
.A1(n_1285),
.A2(n_1337),
.B1(n_1346),
.B2(n_1315),
.Y(n_1364)
);

AOI221x1_ASAP7_75t_L g1365 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_1313),
.B2(n_1349),
.C(n_1352),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1267),
.B(n_1331),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1264),
.B(n_1351),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1220),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1347),
.A2(n_1359),
.B1(n_1222),
.B2(n_1248),
.C(n_1313),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1268),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1345),
.A2(n_1307),
.B1(n_1316),
.B2(n_1357),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1255),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1239),
.A2(n_1329),
.B(n_1348),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1240),
.B(n_1226),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_1217),
.B1(n_1229),
.B2(n_1253),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1293),
.A2(n_1317),
.B1(n_1305),
.B2(n_1315),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1276),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1232),
.A2(n_1291),
.B(n_1236),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1235),
.A2(n_1354),
.B(n_1292),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1253),
.A2(n_1234),
.B1(n_1350),
.B2(n_1243),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1320),
.A2(n_1310),
.B1(n_1321),
.B2(n_1324),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1344),
.B(n_1326),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1301),
.A2(n_1311),
.B1(n_1290),
.B2(n_1355),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1360),
.B(n_1288),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1265),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1294),
.Y(n_1387)
);

AO32x2_ASAP7_75t_L g1388 ( 
.A1(n_1227),
.A2(n_1356),
.A3(n_1353),
.B1(n_1309),
.B2(n_1246),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1221),
.A2(n_1238),
.B(n_1263),
.Y(n_1389)
);

INVx4_ASAP7_75t_SL g1390 ( 
.A(n_1244),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1260),
.B(n_1328),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1271),
.A2(n_1274),
.B(n_1242),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1216),
.B(n_1361),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1293),
.A2(n_1295),
.B(n_1306),
.C(n_1304),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1284),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1287),
.B(n_1286),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1284),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1215),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1275),
.A2(n_1256),
.B(n_1330),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1241),
.A2(n_1237),
.B(n_1299),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1314),
.A2(n_1325),
.B(n_1298),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1332),
.A2(n_1218),
.B(n_1334),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1214),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1218),
.A2(n_1334),
.B(n_1225),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1289),
.A2(n_1323),
.B(n_1327),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1327),
.A2(n_1259),
.B(n_1261),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1278),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1257),
.A2(n_1280),
.B(n_1270),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1259),
.A2(n_1335),
.B(n_1251),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1219),
.A2(n_1319),
.B1(n_1302),
.B2(n_1250),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1333),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1266),
.A2(n_1272),
.B(n_1273),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1296),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1282),
.A2(n_1341),
.B(n_1336),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1340),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_SL g1416 ( 
.A1(n_1343),
.A2(n_1356),
.B(n_1353),
.C(n_1223),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1339),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1338),
.A2(n_1312),
.B(n_1247),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1331),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1258),
.B(n_1219),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1244),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1297),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1300),
.A2(n_1301),
.B1(n_1322),
.B2(n_1308),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1223),
.A2(n_1358),
.B(n_1249),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1353),
.A2(n_1356),
.B(n_1231),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1301),
.B(n_1331),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1318),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1231),
.A2(n_1224),
.B(n_1252),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1318),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1247),
.A2(n_1246),
.B(n_1224),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1214),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1309),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1247),
.A2(n_1246),
.A3(n_1224),
.B(n_1277),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1303),
.B(n_1245),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1267),
.A2(n_1244),
.B(n_1245),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1254),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1267),
.B(n_979),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1220),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1279),
.A2(n_1228),
.B(n_1233),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1346),
.A2(n_1347),
.B(n_1351),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1284),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1283),
.A2(n_1230),
.B(n_1228),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1283),
.A2(n_1230),
.B(n_1228),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1281),
.A2(n_1072),
.B(n_956),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1219),
.B(n_1333),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1331),
.Y(n_1449)
);

CKINVDCx6p67_ASAP7_75t_R g1450 ( 
.A(n_1220),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1220),
.Y(n_1451)
);

INVxp67_ASAP7_75t_SL g1452 ( 
.A(n_1361),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1281),
.A2(n_1072),
.B(n_956),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1240),
.B(n_1172),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1240),
.B(n_1172),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1283),
.A2(n_1230),
.B(n_1228),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1351),
.B(n_1346),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1351),
.B(n_1346),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1346),
.A2(n_1351),
.B1(n_1352),
.B2(n_1349),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1346),
.A2(n_1137),
.B(n_956),
.C(n_1349),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1254),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1254),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1283),
.A2(n_1230),
.B(n_1228),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1346),
.A2(n_1351),
.B1(n_1352),
.B2(n_1349),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1276),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1221),
.A2(n_1165),
.A3(n_1281),
.B(n_1233),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1347),
.A2(n_914),
.B1(n_1351),
.B2(n_756),
.C(n_760),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1254),
.Y(n_1474)
);

INVxp33_ASAP7_75t_L g1475 ( 
.A(n_1240),
.Y(n_1475)
);

CKINVDCx11_ASAP7_75t_R g1476 ( 
.A(n_1220),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1283),
.A2(n_1230),
.B(n_1228),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1219),
.B(n_1333),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1219),
.B(n_1333),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1264),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1264),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1284),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1284),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1357),
.B(n_1226),
.Y(n_1484)
);

AO31x2_ASAP7_75t_L g1485 ( 
.A1(n_1221),
.A2(n_1165),
.A3(n_1281),
.B(n_1233),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1346),
.A2(n_1351),
.B1(n_1352),
.B2(n_1349),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1487)
);

INVx5_ASAP7_75t_L g1488 ( 
.A(n_1244),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1214),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1240),
.B(n_1172),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1253),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_914),
.B2(n_1222),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1222),
.A2(n_914),
.B1(n_1044),
.B2(n_1137),
.Y(n_1495)
);

INVx8_ASAP7_75t_L g1496 ( 
.A(n_1244),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1283),
.A2(n_1228),
.B(n_1233),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1484),
.B(n_1391),
.Y(n_1499)
);

AND2x4_ASAP7_75t_SL g1500 ( 
.A(n_1386),
.B(n_1435),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1473),
.A2(n_1376),
.B1(n_1494),
.B2(n_1492),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1491),
.B(n_1475),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1495),
.A2(n_1463),
.B(n_1459),
.C(n_1458),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1393),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1447),
.B(n_1466),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1376),
.A2(n_1489),
.B1(n_1472),
.B2(n_1447),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1466),
.B(n_1472),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1372),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1494),
.A2(n_1371),
.B1(n_1394),
.B2(n_1369),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1441),
.A2(n_1394),
.B(n_1382),
.C(n_1469),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1480),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1427),
.A2(n_1486),
.B(n_1460),
.Y(n_1515)
);

O2A1O1Ixp5_ASAP7_75t_L g1516 ( 
.A1(n_1383),
.A2(n_1453),
.B(n_1446),
.C(n_1385),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1374),
.A2(n_1364),
.B1(n_1382),
.B2(n_1410),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1421),
.B(n_1381),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1375),
.A2(n_1452),
.B1(n_1377),
.B2(n_1488),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1493),
.B(n_1384),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1479),
.Y(n_1521)
);

OAI22x1_ASAP7_75t_L g1522 ( 
.A1(n_1383),
.A2(n_1433),
.B1(n_1363),
.B2(n_1474),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1479),
.B(n_1367),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1402),
.A2(n_1404),
.B(n_1429),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1377),
.A2(n_1488),
.B1(n_1362),
.B2(n_1437),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1384),
.B(n_1413),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1365),
.A2(n_1366),
.B(n_1420),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1417),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1403),
.B(n_1490),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1377),
.A2(n_1488),
.B1(n_1465),
.B2(n_1467),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1434),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1434),
.B(n_1414),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1366),
.A2(n_1420),
.B(n_1438),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1411),
.B(n_1390),
.Y(n_1534)
);

NOR2xp67_ASAP7_75t_L g1535 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1377),
.A2(n_1488),
.B1(n_1424),
.B2(n_1387),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1481),
.Y(n_1537)
);

NOR2xp67_ASAP7_75t_L g1538 ( 
.A(n_1396),
.B(n_1407),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1396),
.Y(n_1539)
);

AND2x2_ASAP7_75t_SL g1540 ( 
.A(n_1449),
.B(n_1420),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1390),
.B(n_1418),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1415),
.A2(n_1395),
.B1(n_1397),
.B2(n_1482),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1434),
.B(n_1414),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1428),
.Y(n_1544)
);

BUFx4f_ASAP7_75t_L g1545 ( 
.A(n_1378),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1430),
.B(n_1409),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1412),
.B(n_1398),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1412),
.B(n_1378),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1406),
.A2(n_1379),
.B(n_1405),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1409),
.B(n_1378),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1386),
.B(n_1423),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1442),
.A2(n_1483),
.B(n_1416),
.C(n_1395),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1470),
.B(n_1420),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1470),
.B(n_1388),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1470),
.B(n_1388),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1426),
.B(n_1432),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1397),
.A2(n_1482),
.B1(n_1426),
.B2(n_1496),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1388),
.B(n_1425),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1438),
.A2(n_1449),
.B(n_1419),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1426),
.B(n_1431),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1422),
.A2(n_1449),
.B1(n_1423),
.B2(n_1450),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1439),
.A2(n_1451),
.B1(n_1368),
.B2(n_1388),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1406),
.A2(n_1379),
.B(n_1497),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1436),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1476),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1431),
.B(n_1485),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1436),
.B(n_1392),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1408),
.A2(n_1440),
.B(n_1389),
.C(n_1439),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1471),
.B(n_1389),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_L g1570 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1471),
.B(n_1389),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1451),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1471),
.B(n_1399),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1408),
.A2(n_1476),
.B1(n_1400),
.B2(n_1373),
.C(n_1380),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1401),
.B(n_1477),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1576)
);

BUFx4f_ASAP7_75t_SL g1577 ( 
.A(n_1457),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1468),
.B(n_1445),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1454),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1461),
.A2(n_1462),
.B(n_1464),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1487),
.B(n_1455),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1374),
.B(n_1391),
.Y(n_1583)
);

BUFx12f_ASAP7_75t_L g1584 ( 
.A(n_1476),
.Y(n_1584)
);

AOI221x1_ASAP7_75t_SL g1585 ( 
.A1(n_1382),
.A2(n_756),
.B1(n_760),
.B2(n_1351),
.C(n_914),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1393),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1374),
.B(n_1391),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1473),
.A2(n_1072),
.B(n_1248),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1383),
.A2(n_1352),
.B(n_1349),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1393),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1383),
.A2(n_1352),
.B(n_1349),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1383),
.A2(n_1352),
.B(n_1349),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1591),
.A2(n_1594),
.B(n_1593),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1571),
.Y(n_1600)
);

AND2x6_ASAP7_75t_L g1601 ( 
.A(n_1534),
.B(n_1548),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1543),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1544),
.Y(n_1603)
);

BUFx2_ASAP7_75t_SL g1604 ( 
.A(n_1538),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1532),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1590),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1567),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1582),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1532),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1569),
.B(n_1560),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1596),
.B(n_1503),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1560),
.B(n_1566),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1512),
.A2(n_1501),
.B1(n_1508),
.B2(n_1503),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_1562),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1562),
.B(n_1576),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1524),
.Y(n_1618)
);

AO21x2_ASAP7_75t_L g1619 ( 
.A1(n_1568),
.A2(n_1531),
.B(n_1504),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1524),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1563),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1516),
.A2(n_1574),
.B(n_1581),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1578),
.A2(n_1506),
.B(n_1510),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1522),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1550),
.A2(n_1501),
.B(n_1529),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1547),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1587),
.A2(n_1588),
.B(n_1596),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1513),
.A2(n_1512),
.B(n_1508),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1505),
.B(n_1586),
.Y(n_1630)
);

AO21x2_ASAP7_75t_L g1631 ( 
.A1(n_1557),
.A2(n_1509),
.B(n_1506),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1557),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1540),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1592),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1549),
.B(n_1580),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1577),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1509),
.A2(n_1510),
.B(n_1526),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1528),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1525),
.A2(n_1530),
.B(n_1517),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1525),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1515),
.A2(n_1527),
.B(n_1519),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1499),
.B(n_1589),
.Y(n_1643)
);

BUFx12f_ASAP7_75t_L g1644 ( 
.A(n_1565),
.Y(n_1644)
);

AO221x2_ASAP7_75t_L g1645 ( 
.A1(n_1517),
.A2(n_1519),
.B1(n_1585),
.B2(n_1536),
.C(n_1520),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1530),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1539),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1518),
.B(n_1583),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1536),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1502),
.B(n_1507),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1533),
.B(n_1552),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1498),
.B(n_1595),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1602),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1629),
.A2(n_1561),
.B(n_1541),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1599),
.B(n_1521),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1607),
.B(n_1534),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1511),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1599),
.B(n_1523),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1603),
.Y(n_1659)
);

AND2x4_ASAP7_75t_SL g1660 ( 
.A(n_1608),
.B(n_1541),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1603),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1542),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1625),
.B(n_1542),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1601),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1602),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1618),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1610),
.B(n_1553),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1620),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1500),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1597),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1600),
.B(n_1570),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1620),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1621),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1601),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1597),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1600),
.B(n_1572),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1535),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1601),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1605),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1606),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1611),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1644),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1636),
.B(n_1545),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1625),
.B(n_1514),
.Y(n_1686)
);

AOI222xp33_ASAP7_75t_L g1687 ( 
.A1(n_1664),
.A2(n_1629),
.B1(n_1598),
.B2(n_1615),
.C1(n_1642),
.C2(n_1616),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1664),
.A2(n_1598),
.B1(n_1615),
.B2(n_1685),
.C(n_1613),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1658),
.B(n_1650),
.Y(n_1689)
);

OAI33xp33_ASAP7_75t_L g1690 ( 
.A1(n_1685),
.A2(n_1613),
.A3(n_1630),
.B1(n_1647),
.B2(n_1614),
.B3(n_1612),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1677),
.A2(n_1642),
.B1(n_1616),
.B2(n_1647),
.C1(n_1630),
.C2(n_1648),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1678),
.B(n_1628),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1659),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1678),
.B(n_1638),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1627),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1659),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1654),
.A2(n_1670),
.B1(n_1663),
.B2(n_1608),
.C(n_1651),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1663),
.B(n_1633),
.Y(n_1700)
);

INVxp67_ASAP7_75t_SL g1701 ( 
.A(n_1671),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1663),
.B(n_1627),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1653),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1609),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1677),
.A2(n_1648),
.B1(n_1616),
.B2(n_1624),
.C(n_1635),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1686),
.A2(n_1632),
.B(n_1624),
.C(n_1617),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1671),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1658),
.B(n_1672),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1658),
.B(n_1650),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1686),
.A2(n_1645),
.B1(n_1608),
.B2(n_1619),
.Y(n_1715)
);

AOI31xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1681),
.A2(n_1614),
.A3(n_1612),
.B(n_1646),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1683),
.A2(n_1608),
.B1(n_1651),
.B2(n_1633),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1658),
.B(n_1638),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1672),
.A2(n_1645),
.B1(n_1608),
.B2(n_1651),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1656),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1662),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1655),
.B(n_1638),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1608),
.B1(n_1651),
.B2(n_1633),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1645),
.C(n_1638),
.Y(n_1725)
);

OR2x2_ASAP7_75t_SL g1726 ( 
.A(n_1666),
.B(n_1643),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1662),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1665),
.B(n_1609),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1672),
.A2(n_1651),
.B1(n_1632),
.B2(n_1641),
.C(n_1617),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1676),
.B(n_1627),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1645),
.C(n_1638),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1677),
.A2(n_1645),
.B1(n_1619),
.B2(n_1631),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1672),
.B(n_1650),
.Y(n_1734)
);

BUFx10_ASAP7_75t_L g1735 ( 
.A(n_1660),
.Y(n_1735)
);

OAI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1677),
.A2(n_1641),
.B(n_1635),
.C(n_1622),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1676),
.B(n_1623),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1684),
.A2(n_1649),
.B(n_1617),
.C(n_1634),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1675),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1680),
.B(n_1649),
.C(n_1622),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1657),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1662),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1722),
.B(n_1682),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

INVx4_ASAP7_75t_SL g1746 ( 
.A(n_1740),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1742),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1688),
.B(n_1655),
.Y(n_1748)
);

OA21x2_ASAP7_75t_L g1749 ( 
.A1(n_1741),
.A2(n_1673),
.B(n_1669),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1695),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1712),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1698),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1718),
.B(n_1682),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1699),
.A2(n_1651),
.B(n_1619),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1740),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1717),
.A2(n_1619),
.B(n_1640),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1740),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1687),
.A2(n_1660),
.B(n_1637),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1709),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1721),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1728),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1736),
.A2(n_1667),
.B(n_1673),
.Y(n_1764)
);

INVx4_ASAP7_75t_SL g1765 ( 
.A(n_1740),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1714),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1691),
.B(n_1634),
.C(n_1622),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1668),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1743),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1692),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1723),
.Y(n_1771)
);

AND2x6_ASAP7_75t_SL g1772 ( 
.A(n_1692),
.B(n_1584),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1695),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1742),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1703),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1723),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1707),
.B(n_1655),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1727),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1703),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1704),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1704),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1735),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1727),
.Y(n_1784)
);

AND2x4_ASAP7_75t_SL g1785 ( 
.A(n_1735),
.B(n_1656),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1701),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1692),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_SL g1788 ( 
.A(n_1715),
.B(n_1643),
.C(n_1637),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1689),
.B(n_1713),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1710),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1747),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1767),
.A2(n_1715),
.B1(n_1733),
.B2(n_1724),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1773),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1785),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1774),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1745),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1759),
.A2(n_1738),
.B(n_1733),
.C(n_1732),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1772),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1770),
.B(n_1739),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1770),
.B(n_1739),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1786),
.Y(n_1803)
);

NOR3xp33_ASAP7_75t_L g1804 ( 
.A(n_1788),
.B(n_1755),
.C(n_1724),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1786),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1744),
.B(n_1693),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1744),
.B(n_1696),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1753),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1753),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1748),
.B(n_1734),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1777),
.A2(n_1690),
.B1(n_1719),
.B2(n_1725),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_SL g1812 ( 
.A(n_1778),
.B(n_1700),
.C(n_1737),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1790),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1790),
.B(n_1657),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1754),
.B(n_1726),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1789),
.B(n_1668),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1760),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1760),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1762),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1756),
.B(n_1668),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1787),
.B(n_1739),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1757),
.B(n_1716),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1754),
.B(n_1702),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1787),
.A2(n_1700),
.B1(n_1631),
.B2(n_1640),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1763),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1785),
.B(n_1746),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1749),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1769),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1775),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1756),
.B(n_1668),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1757),
.A2(n_1730),
.B(n_1697),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1775),
.B(n_1731),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1780),
.B(n_1626),
.Y(n_1833)
);

NOR3xp33_ASAP7_75t_SL g1834 ( 
.A(n_1780),
.B(n_1537),
.C(n_1781),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1781),
.B(n_1626),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1809),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1809),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1810),
.B(n_1782),
.Y(n_1838)
);

NAND2x1p5_ASAP7_75t_L g1839 ( 
.A(n_1822),
.B(n_1783),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_SL g1840 ( 
.A1(n_1798),
.A2(n_1758),
.B(n_1751),
.C(n_1782),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1814),
.B(n_1758),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1797),
.Y(n_1842)
);

INVxp33_ASAP7_75t_SL g1843 ( 
.A(n_1800),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1801),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1801),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1821),
.B(n_1746),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1811),
.B(n_1750),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1799),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1803),
.B(n_1750),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1808),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1817),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1826),
.B(n_1746),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1821),
.B(n_1746),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1794),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1818),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1805),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1813),
.B(n_1752),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1819),
.B(n_1752),
.Y(n_1858)
);

AND3x2_ASAP7_75t_L g1859 ( 
.A(n_1826),
.B(n_1765),
.C(n_1639),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1793),
.A2(n_1764),
.B1(n_1604),
.B2(n_1749),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1802),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1802),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1825),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1828),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1792),
.B(n_1768),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1816),
.B(n_1631),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_SL g1867 ( 
.A(n_1796),
.B(n_1644),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1829),
.B(n_1761),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1815),
.B(n_1631),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1832),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1798),
.B(n_1761),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1832),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1831),
.A2(n_1783),
.B(n_1675),
.C(n_1679),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1820),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1795),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1843),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1853),
.B(n_1852),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1836),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1854),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1837),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1852),
.B(n_1795),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1861),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1839),
.A2(n_1824),
.B1(n_1804),
.B2(n_1834),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1839),
.B(n_1765),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1862),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1842),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1867),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1856),
.B(n_1806),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1870),
.B(n_1806),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1848),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1859),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1844),
.B(n_1765),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1847),
.A2(n_1812),
.B1(n_1764),
.B2(n_1815),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1845),
.B(n_1765),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1872),
.Y(n_1895)
);

NOR2x1_ASAP7_75t_L g1896 ( 
.A(n_1860),
.B(n_1791),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1850),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1873),
.B(n_1783),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1865),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1838),
.B(n_1823),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.B(n_1823),
.Y(n_1901)
);

INVx4_ASAP7_75t_L g1902 ( 
.A(n_1863),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1851),
.Y(n_1903)
);

NAND3xp33_ASAP7_75t_L g1904 ( 
.A(n_1896),
.B(n_1840),
.C(n_1860),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1879),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1876),
.B(n_1644),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1876),
.B(n_1864),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1878),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1878),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1883),
.A2(n_1847),
.B1(n_1871),
.B2(n_1874),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1880),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1885),
.B(n_1871),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1885),
.B(n_1855),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1880),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1895),
.Y(n_1915)
);

OAI211xp5_ASAP7_75t_L g1916 ( 
.A1(n_1896),
.A2(n_1869),
.B(n_1849),
.C(n_1857),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1887),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1877),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1881),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1893),
.A2(n_1857),
.B1(n_1858),
.B2(n_1791),
.C(n_1827),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1883),
.A2(n_1764),
.B1(n_1749),
.B2(n_1640),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1887),
.A2(n_1858),
.B(n_1868),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1895),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1885),
.B(n_1841),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1895),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1899),
.B(n_1830),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1891),
.B(n_1783),
.Y(n_1927)
);

NOR2xp67_ASAP7_75t_L g1928 ( 
.A(n_1904),
.B(n_1882),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1906),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1917),
.B(n_1899),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1915),
.Y(n_1931)
);

AND2x4_ASAP7_75t_SL g1932 ( 
.A(n_1906),
.B(n_1877),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1923),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1919),
.B(n_1875),
.Y(n_1934)
);

NAND2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1927),
.B(n_1884),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1907),
.B(n_1875),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1918),
.B(n_1881),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1919),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1905),
.B(n_1881),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1925),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_SL g1941 ( 
.A(n_1912),
.B(n_1891),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1910),
.B(n_1881),
.Y(n_1942)
);

AOI321xp33_ASAP7_75t_L g1943 ( 
.A1(n_1942),
.A2(n_1920),
.A3(n_1927),
.B1(n_1916),
.B2(n_1921),
.C(n_1922),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1941),
.B(n_1884),
.Y(n_1944)
);

NOR2x1_ASAP7_75t_L g1945 ( 
.A(n_1930),
.B(n_1902),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1928),
.B(n_1924),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1941),
.A2(n_1921),
.B(n_1913),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1936),
.A2(n_1898),
.B1(n_1892),
.B2(n_1894),
.Y(n_1948)
);

O2A1O1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1935),
.A2(n_1909),
.B(n_1911),
.C(n_1914),
.Y(n_1949)
);

NOR3xp33_ASAP7_75t_L g1950 ( 
.A(n_1929),
.B(n_1908),
.C(n_1902),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1934),
.A2(n_1888),
.B(n_1926),
.Y(n_1951)
);

AOI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1939),
.A2(n_1902),
.B1(n_1888),
.B2(n_1886),
.C(n_1903),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_SL g1953 ( 
.A1(n_1938),
.A2(n_1903),
.B(n_1890),
.C(n_1897),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1953),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1949),
.Y(n_1955)
);

O2A1O1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1944),
.A2(n_1935),
.B(n_1940),
.C(n_1933),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1947),
.A2(n_1932),
.B(n_1937),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1945),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1946),
.B(n_1931),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1948),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_SL g1961 ( 
.A(n_1954),
.B(n_1902),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_L g1962 ( 
.A(n_1958),
.B(n_1950),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1955),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1959),
.Y(n_1964)
);

OAI21xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1960),
.A2(n_1952),
.B(n_1943),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1956),
.Y(n_1966)
);

NOR2x1_ASAP7_75t_L g1967 ( 
.A(n_1957),
.B(n_1951),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1960),
.B(n_1898),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1967),
.A2(n_1901),
.B1(n_1889),
.B2(n_1900),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1965),
.A2(n_1892),
.B1(n_1894),
.B2(n_1897),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1966),
.B(n_1968),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1963),
.B(n_1886),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1964),
.A2(n_1901),
.B1(n_1889),
.B2(n_1900),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1962),
.B(n_1890),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_SL g1975 ( 
.A1(n_1970),
.A2(n_1961),
.B(n_1868),
.Y(n_1975)
);

AOI221xp5_ASAP7_75t_L g1976 ( 
.A1(n_1969),
.A2(n_1961),
.B1(n_1827),
.B2(n_1783),
.C(n_1833),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1974),
.B(n_1807),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1972),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1978),
.B(n_1971),
.Y(n_1979)
);

NOR3xp33_ASAP7_75t_SL g1980 ( 
.A(n_1975),
.B(n_1973),
.C(n_1604),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1979),
.A2(n_1977),
.B1(n_1976),
.B2(n_1764),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1980),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1982),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1981),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1983),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_L g1986 ( 
.A(n_1984),
.B(n_1835),
.C(n_1833),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1985),
.A2(n_1866),
.B1(n_1835),
.B2(n_1807),
.Y(n_1987)
);

AOI22x1_ASAP7_75t_L g1988 ( 
.A1(n_1986),
.A2(n_1784),
.B1(n_1779),
.B2(n_1776),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1988),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1989),
.A2(n_1987),
.B1(n_1784),
.B2(n_1779),
.C(n_1776),
.Y(n_1990)
);

AOI222xp33_ASAP7_75t_L g1991 ( 
.A1(n_1990),
.A2(n_1771),
.B1(n_1766),
.B2(n_1768),
.C1(n_1639),
.C2(n_1711),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_SL g1992 ( 
.A1(n_1991),
.A2(n_1771),
.B1(n_1766),
.B2(n_1705),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1992),
.A2(n_1705),
.B1(n_1706),
.B2(n_1729),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_L g1994 ( 
.A1(n_1993),
.A2(n_1652),
.B(n_1684),
.C(n_1729),
.Y(n_1994)
);


endmodule