module fake_jpeg_7595_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_30),
.B1(n_24),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_47),
.B1(n_22),
.B2(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_30),
.B1(n_15),
.B2(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_15),
.B1(n_17),
.B2(n_28),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_66),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_76),
.Y(n_82)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_77),
.B1(n_27),
.B2(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_60),
.B1(n_51),
.B2(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_92),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_90),
.B1(n_100),
.B2(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_59),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_2),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_50),
.B1(n_26),
.B2(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_80),
.B1(n_63),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_95),
.B1(n_81),
.B2(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_64),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_115),
.C(n_13),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_70),
.B1(n_46),
.B2(n_66),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_67),
.C(n_53),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_119),
.C(n_81),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_117),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_25),
.C(n_31),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_128),
.Y(n_151)
);

NOR4xp25_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_85),
.C(n_84),
.D(n_93),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_127),
.C(n_115),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_105),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_105),
.C(n_111),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_67),
.B(n_35),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_119),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_35),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_103),
.C(n_107),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_70),
.C(n_25),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_14),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_89),
.B(n_86),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_103),
.C(n_113),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_146),
.B1(n_124),
.B2(n_35),
.C(n_13),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_115),
.C(n_108),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_149),
.C(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_132),
.C(n_125),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_131),
.B1(n_133),
.B2(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_159),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_124),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_163),
.Y(n_165)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_57),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_3),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_144),
.B1(n_140),
.B2(n_141),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_55),
.B(n_4),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_159),
.A2(n_3),
.B(n_4),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_152),
.C(n_157),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_3),
.B(n_4),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_5),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_173),
.C(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_165),
.Y(n_182)
);

AOI31xp33_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_161),
.A3(n_152),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

OAI211xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_6),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_185),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_177),
.B1(n_55),
.B2(n_7),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_180),
.B(n_6),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_190),
.B(n_186),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_191),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_193),
.Y(n_194)
);


endmodule