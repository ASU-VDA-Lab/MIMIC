module fake_aes_7593_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_SL g3 ( .A(n_2), .B(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_5), .B(n_2), .Y(n_6) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_5), .Y(n_8) );
OAI211xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_4), .B(n_1), .C(n_2), .Y(n_9) );
AOI22xp5_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_10) );
AO22x1_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_8), .B1(n_9), .B2(n_0), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B1(n_9), .B2(n_2), .Y(n_15) );
endmodule