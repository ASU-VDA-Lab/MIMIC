module fake_jpeg_25753_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_18),
.B1(n_21),
.B2(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_24),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_22),
.Y(n_35)
);

NOR2xp67_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_33),
.B(n_26),
.Y(n_38)
);


endmodule