module real_jpeg_23376_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_35),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_1),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_153),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_3),
.A2(n_69),
.B1(n_153),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_67),
.B1(n_70),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_113),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_113),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_162),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_6),
.A2(n_77),
.B1(n_162),
.B2(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_52),
.B1(n_67),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_9),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_68),
.B1(n_85),
.B2(n_124),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_85),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_11),
.A2(n_28),
.B(n_43),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_11),
.B(n_91),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_25),
.B1(n_32),
.B2(n_180),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_62),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_11),
.B(n_78),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_139),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_20),
.B(n_118),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_100),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_21),
.A2(n_80),
.B1(n_81),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_21),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_53),
.B2(n_79),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_22),
.A2(n_54),
.B(n_56),
.Y(n_137)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_24),
.A2(n_36),
.B1(n_54),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_25),
.A2(n_106),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_25),
.A2(n_108),
.B1(n_170),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_25),
.A2(n_33),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_25),
.A2(n_206),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_26),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_26),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_27),
.B(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_32),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_34),
.B(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_36),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_47),
.B(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_37),
.A2(n_46),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_37),
.A2(n_94),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_38),
.A2(n_95),
.B(n_96),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_38),
.A2(n_96),
.B1(n_152),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_38),
.A2(n_96),
.B1(n_161),
.B2(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_38),
.A2(n_50),
.B(n_95),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_41),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_40),
.B(n_89),
.Y(n_204)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_41),
.A2(n_45),
.B(n_150),
.C(n_155),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_41),
.A2(n_62),
.A3(n_88),
.B1(n_195),
.B2(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_46),
.B(n_150),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_46),
.A2(n_97),
.B(n_110),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_71),
.B(n_75),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_57),
.A2(n_58),
.B1(n_112),
.B2(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_70),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_59),
.A2(n_63),
.A3(n_69),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_60),
.B(n_62),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_63),
.B(n_150),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_70),
.A2(n_150),
.B(n_241),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_78),
.Y(n_114)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_73),
.B(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_77),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_78),
.A2(n_126),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_78),
.A2(n_126),
.B1(n_259),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_93),
.B(n_99),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_93),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_87),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_92),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_86),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_86),
.A2(n_91),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_86),
.A2(n_91),
.B1(n_220),
.B2(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_86),
.A2(n_255),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_87),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_87),
.B(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_117),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_120),
.B1(n_135),
.B2(n_136),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_100),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.C(n_115),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_101),
.A2(n_102),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_103),
.B(n_109),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_104),
.A2(n_173),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_105),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_111),
.B(n_115),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_137),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_134),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_132),
.A2(n_196),
.B(n_271),
.Y(n_289)
);

AOI311xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_301),
.A3(n_313),
.B(n_317),
.C(n_318),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_262),
.C(n_296),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_235),
.B(n_261),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_213),
.B(n_234),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_188),
.B(n_212),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_166),
.B(n_187),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_148),
.B1(n_154),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_163),
.C(n_164),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_165),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_176),
.B(n_186),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_174),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_185),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_202),
.B1(n_210),
.B2(n_211),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.C(n_210),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_205),
.Y(n_229)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_227),
.B2(n_228),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_230),
.C(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_223),
.C(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_252),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_251),
.C(n_252),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_263),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_264),
.B(n_281),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_276),
.C(n_277),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_265),
.A2(n_266),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_269),
.C(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_277),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_291),
.B2(n_292),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_292),
.C(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_290),
.Y(n_284)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_314),
.B(n_319),
.C(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_310),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.C(n_309),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_307),
.CI(n_309),
.CON(n_316),
.SN(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_316),
.Y(n_324)
);


endmodule