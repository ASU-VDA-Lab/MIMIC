module fake_jpeg_17836_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_2),
.Y(n_72)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_41),
.B1(n_53),
.B2(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_57),
.B1(n_49),
.B2(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_79),
.B1(n_80),
.B2(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_3),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_57),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_51),
.B1(n_45),
.B2(n_41),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_40),
.B(n_6),
.C(n_7),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_42),
.B1(n_51),
.B2(n_5),
.Y(n_79)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_98),
.B1(n_9),
.B2(n_10),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_4),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_91),
.B(n_93),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_52),
.B(n_50),
.C(n_44),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_89),
.C(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_4),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_99),
.B(n_9),
.C(n_14),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_86),
.B(n_88),
.C(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_18),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_87),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_106),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_101),
.C(n_107),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_87),
.B(n_20),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_105),
.B1(n_96),
.B2(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_119),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_130),
.B1(n_125),
.B2(n_21),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_129),
.C(n_131),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_19),
.C(n_22),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_23),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_24),
.B(n_25),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_26),
.B(n_30),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_37),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_31),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_35),
.Y(n_142)
);


endmodule