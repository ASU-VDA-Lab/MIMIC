module fake_ibex_304_n_1499 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1499);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1499;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1421;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_1115;
wire n_998;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1361;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_74),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_15),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_157),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_144),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_13),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_161),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_189),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_150),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_260),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_43),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_58),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_188),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_124),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_57),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_89),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_169),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_230),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_175),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_168),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_156),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_266),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g305 ( 
.A(n_248),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_252),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_193),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_71),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_179),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_245),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_126),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_267),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_121),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_198),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_93),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_159),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_208),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_180),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_239),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_187),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_214),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_53),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_241),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_31),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_203),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_99),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_64),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_145),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_17),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_74),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_23),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_213),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_35),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_128),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_268),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_71),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_3),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_197),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_192),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_215),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_224),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_123),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_221),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_243),
.B(n_44),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_54),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_134),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_153),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_51),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_132),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_250),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_100),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_49),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_19),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_13),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_100),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_227),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_42),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_51),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_185),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_226),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_151),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_242),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_235),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_256),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_2),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_207),
.B(n_56),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_65),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_212),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_190),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_238),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_124),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_135),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_24),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_33),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_86),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_123),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_135),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_43),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_113),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_85),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_165),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_58),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_132),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_82),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_70),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_69),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_2),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_184),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_158),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_155),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_33),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_56),
.B(n_173),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_255),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_247),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_183),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_233),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_234),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_205),
.Y(n_413)
);

BUFx2_ASAP7_75t_SL g414 ( 
.A(n_37),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_194),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_170),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_237),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_7),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_116),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_167),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_178),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_62),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_254),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_219),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_160),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_139),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_81),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_164),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_196),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_228),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_17),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_209),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_77),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_50),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_49),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_166),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_114),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_69),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_103),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_61),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_62),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_206),
.B(n_191),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_4),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_119),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_5),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_6),
.B(n_120),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_47),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_218),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_65),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_116),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_96),
.B(n_176),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_59),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_120),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_29),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_232),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_107),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_103),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_77),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_60),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_174),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_24),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_154),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_259),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_73),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_118),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_202),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_220),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_57),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_133),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_98),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_16),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_142),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_75),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_36),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_133),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_114),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_95),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_8),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_35),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_334),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_403),
.Y(n_482)
);

BUFx12f_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_295),
.B(n_0),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_354),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_273),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_354),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_334),
.B(n_1),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_368),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_368),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_332),
.B(n_4),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_362),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_394),
.B(n_363),
.Y(n_497)
);

INVx6_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_299),
.B(n_309),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_273),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_324),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_294),
.B(n_9),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_365),
.B(n_9),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_276),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_427),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_276),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_286),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_480),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_435),
.B(n_10),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_395),
.B(n_463),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_388),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_480),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_388),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_442),
.B(n_11),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_286),
.A2(n_146),
.B(n_143),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_293),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_293),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_290),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_446),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_284),
.B(n_14),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_350),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_318),
.B(n_16),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_379),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_296),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_322),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_375),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_275),
.B(n_21),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_350),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_360),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_360),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_383),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_327),
.B(n_22),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_471),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_409),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_422),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_308),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_471),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_289),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_479),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_308),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_555)
);

BUFx8_ASAP7_75t_L g556 ( 
.A(n_452),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_344),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_344),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_422),
.B(n_460),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_409),
.B(n_25),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_313),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_269),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_344),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_379),
.A2(n_316),
.B1(n_359),
.B2(n_313),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_362),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_316),
.B(n_28),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_270),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_431),
.B(n_29),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_402),
.A2(n_148),
.B(n_147),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_402),
.Y(n_572)
);

OA21x2_ASAP7_75t_L g573 ( 
.A1(n_408),
.A2(n_152),
.B(n_149),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_310),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_344),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_271),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_L g580 ( 
.A(n_511),
.B(n_459),
.C(n_423),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_498),
.B(n_420),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_498),
.B(n_420),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_498),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_498),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_536),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_490),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_536),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_482),
.B(n_278),
.Y(n_591)
);

CKINVDCx6p67_ASAP7_75t_R g592 ( 
.A(n_519),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_482),
.B(n_282),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_525),
.Y(n_595)
);

BUFx6f_ASAP7_75t_SL g596 ( 
.A(n_505),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_537),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_497),
.B(n_423),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_490),
.Y(n_600)
);

AND3x2_ASAP7_75t_L g601 ( 
.A(n_499),
.B(n_425),
.C(n_370),
.Y(n_601)
);

CKINVDCx11_ASAP7_75t_R g602 ( 
.A(n_567),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_548),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_428),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_520),
.B(n_428),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_556),
.B(n_282),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_548),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_521),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_520),
.B(n_432),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_510),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_505),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_525),
.B(n_432),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_564),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_556),
.B(n_283),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_559),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_564),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_567),
.B(n_552),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_526),
.B(n_355),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_519),
.B(n_414),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_488),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_488),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_575),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_559),
.B(n_285),
.Y(n_627)
);

CKINVDCx6p67_ASAP7_75t_R g628 ( 
.A(n_483),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_575),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_575),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_575),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_485),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_553),
.A2(n_287),
.B1(n_288),
.B2(n_280),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_560),
.B(n_418),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_510),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

AOI22x1_ASAP7_75t_L g637 ( 
.A1(n_512),
.A2(n_411),
.B1(n_279),
.B2(n_281),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_539),
.B(n_289),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_514),
.B(n_277),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_514),
.B(n_285),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_512),
.Y(n_641)
);

BUFx6f_ASAP7_75t_SL g642 ( 
.A(n_561),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_553),
.B(n_516),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_483),
.B(n_516),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_578),
.Y(n_645)
);

BUFx6f_ASAP7_75t_SL g646 ( 
.A(n_561),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_578),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_485),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_566),
.A2(n_440),
.B1(n_441),
.B2(n_438),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_570),
.B(n_291),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_513),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_485),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_513),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_539),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_533),
.A2(n_440),
.B1(n_441),
.B2(n_438),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_550),
.A2(n_453),
.B1(n_457),
.B2(n_451),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_570),
.B(n_291),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_492),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_570),
.B(n_298),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_492),
.Y(n_661)
);

CKINVDCx11_ASAP7_75t_R g662 ( 
.A(n_523),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_563),
.B(n_298),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_504),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_527),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_568),
.A2(n_311),
.B1(n_330),
.B2(n_292),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_492),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_569),
.B(n_451),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_447),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_568),
.B(n_453),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_579),
.B(n_457),
.Y(n_672)
);

AND3x2_ASAP7_75t_L g673 ( 
.A(n_515),
.B(n_467),
.C(n_331),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_SL g674 ( 
.A(n_515),
.B(n_302),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_576),
.B(n_304),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_501),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_530),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_576),
.B(n_304),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_576),
.B(n_306),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_501),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_538),
.B(n_475),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_549),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_502),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_573),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_549),
.B(n_306),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_297),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_532),
.B(n_300),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_484),
.A2(n_475),
.B1(n_323),
.B2(n_378),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_543),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_549),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_524),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_538),
.B(n_551),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_495),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_545),
.B(n_312),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_517),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_524),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_551),
.B(n_315),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_486),
.B(n_301),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_572),
.B(n_315),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_507),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_486),
.B(n_303),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_489),
.B(n_491),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_524),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_517),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_572),
.B(n_356),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_524),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_524),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_574),
.B(n_356),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_496),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_660),
.B(n_424),
.Y(n_714)
);

AO22x2_ASAP7_75t_L g715 ( 
.A1(n_580),
.A2(n_555),
.B1(n_562),
.B2(n_535),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_671),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_708),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_681),
.B(n_426),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_589),
.A2(n_571),
.B(n_522),
.C(n_493),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_581),
.A2(n_493),
.B1(n_494),
.B2(n_491),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_619),
.B(n_429),
.Y(n_721)
);

BUFx8_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_671),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_634),
.B(n_429),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_582),
.B(n_583),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_591),
.B(n_494),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_643),
.A2(n_481),
.B1(n_323),
.B2(n_378),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_599),
.A2(n_571),
.B(n_506),
.C(n_508),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_595),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_623),
.B(n_302),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_672),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_704),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_712),
.B(n_274),
.C(n_272),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_594),
.B(n_500),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_598),
.A2(n_417),
.B1(n_433),
.B2(n_410),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_704),
.B(n_430),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_697),
.B(n_468),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_636),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_L g742 ( 
.A1(n_600),
.A2(n_340),
.B(n_337),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_640),
.B(n_500),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_706),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_604),
.B(n_338),
.Y(n_745)
);

AND2x6_ASAP7_75t_SL g746 ( 
.A(n_602),
.B(n_341),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_624),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_623),
.B(n_410),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_669),
.B(n_506),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_607),
.B(n_508),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_625),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_509),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_581),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_639),
.B(n_509),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_581),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_654),
.B(n_528),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_664),
.B(n_528),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_650),
.B(n_540),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_656),
.B(n_540),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_687),
.B(n_688),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_657),
.B(n_542),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_712),
.B(n_348),
.C(n_345),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_655),
.A2(n_554),
.B(n_547),
.C(n_347),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_615),
.B(n_366),
.C(n_358),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_592),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

NAND2x1_ASAP7_75t_L g767 ( 
.A(n_614),
.B(n_616),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_611),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_649),
.B(n_638),
.C(n_674),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_611),
.A2(n_361),
.B1(n_364),
.B2(n_342),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

NOR2x1p5_ASAP7_75t_L g772 ( 
.A(n_592),
.B(n_371),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_701),
.B(n_622),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_628),
.B(n_372),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_305),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_606),
.A2(n_387),
.B1(n_389),
.B2(n_367),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_628),
.B(n_390),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_307),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_698),
.B(n_314),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_588),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_638),
.B(n_398),
.C(n_393),
.Y(n_781)
);

AOI221xp5_ASAP7_75t_L g782 ( 
.A1(n_633),
.A2(n_391),
.B1(n_401),
.B2(n_399),
.C(n_396),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_616),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_667),
.A2(n_461),
.B1(n_473),
.B2(n_433),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_584),
.B(n_335),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_584),
.B(n_349),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_623),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_605),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_461),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_677),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_665),
.B(n_400),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_703),
.B(n_317),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_585),
.B(n_352),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_602),
.B(n_404),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_644),
.A2(n_473),
.B1(n_462),
.B2(n_465),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_609),
.B(n_382),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_709),
.B(n_319),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_618),
.B(n_412),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_613),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_596),
.A2(n_466),
.B1(n_472),
.B2(n_406),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_678),
.B(n_419),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_627),
.B(n_320),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_674),
.B(n_477),
.C(n_436),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_596),
.B(n_321),
.Y(n_804)
);

INVx8_ASAP7_75t_L g805 ( 
.A(n_642),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_642),
.B(n_325),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_635),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_663),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_670),
.B(n_416),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_670),
.B(n_326),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_670),
.B(n_328),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_679),
.B(n_329),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_686),
.B(n_333),
.Y(n_813)
);

NOR2xp67_ASAP7_75t_L g814 ( 
.A(n_690),
.B(n_557),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_686),
.B(n_336),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_673),
.Y(n_816)
);

NOR3xp33_ASAP7_75t_L g817 ( 
.A(n_662),
.B(n_444),
.C(n_434),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_685),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_635),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_641),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_646),
.B(n_339),
.Y(n_821)
);

BUFx6f_ASAP7_75t_SL g822 ( 
.A(n_641),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_651),
.B(n_653),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_653),
.B(n_343),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_637),
.A2(n_448),
.B1(n_450),
.B2(n_445),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_662),
.B(n_455),
.C(n_454),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_637),
.A2(n_469),
.B1(n_474),
.B2(n_458),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_689),
.B(n_385),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_646),
.A2(n_476),
.B1(n_392),
.B2(n_439),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_689),
.B(n_346),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_691),
.A2(n_696),
.B1(n_693),
.B2(n_666),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_691),
.B(n_351),
.Y(n_832)
);

AO221x1_ASAP7_75t_L g833 ( 
.A1(n_621),
.A2(n_392),
.B1(n_397),
.B2(n_439),
.C(n_478),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_693),
.B(n_353),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_601),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_702),
.B(n_369),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_705),
.B(n_373),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_692),
.B(n_374),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_683),
.B(n_357),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_621),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_708),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_713),
.A2(n_397),
.B1(n_380),
.B2(n_376),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_377),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_708),
.B(n_384),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_586),
.B(n_407),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_L g846 ( 
.A1(n_713),
.A2(n_478),
.B1(n_415),
.B2(n_421),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_587),
.A2(n_573),
.B(n_590),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_590),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_593),
.B(n_443),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_593),
.A2(n_478),
.B1(n_449),
.B2(n_456),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_808),
.B(n_30),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_799),
.A2(n_464),
.B1(n_558),
.B2(n_557),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_799),
.Y(n_853)
);

BUFx2_ASAP7_75t_SL g854 ( 
.A(n_822),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_733),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_722),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_828),
.B(n_31),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_725),
.A2(n_565),
.B(n_577),
.C(n_558),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_741),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_716),
.B(n_32),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_717),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_831),
.A2(n_577),
.B1(n_603),
.B2(n_597),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_806),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_773),
.A2(n_610),
.B(n_608),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_744),
.B(n_32),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_726),
.A2(n_620),
.B(n_617),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_760),
.A2(n_629),
.B(n_626),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_722),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_34),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_725),
.B(n_34),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_783),
.A2(n_767),
.B(n_847),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_787),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_754),
.A2(n_630),
.B(n_631),
.C(n_629),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_806),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_732),
.B(n_36),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_738),
.B(n_38),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_714),
.B(n_38),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_723),
.B(n_39),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_730),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_758),
.A2(n_761),
.B(n_757),
.C(n_755),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_723),
.B(n_39),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_763),
.A2(n_647),
.B(n_645),
.C(n_648),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_846),
.A2(n_661),
.B(n_668),
.C(n_658),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_766),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_753),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_739),
.B(n_40),
.Y(n_887)
);

AND2x2_ASAP7_75t_SL g888 ( 
.A(n_731),
.B(n_41),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_745),
.B(n_45),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_761),
.A2(n_531),
.B(n_534),
.C(n_707),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_769),
.A2(n_531),
.B1(n_534),
.B2(n_699),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_765),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_759),
.B(n_46),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_750),
.B(n_752),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_784),
.B(n_680),
.C(n_676),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_846),
.A2(n_711),
.B(n_700),
.C(n_694),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_737),
.B(n_46),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_771),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_728),
.B(n_682),
.C(n_680),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_823),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_813),
.A2(n_815),
.B(n_838),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_770),
.B(n_47),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_829),
.B(n_48),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_770),
.B(n_48),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_838),
.A2(n_749),
.B(n_740),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_778),
.B(n_50),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_778),
.B(n_776),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_805),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_776),
.B(n_52),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_802),
.B(n_53),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_751),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_734),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_731),
.B(n_748),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_720),
.A2(n_825),
.B1(n_827),
.B2(n_769),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_791),
.B(n_789),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_802),
.B(n_54),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_805),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_774),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_748),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_801),
.B(n_55),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_816),
.B(n_55),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_841),
.A2(n_652),
.B(n_632),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_720),
.A2(n_827),
.B1(n_825),
.B2(n_780),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_801),
.B(n_60),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_822),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_757),
.A2(n_710),
.B(n_684),
.C(n_64),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_775),
.B(n_61),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_727),
.B(n_63),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_800),
.B(n_63),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_804),
.B(n_66),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_727),
.B(n_66),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_728),
.B(n_67),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_789),
.B(n_67),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_804),
.A2(n_182),
.B(n_263),
.C(n_262),
.Y(n_936)
);

CKINVDCx10_ASAP7_75t_R g937 ( 
.A(n_746),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_788),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_756),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_809),
.B(n_68),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_736),
.B(n_70),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_736),
.B(n_72),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_743),
.B(n_72),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_806),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_743),
.B(n_73),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_794),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_724),
.A2(n_75),
.B(n_76),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_807),
.A2(n_820),
.B(n_819),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_790),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_735),
.A2(n_762),
.B(n_779),
.Y(n_950)
);

OA22x2_ASAP7_75t_L g951 ( 
.A1(n_833),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_777),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_772),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_803),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_803),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_821),
.B(n_835),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_814),
.B(n_83),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_781),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_818),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_845),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_812),
.B(n_84),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_781),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_795),
.B(n_842),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_742),
.A2(n_87),
.B(n_88),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_779),
.B(n_89),
.Y(n_965)
);

OAI321xp33_ASAP7_75t_L g966 ( 
.A1(n_810),
.A2(n_90),
.A3(n_91),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_824),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_792),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_817),
.B(n_97),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_830),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_832),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_792),
.B(n_797),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_797),
.B(n_98),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_715),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_821),
.A2(n_101),
.B(n_102),
.C(n_104),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_764),
.B(n_105),
.Y(n_976)
);

AND2x6_ASAP7_75t_L g977 ( 
.A(n_818),
.B(n_171),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_836),
.A2(n_837),
.B(n_844),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_796),
.B(n_106),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_811),
.B(n_106),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_782),
.B(n_107),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_817),
.B(n_108),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_834),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_826),
.B(n_109),
.C(n_110),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_826),
.A2(n_111),
.B(n_112),
.C(n_113),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_843),
.B(n_111),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_798),
.B(n_112),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_721),
.B(n_115),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_715),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_715),
.B(n_121),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_839),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_849),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_849),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_850),
.A2(n_122),
.B(n_125),
.C(n_126),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_785),
.B(n_125),
.Y(n_995)
);

CKINVDCx11_ASAP7_75t_R g996 ( 
.A(n_840),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_786),
.B(n_127),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_919),
.B(n_793),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_888),
.B(n_129),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_895),
.A2(n_848),
.B1(n_131),
.B2(n_134),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_869),
.Y(n_1001)
);

AND2x6_ASAP7_75t_L g1002 ( 
.A(n_864),
.B(n_848),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_881),
.A2(n_848),
.B(n_131),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_862),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_917),
.A2(n_130),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_920),
.B(n_136),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_855),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_868),
.A2(n_137),
.A3(n_138),
.B(n_139),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_948),
.A2(n_140),
.B(n_141),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_140),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_902),
.A2(n_907),
.B(n_925),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_919),
.B(n_265),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_963),
.B(n_217),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_910),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_SL g1015 ( 
.A1(n_944),
.A2(n_229),
.B(n_231),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_865),
.A2(n_924),
.B(n_867),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_925),
.A2(n_240),
.B(n_874),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_SL g1018 ( 
.A1(n_856),
.A2(n_946),
.B1(n_920),
.B2(n_990),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_SL g1019 ( 
.A(n_873),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_910),
.B(n_880),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_952),
.B(n_898),
.Y(n_1021)
);

O2A1O1Ixp5_ASAP7_75t_L g1022 ( 
.A1(n_932),
.A2(n_986),
.B(n_956),
.C(n_912),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_904),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_990),
.A2(n_916),
.B1(n_971),
.B2(n_970),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_913),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_916),
.B(n_914),
.Y(n_1026)
);

AOI211x1_ASAP7_75t_L g1027 ( 
.A1(n_981),
.A2(n_931),
.B(n_911),
.C(n_906),
.Y(n_1027)
);

AOI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_958),
.A2(n_892),
.B(n_954),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_883),
.A2(n_882),
.B(n_879),
.C(n_890),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_866),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_878),
.A2(n_965),
.B(n_973),
.C(n_870),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_929),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_921),
.A2(n_935),
.B1(n_929),
.B2(n_915),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_918),
.A2(n_908),
.B(n_945),
.C(n_943),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_959),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_893),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_871),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_996),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_860),
.B(n_857),
.Y(n_1039)
);

OA22x2_ASAP7_75t_L g1040 ( 
.A1(n_990),
.A2(n_989),
.B1(n_974),
.B2(n_957),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_886),
.B(n_889),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_984),
.B(n_985),
.C(n_962),
.Y(n_1042)
);

CKINVDCx11_ASAP7_75t_R g1043 ( 
.A(n_937),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_851),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_899),
.B(n_922),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_926),
.B(n_950),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_960),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_950),
.B(n_877),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_887),
.B(n_934),
.Y(n_1049)
);

AND3x4_ASAP7_75t_L g1050 ( 
.A(n_957),
.B(n_923),
.C(n_979),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_936),
.A2(n_891),
.B(n_928),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_927),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_900),
.B(n_947),
.C(n_987),
.Y(n_1053)
);

NOR2x1_ASAP7_75t_L g1054 ( 
.A(n_905),
.B(n_976),
.Y(n_1054)
);

AOI221x1_ASAP7_75t_L g1055 ( 
.A1(n_964),
.A2(n_975),
.B1(n_967),
.B2(n_983),
.C(n_968),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_876),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_997),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_980),
.B(n_903),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_930),
.A2(n_941),
.B1(n_942),
.B2(n_933),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_858),
.A2(n_940),
.B(n_994),
.C(n_884),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_955),
.A2(n_983),
.B1(n_967),
.B2(n_894),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_979),
.B(n_982),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_897),
.A2(n_852),
.B(n_863),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_991),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_953),
.Y(n_1065)
);

OA22x2_ASAP7_75t_L g1066 ( 
.A1(n_969),
.A2(n_997),
.B1(n_976),
.B2(n_961),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_961),
.B(n_885),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_859),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_988),
.B(n_995),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_852),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_992),
.B(n_993),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_992),
.B(n_966),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_861),
.B(n_949),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_896),
.B(n_951),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_910),
.Y(n_1075)
);

AO32x2_ASAP7_75t_L g1076 ( 
.A1(n_916),
.A2(n_983),
.A3(n_967),
.B1(n_925),
.B2(n_852),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_910),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_901),
.B(n_895),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_910),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_904),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_855),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1083)
);

NOR4xp25_ASAP7_75t_L g1084 ( 
.A(n_966),
.B(n_954),
.C(n_958),
.D(n_985),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_904),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_904),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_910),
.B(n_808),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_869),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_888),
.B(n_733),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_904),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1092)
);

NOR4xp25_ASAP7_75t_L g1093 ( 
.A(n_966),
.B(n_954),
.C(n_958),
.D(n_985),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_919),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_978),
.A2(n_726),
.B(n_895),
.C(n_972),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_R g1098 ( 
.A(n_869),
.B(n_602),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_910),
.B(n_808),
.Y(n_1099)
);

BUFx4_ASAP7_75t_SL g1100 ( 
.A(n_856),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_928),
.B(n_576),
.C(n_892),
.Y(n_1101)
);

BUFx4_ASAP7_75t_SL g1102 ( 
.A(n_856),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_895),
.A2(n_901),
.B1(n_990),
.B2(n_853),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_919),
.B(n_910),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_855),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_938),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_895),
.B(n_939),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_904),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_869),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_895),
.A2(n_901),
.B1(n_990),
.B2(n_853),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_895),
.B(n_939),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_855),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_904),
.Y(n_1117)
);

NAND3x1_ASAP7_75t_L g1118 ( 
.A(n_984),
.B(n_769),
.C(n_817),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_862),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_959),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_910),
.B(n_808),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_869),
.B(n_787),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_869),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_895),
.A2(n_901),
.B1(n_990),
.B2(n_853),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_888),
.B(n_733),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_901),
.B(n_895),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_904),
.Y(n_1127)
);

AOI211x1_ASAP7_75t_L g1128 ( 
.A1(n_909),
.A2(n_916),
.B(n_981),
.C(n_931),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_978),
.A2(n_726),
.B(n_895),
.C(n_972),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_SL g1131 ( 
.A(n_984),
.B(n_665),
.C(n_552),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_855),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_895),
.A2(n_901),
.B1(n_990),
.B2(n_853),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_901),
.B(n_895),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_944),
.A2(n_875),
.B(n_864),
.Y(n_1135)
);

INVx6_ASAP7_75t_SL g1136 ( 
.A(n_929),
.Y(n_1136)
);

OAI21xp33_ASAP7_75t_SL g1137 ( 
.A1(n_888),
.A2(n_895),
.B(n_901),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_895),
.B(n_939),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_872),
.A2(n_729),
.B(n_719),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_904),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_862),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_895),
.B(n_939),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_888),
.B(n_733),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_917),
.A2(n_784),
.B1(n_552),
.B2(n_674),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_854),
.B(n_805),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_895),
.B(n_939),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_868),
.A2(n_729),
.A3(n_719),
.B(n_928),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_869),
.B(n_787),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_904),
.Y(n_1151)
);

BUFx2_ASAP7_75t_SL g1152 ( 
.A(n_1122),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1078),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1062),
.B(n_1078),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1128),
.B(n_1027),
.C(n_1137),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1094),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1104),
.B(n_1114),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_SL g1158 ( 
.A(n_1094),
.B(n_1147),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1113),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1104),
.Y(n_1160)
);

BUFx2_ASAP7_75t_SL g1161 ( 
.A(n_1150),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1080),
.A2(n_1088),
.B(n_1083),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1080),
.A2(n_1088),
.B(n_1083),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1053),
.B(n_1005),
.C(n_1055),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1034),
.A2(n_1031),
.B(n_1016),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1096),
.A2(n_1130),
.B(n_1011),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1011),
.A2(n_1026),
.B(n_1046),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1094),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1095),
.A2(n_1108),
.B(n_1105),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_1094),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1110),
.A2(n_1115),
.B1(n_1138),
.B2(n_1144),
.C(n_1148),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1040),
.A2(n_1042),
.B1(n_1066),
.B2(n_1054),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1114),
.A2(n_1124),
.B1(n_1133),
.B2(n_1066),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1017),
.A2(n_1140),
.B(n_1111),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1111),
.A2(n_1141),
.B(n_1140),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1126),
.A2(n_1134),
.B1(n_1118),
.B2(n_1125),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1141),
.A2(n_1058),
.B(n_1048),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1007),
.Y(n_1178)
);

AO32x2_ASAP7_75t_L g1179 ( 
.A1(n_1024),
.A2(n_1133),
.A3(n_1124),
.B1(n_1000),
.B2(n_1061),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1049),
.B(n_1023),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1062),
.B(n_1146),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1018),
.A2(n_999),
.B1(n_1040),
.B2(n_1057),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1007),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1136),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1025),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1081),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1100),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1049),
.B(n_1085),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1021),
.B(n_1090),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1086),
.B(n_1091),
.Y(n_1190)
);

OAI222xp33_ASAP7_75t_L g1191 ( 
.A1(n_1061),
.A2(n_1000),
.B1(n_1072),
.B2(n_1074),
.C1(n_1070),
.C2(n_1010),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1145),
.B(n_1033),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1132),
.B(n_1082),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1060),
.A2(n_1028),
.B(n_1059),
.C(n_1029),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1112),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1084),
.A2(n_1093),
.B1(n_1151),
.B2(n_1142),
.C(n_1117),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1132),
.B(n_1107),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1116),
.B(n_1032),
.Y(n_1200)
);

AO21x2_ASAP7_75t_L g1201 ( 
.A1(n_1051),
.A2(n_1003),
.B(n_1063),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1127),
.B(n_1041),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_SL g1204 ( 
.A(n_1147),
.B(n_1035),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1101),
.B(n_1009),
.C(n_1074),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1057),
.Y(n_1206)
);

OR2x2_ASAP7_75t_SL g1207 ( 
.A(n_1098),
.B(n_1131),
.Y(n_1207)
);

BUFx4f_ASAP7_75t_SL g1208 ( 
.A(n_1038),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1019),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1147),
.B(n_1012),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1089),
.A2(n_1001),
.B1(n_1123),
.B2(n_1012),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1064),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1050),
.A2(n_1013),
.B1(n_1006),
.B2(n_1044),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1039),
.A2(n_1065),
.B1(n_1056),
.B2(n_1059),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1022),
.A2(n_1028),
.B(n_1069),
.C(n_1045),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1047),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1036),
.Y(n_1218)
);

AO21x2_ASAP7_75t_L g1219 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1015),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1067),
.B(n_1045),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1014),
.B(n_1075),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1135),
.A2(n_1073),
.B(n_1068),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_998),
.B(n_1071),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1092),
.A2(n_1149),
.A3(n_1139),
.B(n_1129),
.Y(n_1224)
);

BUFx8_ASAP7_75t_L g1225 ( 
.A(n_1102),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1068),
.A2(n_1143),
.B(n_1004),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1020),
.A2(n_1121),
.B1(n_1099),
.B2(n_1087),
.C(n_1052),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1106),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1008),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1002),
.A2(n_1119),
.B(n_1076),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1008),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1092),
.A2(n_1097),
.B(n_1129),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1043),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1097),
.A2(n_1103),
.B(n_1129),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1097),
.B(n_1149),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1103),
.B(n_1120),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_1147),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1062),
.B(n_963),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_R g1239 ( 
.A(n_1113),
.B(n_869),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1104),
.A2(n_1124),
.B(n_1114),
.Y(n_1240)
);

NAND2x1_ASAP7_75t_L g1241 ( 
.A(n_1002),
.B(n_977),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1113),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1096),
.A2(n_1130),
.B(n_1011),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1080),
.A2(n_1088),
.B(n_1083),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1104),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1094),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1094),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_SL g1248 ( 
.A(n_1113),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1034),
.A2(n_1031),
.B(n_685),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1137),
.A2(n_784),
.B1(n_567),
.B2(n_552),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1170),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1170),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1170),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1225),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1153),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1170),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1166),
.A2(n_1243),
.B(n_1165),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1182),
.A2(n_1238),
.B1(n_1172),
.B2(n_1181),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1182),
.A2(n_1238),
.B1(n_1172),
.B2(n_1181),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1246),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1216),
.A2(n_1249),
.B(n_1164),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1249),
.A2(n_1195),
.B(n_1205),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1229),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1231),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1177),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1177),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1155),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1190),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1185),
.Y(n_1269)
);

AO221x2_ASAP7_75t_L g1270 ( 
.A1(n_1173),
.A2(n_1191),
.B1(n_1230),
.B2(n_1174),
.C(n_1157),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1186),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1193),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1196),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1202),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1165),
.A2(n_1175),
.B(n_1169),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1246),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1199),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1237),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1237),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1171),
.B(n_1154),
.Y(n_1280)
);

BUFx8_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1236),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1195),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1241),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1212),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1178),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1171),
.A2(n_1215),
.B1(n_1210),
.B2(n_1176),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1156),
.B(n_1247),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1217),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1154),
.B(n_1220),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1179),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1213),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1243),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1237),
.Y(n_1294)
);

AND2x2_ASAP7_75t_SL g1295 ( 
.A(n_1157),
.B(n_1210),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1226),
.B(n_1222),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1168),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1250),
.A2(n_1245),
.B1(n_1160),
.B2(n_1173),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1178),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1263),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1274),
.B(n_1198),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1282),
.B(n_1235),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1274),
.B(n_1198),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1282),
.B(n_1232),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1257),
.B(n_1232),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1258),
.A2(n_1240),
.B1(n_1192),
.B2(n_1160),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1257),
.B(n_1234),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1257),
.B(n_1162),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1264),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1280),
.A2(n_1192),
.B1(n_1245),
.B2(n_1214),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1293),
.B(n_1163),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1286),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1300),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1297),
.B(n_1224),
.Y(n_1316)
);

INVxp33_ASAP7_75t_L g1317 ( 
.A(n_1288),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1291),
.B(n_1201),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1291),
.B(n_1167),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1251),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1281),
.B(n_1225),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1251),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1275),
.B(n_1219),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1251),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1259),
.A2(n_1189),
.B1(n_1188),
.B2(n_1180),
.Y(n_1325)
);

BUFx2_ASAP7_75t_SL g1326 ( 
.A(n_1252),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1284),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1255),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1315),
.B(n_1308),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1325),
.A2(n_1295),
.B1(n_1287),
.B2(n_1292),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1301),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1316),
.B(n_1283),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1328),
.B(n_1265),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1328),
.B(n_1265),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1306),
.B(n_1295),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1306),
.B(n_1295),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1266),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1322),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1322),
.B(n_1252),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1313),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1305),
.B(n_1266),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1316),
.B(n_1302),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_SL g1343 ( 
.A(n_1326),
.B(n_1320),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1326),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1305),
.B(n_1270),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1322),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1310),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1303),
.B(n_1277),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1316),
.B(n_1268),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1319),
.B(n_1270),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1319),
.B(n_1270),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1313),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1302),
.B(n_1268),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1303),
.B(n_1272),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1303),
.B(n_1314),
.Y(n_1355)
);

NAND4xp25_ASAP7_75t_L g1356 ( 
.A(n_1325),
.B(n_1211),
.C(n_1290),
.D(n_1299),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1314),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1355),
.B(n_1312),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1342),
.B(n_1304),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1355),
.B(n_1312),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1342),
.B(n_1304),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1340),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1329),
.B(n_1315),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1345),
.B(n_1319),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1356),
.A2(n_1311),
.B1(n_1307),
.B2(n_1270),
.Y(n_1365)
);

NAND2x1_ASAP7_75t_L g1366 ( 
.A(n_1346),
.B(n_1327),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1337),
.B(n_1329),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1352),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1344),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1329),
.B(n_1315),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1344),
.B(n_1252),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_L g1373 ( 
.A(n_1346),
.B(n_1322),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1337),
.B(n_1309),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_L g1375 ( 
.A(n_1346),
.B(n_1253),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1329),
.B(n_1309),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1357),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1333),
.B(n_1334),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1343),
.Y(n_1379)
);

NAND2x1_ASAP7_75t_L g1380 ( 
.A(n_1346),
.B(n_1327),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_SL g1381 ( 
.A(n_1339),
.B(n_1281),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1331),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1374),
.B(n_1350),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1378),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1373),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1378),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1379),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1362),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1372),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1369),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1377),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1358),
.B(n_1333),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1374),
.B(n_1350),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1358),
.B(n_1334),
.Y(n_1394)
);

OAI31xp67_ASAP7_75t_L g1395 ( 
.A1(n_1365),
.A2(n_1356),
.A3(n_1321),
.B(n_1207),
.Y(n_1395)
);

NOR2x1_ASAP7_75t_L g1396 ( 
.A(n_1375),
.B(n_1233),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1359),
.B(n_1351),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1360),
.B(n_1332),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1367),
.B(n_1376),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1332),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1367),
.B(n_1335),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1366),
.B(n_1380),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1370),
.Y(n_1403)
);

INVxp33_ASAP7_75t_L g1404 ( 
.A(n_1381),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1392),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1396),
.A2(n_1330),
.B(n_1368),
.C(n_1191),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1392),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1403),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1399),
.B(n_1376),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1404),
.A2(n_1330),
.B(n_1372),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1384),
.B(n_1361),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1394),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1394),
.B(n_1364),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1398),
.Y(n_1414)
);

AOI211x1_ASAP7_75t_SL g1415 ( 
.A1(n_1395),
.A2(n_1353),
.B(n_1261),
.C(n_1262),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1402),
.A2(n_1351),
.B(n_1336),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1404),
.A2(n_1371),
.B1(n_1363),
.B2(n_1339),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1388),
.A2(n_1187),
.B(n_1267),
.C(n_1353),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1398),
.B(n_1354),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1397),
.A2(n_1307),
.B1(n_1382),
.B2(n_1267),
.C(n_1321),
.Y(n_1420)
);

AOI332xp33_ASAP7_75t_L g1421 ( 
.A1(n_1386),
.A2(n_1271),
.A3(n_1289),
.B1(n_1285),
.B2(n_1269),
.B3(n_1273),
.C1(n_1341),
.C2(n_1347),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1390),
.B(n_1354),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1400),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1402),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1391),
.B(n_1348),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1409),
.B(n_1399),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1405),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1415),
.A2(n_1387),
.B1(n_1385),
.B2(n_1281),
.C1(n_1389),
.C2(n_1239),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1407),
.B(n_1383),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1417),
.A2(n_1402),
.B1(n_1387),
.B2(n_1393),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1416),
.A2(n_1389),
.B(n_1254),
.C(n_1279),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1412),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1414),
.B(n_1400),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1408),
.Y(n_1434)
);

XNOR2x2_ASAP7_75t_L g1435 ( 
.A(n_1410),
.B(n_1281),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1419),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1419),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1411),
.B(n_1401),
.Y(n_1438)
);

AOI211xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1431),
.A2(n_1208),
.B(n_1420),
.C(n_1248),
.Y(n_1439)
);

NOR4xp25_ASAP7_75t_L g1440 ( 
.A(n_1434),
.B(n_1406),
.C(n_1418),
.D(n_1424),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1431),
.A2(n_1402),
.B(n_1424),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1436),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1428),
.B(n_1422),
.C(n_1425),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1437),
.B(n_1254),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1430),
.A2(n_1423),
.B(n_1422),
.C(n_1425),
.Y(n_1445)
);

AOI31xp33_ASAP7_75t_L g1446 ( 
.A1(n_1435),
.A2(n_1242),
.A3(n_1208),
.B(n_1339),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1427),
.A2(n_1409),
.B1(n_1401),
.B2(n_1371),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1438),
.B(n_1413),
.Y(n_1448)
);

OAI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1435),
.A2(n_1421),
.B(n_1209),
.C(n_1184),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1432),
.A2(n_1371),
.B1(n_1363),
.B2(n_1413),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1438),
.A2(n_1317),
.B(n_1256),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1433),
.B(n_1248),
.Y(n_1452)
);

AOI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1429),
.A2(n_1335),
.B1(n_1336),
.B2(n_1363),
.C(n_1349),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1440),
.B(n_1426),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1446),
.A2(n_1343),
.B(n_1158),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1341),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1449),
.B(n_1227),
.C(n_1218),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1449),
.A2(n_1279),
.B(n_1278),
.C(n_1294),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1451),
.A2(n_1338),
.B1(n_1320),
.B2(n_1324),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_SL g1460 ( 
.A(n_1439),
.B(n_1228),
.C(n_1183),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1441),
.B(n_1338),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1450),
.B(n_1318),
.Y(n_1462)
);

XOR2x2_ASAP7_75t_L g1463 ( 
.A(n_1444),
.B(n_1194),
.Y(n_1463)
);

NOR3x1_ASAP7_75t_L g1464 ( 
.A(n_1443),
.B(n_1294),
.C(n_1278),
.Y(n_1464)
);

NOR3xp33_ASAP7_75t_L g1465 ( 
.A(n_1460),
.B(n_1445),
.C(n_1452),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1454),
.Y(n_1466)
);

AOI211x1_ASAP7_75t_L g1467 ( 
.A1(n_1454),
.A2(n_1448),
.B(n_1442),
.C(n_1453),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1458),
.B(n_1227),
.C(n_1298),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1457),
.B(n_1298),
.C(n_1271),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1456),
.B(n_1323),
.Y(n_1470)
);

AND2x2_ASAP7_75t_SL g1471 ( 
.A(n_1464),
.B(n_1455),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1463),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1461),
.B(n_1152),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1462),
.Y(n_1474)
);

NAND4xp25_ASAP7_75t_L g1475 ( 
.A(n_1459),
.B(n_1161),
.C(n_1183),
.D(n_1228),
.Y(n_1475)
);

NAND4xp75_ASAP7_75t_L g1476 ( 
.A(n_1464),
.B(n_1324),
.C(n_1320),
.D(n_1276),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1466),
.B(n_1331),
.Y(n_1477)
);

NOR2x1_ASAP7_75t_L g1478 ( 
.A(n_1472),
.B(n_1469),
.Y(n_1478)
);

NAND2x1_ASAP7_75t_SL g1479 ( 
.A(n_1473),
.B(n_1253),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1467),
.B(n_1221),
.C(n_1200),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1468),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1465),
.B(n_1206),
.C(n_1256),
.D(n_1253),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1474),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1471),
.Y(n_1484)
);

NAND4xp75_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1203),
.C(n_1324),
.D(n_1204),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1481),
.B(n_1470),
.Y(n_1486)
);

NAND4xp75_ASAP7_75t_L g1487 ( 
.A(n_1478),
.B(n_1475),
.C(n_1197),
.D(n_1194),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1477),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1483),
.Y(n_1489)
);

NOR2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1484),
.B(n_1475),
.Y(n_1490)
);

NOR2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1487),
.B(n_1482),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1489),
.B(n_1480),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1492),
.A2(n_1486),
.B1(n_1488),
.B2(n_1490),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1493),
.Y(n_1494)
);

AOI22x1_ASAP7_75t_L g1495 ( 
.A1(n_1494),
.A2(n_1491),
.B1(n_1486),
.B2(n_1479),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1495),
.A2(n_1485),
.B1(n_1221),
.B2(n_1197),
.C(n_1206),
.Y(n_1496)
);

OAI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1496),
.A2(n_1256),
.B(n_1223),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1497),
.B(n_1260),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1498),
.A2(n_1260),
.B1(n_1338),
.B2(n_1223),
.Y(n_1499)
);


endmodule