module fake_jpeg_15846_n_300 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_247;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_25),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_20),
.C(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_49),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_26),
.B1(n_18),
.B2(n_22),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_60),
.B1(n_22),
.B2(n_16),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_76),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_80),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_38),
.B1(n_31),
.B2(n_18),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_54),
.B1(n_81),
.B2(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_38),
.B1(n_31),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_83),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_20),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_23),
.B1(n_16),
.B2(n_29),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_24),
.B1(n_23),
.B2(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_97),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_56),
.C(n_36),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_72),
.C(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_17),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_17),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_75),
.B1(n_105),
.B2(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_92),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_117),
.C(n_127),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_71),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_121),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_83),
.B(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_83),
.B1(n_77),
.B2(n_66),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_77),
.B1(n_73),
.B2(n_66),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_13),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_92),
.Y(n_147)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_147),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_89),
.B(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_149),
.B1(n_111),
.B2(n_29),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_88),
.B(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_144),
.B1(n_146),
.B2(n_152),
.Y(n_172)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_86),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_95),
.B1(n_94),
.B2(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_95),
.B1(n_94),
.B2(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_131),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_91),
.B(n_98),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_94),
.B1(n_91),
.B2(n_99),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_97),
.C(n_56),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_27),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_131),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_121),
.B1(n_116),
.B2(n_109),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_165),
.B1(n_176),
.B2(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_161),
.B(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_156),
.B(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_122),
.B1(n_130),
.B2(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_127),
.C(n_124),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_174),
.C(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_111),
.B1(n_64),
.B2(n_61),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_56),
.C(n_58),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_64),
.B1(n_61),
.B2(n_23),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_41),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_42),
.CI(n_45),
.CON(n_183),
.SN(n_183)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_144),
.B1(n_140),
.B2(n_158),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_189),
.B1(n_190),
.B2(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_140),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_162),
.B(n_159),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_137),
.B1(n_155),
.B2(n_151),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_137),
.B1(n_148),
.B2(n_153),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_200),
.B(n_27),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_136),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_153),
.B1(n_61),
.B2(n_15),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_207),
.B1(n_186),
.B2(n_161),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_63),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_24),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_63),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_183),
.C(n_181),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_163),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_225),
.B(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_178),
.B1(n_169),
.B2(n_173),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_167),
.B1(n_183),
.B2(n_168),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_220),
.B1(n_226),
.B2(n_10),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_170),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_58),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_173),
.C(n_164),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_188),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_193),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_164),
.B1(n_81),
.B2(n_3),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_208),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_189),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_227),
.C(n_58),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_19),
.B1(n_15),
.B2(n_63),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_42),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_205),
.B(n_192),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_241),
.B(n_11),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_242),
.C(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_210),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_193),
.B1(n_195),
.B2(n_19),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_243),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_10),
.B(n_13),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_42),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_249),
.C(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_218),
.C(n_215),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_254),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_216),
.C(n_227),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_225),
.C(n_50),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_260),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_261),
.Y(n_265)
);

AOI31xp33_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_11),
.A3(n_10),
.B(n_3),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_266),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_229),
.B(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_245),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_0),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_275),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_255),
.B(n_259),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_284),
.B(n_285),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_50),
.A3(n_46),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_50),
.B(n_46),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_1),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_8),
.B1(n_9),
.B2(n_287),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_264),
.B(n_274),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.C(n_291),
.Y(n_293)
);

OAI31xp33_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_273),
.A3(n_269),
.B(n_5),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_3),
.B(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_276),
.B(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_8),
.C(n_9),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_298),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_296),
.Y(n_300)
);


endmodule