module fake_netlist_6_1470_n_103 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_103);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_103;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp67_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_21),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2x1p5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_30),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_39),
.B(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_36),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_40),
.B(n_37),
.C(n_42),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_39),
.B(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_39),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_37),
.B(n_23),
.C(n_22),
.Y(n_59)
);

AO31x2_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_20),
.A3(n_22),
.B(n_51),
.Y(n_60)
);

OAI21x1_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_51),
.B(n_48),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_52),
.B(n_44),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_44),
.B(n_33),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_48),
.B1(n_44),
.B2(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_61),
.B1(n_62),
.B2(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_68),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_49),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_59),
.B1(n_73),
.B2(n_53),
.C(n_46),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_71),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_68),
.B1(n_74),
.B2(n_53),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_69),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_66),
.B1(n_81),
.B2(n_46),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_84),
.B1(n_86),
.B2(n_85),
.Y(n_92)
);

AOI211x1_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_90),
.B(n_6),
.C(n_7),
.Y(n_93)
);

OAI211xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_88),
.B(n_6),
.C(n_7),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_4),
.C(n_8),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI31xp33_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_94),
.A3(n_8),
.B(n_9),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OAI322xp33_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_98),
.A3(n_97),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_4),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_99),
.B1(n_13),
.B2(n_11),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_11),
.B1(n_46),
.B2(n_39),
.C(n_58),
.Y(n_103)
);


endmodule