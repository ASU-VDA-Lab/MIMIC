module fake_jpeg_11049_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_23),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_11),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_36),
.B1(n_40),
.B2(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_56),
.B1(n_51),
.B2(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_38),
.B1(n_40),
.B2(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_63),
.B1(n_6),
.B2(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_49),
.B1(n_47),
.B2(n_33),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_65),
.B(n_5),
.C(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_7),
.B1(n_8),
.B2(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_15),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_2),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_52),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_77),
.C(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_17),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_80),
.B(n_9),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_4),
.C(n_5),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_82),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_86),
.B(n_76),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_79),
.C(n_84),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_74),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_75),
.A3(n_78),
.B1(n_24),
.B2(n_25),
.C1(n_27),
.C2(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_18),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_81),
.C(n_92),
.Y(n_96)
);


endmodule