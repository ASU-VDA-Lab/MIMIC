module fake_netlist_1_7745_n_701 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_701);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_701;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_0), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_49), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_5), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_73), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_75), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_18), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_61), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_70), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_69), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_23), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_20), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_12), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_3), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_19), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_30), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_62), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_51), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_38), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_4), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_16), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_27), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_25), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_48), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_10), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_9), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_12), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_63), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_8), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_40), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_35), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_65), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_3), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_18), .B(n_76), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_39), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_121), .B(n_0), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_101), .Y(n_127) );
AND2x6_ASAP7_75t_L g128 ( .A(n_83), .B(n_34), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_121), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_79), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_114), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_120), .B(n_36), .Y(n_136) );
XOR2xp5_ASAP7_75t_L g137 ( .A(n_113), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_96), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_78), .B(n_2), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_120), .B(n_41), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_81), .B(n_2), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_103), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_88), .B(n_4), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_103), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_103), .B(n_42), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_84), .Y(n_157) );
NOR3xp33_ASAP7_75t_L g158 ( .A(n_110), .B(n_6), .C(n_7), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_113), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_86), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_77), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_85), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_124), .B(n_6), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_116), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_129), .B(n_91), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_166), .B(n_108), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_167), .B(n_123), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_166), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_126), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_136), .A2(n_97), .B1(n_112), .B2(n_91), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_126), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_126), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_164), .B(n_87), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_162), .B(n_93), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_164), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_127), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_166), .B(n_87), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_156), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_129), .B(n_108), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_164), .B(n_104), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_129), .B(n_167), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_125), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_132), .B(n_112), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_153), .B(n_86), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
NAND3x1_ASAP7_75t_L g207 ( .A(n_158), .B(n_117), .C(n_115), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
BUFx10_ASAP7_75t_L g209 ( .A(n_127), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_151), .B(n_94), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_151), .B(n_106), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_132), .B(n_97), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_156), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_130), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
INVx1_ASAP7_75t_SL g217 ( .A(n_153), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_137), .A2(n_139), .B1(n_152), .B2(n_141), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_156), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_161), .B(n_105), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_135), .B(n_100), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_128), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
BUFx4f_ASAP7_75t_L g226 ( .A(n_136), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_135), .B(n_99), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_138), .B(n_106), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_160), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_149), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g232 ( .A(n_175), .B(n_136), .C(n_165), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_221), .B(n_139), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_221), .B(n_141), .Y(n_236) );
BUFx12f_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
NAND2xp33_ASAP7_75t_SL g238 ( .A(n_189), .B(n_228), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_185), .B(n_160), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_198), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_201), .B(n_143), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_212), .B(n_143), .Y(n_242) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_185), .B(n_131), .C(n_148), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_217), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_226), .A2(n_152), .B1(n_138), .B2(n_140), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_171), .B(n_163), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_226), .A2(n_140), .B1(n_147), .B2(n_150), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_226), .A2(n_142), .B1(n_163), .B2(n_161), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_172), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_189), .B(n_137), .C(n_117), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_196), .B(n_154), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_171), .B(n_157), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_179), .B(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_179), .B(n_150), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_190), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_215), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_169), .B(n_193), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_184), .A2(n_157), .B(n_155), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_211), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_222), .B(n_128), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_200), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_224), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_211), .B(n_159), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_195), .B(n_186), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_190), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_180), .B(n_146), .Y(n_272) );
OR2x6_ASAP7_75t_L g273 ( .A(n_211), .B(n_115), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_190), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_180), .B(n_146), .Y(n_275) );
INVx5_ASAP7_75t_L g276 ( .A(n_192), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_183), .B(n_146), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_202), .A2(n_146), .B1(n_128), .B2(n_156), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_209), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_218), .B(n_7), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_183), .A2(n_155), .B(n_149), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_186), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_187), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_227), .B(n_146), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_202), .A2(n_146), .B1(n_128), .B2(n_156), .Y(n_288) );
INVx5_ASAP7_75t_L g289 ( .A(n_192), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_210), .B(n_146), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_187), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_172), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_216), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_199), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_174), .B(n_128), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_199), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_171), .B(n_155), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_245), .A2(n_205), .B1(n_208), .B2(n_218), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_241), .A2(n_205), .B1(n_208), .B2(n_218), .Y(n_300) );
BUFx12f_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
BUFx2_ASAP7_75t_SL g302 ( .A(n_282), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_244), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_272), .A2(n_194), .B(n_181), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_256), .A2(n_223), .B(n_216), .C(n_220), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_257), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_260), .A2(n_223), .B(n_220), .C(n_191), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_269), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_235), .B(n_202), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_235), .B(n_202), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_236), .B(n_248), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_273), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_241), .A2(n_218), .B1(n_207), .B2(n_181), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_276), .Y(n_318) );
AOI21x1_ASAP7_75t_L g319 ( .A1(n_272), .A2(n_170), .B(n_168), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_231), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_236), .B(n_202), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_270), .B(n_181), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_231), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_231), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_258), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_246), .B(n_229), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_286), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_242), .A2(n_207), .B(n_213), .C(n_230), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_263), .A2(n_194), .B1(n_219), .B2(n_214), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_242), .A2(n_230), .B(n_213), .C(n_206), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_275), .A2(n_194), .B(n_219), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_239), .B(n_8), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_232), .B(n_219), .Y(n_334) );
O2A1O1Ixp5_ASAP7_75t_L g335 ( .A1(n_268), .A2(n_188), .B(n_173), .C(n_206), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_233), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_273), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_273), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_283), .A2(n_219), .B1(n_214), .B2(n_192), .Y(n_339) );
CKINVDCx8_ASAP7_75t_R g340 ( .A(n_246), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_233), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_233), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_267), .B(n_9), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_252), .B(n_219), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_285), .B(n_214), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_252), .Y(n_347) );
BUFx4f_ASAP7_75t_SL g348 ( .A(n_254), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_337), .A2(n_243), .B1(n_254), .B2(n_285), .Y(n_351) );
BUFx8_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
INVx6_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_300), .A2(n_238), .B1(n_251), .B2(n_253), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_319), .A2(n_262), .B(n_284), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_335), .A2(n_279), .B(n_275), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_347), .B(n_261), .Y(n_357) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_334), .A2(n_264), .B(n_287), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_303), .B(n_294), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_306), .B(n_297), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_300), .A2(n_297), .B(n_280), .C(n_247), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_347), .B(n_296), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_306), .B(n_234), .Y(n_363) );
AO31x2_ASAP7_75t_L g364 ( .A1(n_298), .A2(n_279), .A3(n_295), .B(n_290), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_316), .A2(n_250), .B1(n_277), .B2(n_281), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_299), .B(n_277), .Y(n_368) );
OR2x6_ASAP7_75t_L g369 ( .A(n_302), .B(n_295), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_307), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_333), .A2(n_288), .B1(n_265), .B2(n_240), .C(n_278), .Y(n_371) );
OAI21x1_ASAP7_75t_SL g372 ( .A1(n_317), .A2(n_255), .B(n_293), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_328), .B(n_292), .C(n_249), .Y(n_373) );
INVx8_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_325), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_314), .B(n_289), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_348), .Y(n_377) );
BUFx12f_ASAP7_75t_L g378 ( .A(n_309), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_316), .A2(n_149), .B1(n_155), .B2(n_192), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_320), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_376), .A2(n_330), .B(n_334), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_298), .B1(n_338), .B2(n_344), .C(n_326), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_315), .B1(n_326), .B2(n_321), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_366), .A2(n_321), .B1(n_313), .B2(n_310), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_370), .B(n_341), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_350), .A2(n_311), .B1(n_340), .B2(n_318), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_375), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_374), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_322), .B1(n_345), .B2(n_311), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_352), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_359), .A2(n_308), .B(n_305), .C(n_322), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_352), .A2(n_345), .B1(n_346), .B2(n_343), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_359), .B(n_339), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_331), .B1(n_304), .B2(n_155), .C(n_149), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g398 ( .A1(n_380), .A2(n_168), .B(n_173), .C(n_176), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_346), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_362), .A2(n_329), .B1(n_342), .B2(n_336), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_352), .A2(n_320), .B1(n_342), .B2(n_336), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_377), .B(n_11), .C(n_13), .D(n_15), .Y(n_404) );
AOI211xp5_ASAP7_75t_SL g405 ( .A1(n_371), .A2(n_11), .B(n_15), .C(n_16), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_368), .B(n_17), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
BUFx6f_ASAP7_75t_SL g408 ( .A(n_369), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_389), .B(n_364), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_383), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_401), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_403), .B(n_364), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_407), .B(n_363), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_392), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_403), .B(n_364), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_404), .B(n_373), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_407), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_390), .B(n_369), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_382), .B(n_364), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_386), .B(n_379), .Y(n_430) );
AOI33xp33_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_379), .A3(n_361), .B1(n_182), .B2(n_204), .B3(n_197), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_408), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_393), .B(n_378), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_405), .B(n_353), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_385), .B(n_353), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_391), .B(n_353), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_411), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_424), .B(n_381), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g447 ( .A1(n_441), .A2(n_394), .A3(n_393), .B(n_387), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_437), .B(n_369), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_421), .B(n_395), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_423), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_411), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_437), .B(n_369), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_423), .B(n_402), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_397), .A3(n_17), .B1(n_182), .B2(n_204), .B3(n_197), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_358), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_422), .B(n_176), .C(n_188), .D(n_178), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_417), .B(n_380), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_422), .A2(n_358), .B1(n_177), .B2(n_178), .C(n_378), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_426), .A2(n_374), .B1(n_358), .B2(n_323), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_424), .B(n_356), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_420), .B(n_356), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_410), .A2(n_374), .B(n_372), .Y(n_468) );
NAND2xp33_ASAP7_75t_L g469 ( .A(n_425), .B(n_374), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_412), .B(n_355), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_434), .B(n_177), .C(n_22), .D(n_24), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g472 ( .A1(n_441), .A2(n_430), .B1(n_429), .B2(n_416), .C1(n_413), .C2(n_434), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
AOI211x1_ASAP7_75t_L g474 ( .A1(n_416), .A2(n_21), .B(n_26), .C(n_28), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_410), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_423), .B(n_355), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_418), .B(n_343), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_409), .B(n_32), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_419), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_409), .B(n_33), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_415), .B(n_43), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_418), .B(n_343), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_440), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_428), .B(n_44), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_427), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_430), .B(n_45), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_434), .B(n_342), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_455), .B(n_429), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_487), .B(n_435), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_483), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_456), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_484), .B(n_432), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_449), .B(n_433), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_455), .B(n_439), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_473), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_465), .B(n_439), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_465), .B(n_438), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_467), .B(n_438), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_493), .B(n_433), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_483), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_473), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_459), .Y(n_513) );
OAI211xp5_ASAP7_75t_SL g514 ( .A1(n_447), .A2(n_431), .B(n_425), .C(n_436), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_467), .B(n_438), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_463), .B(n_444), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g517 ( .A(n_472), .B(n_442), .C(n_444), .D(n_433), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_463), .B(n_442), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_436), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_436), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_489), .B(n_432), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_492), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_492), .B(n_432), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_489), .B(n_426), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_459), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_476), .B(n_426), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g527 ( .A(n_471), .B(n_443), .C(n_47), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
AND2x4_ASAP7_75t_SL g529 ( .A(n_491), .B(n_443), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_443), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_490), .B(n_46), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_461), .B(n_50), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_461), .B(n_52), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_461), .B(n_54), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_55), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_490), .B(n_56), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_458), .B(n_58), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_484), .B(n_336), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_458), .B(n_64), .Y(n_541) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_464), .A2(n_324), .B(n_323), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_479), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_481), .B(n_66), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_466), .B(n_67), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_482), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_445), .B(n_72), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_486), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_481), .B(n_74), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_446), .B(n_324), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_503), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_510), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_548), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_499), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_535), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_497), .B(n_494), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_540), .B(n_500), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
NOR3xp33_ASAP7_75t_SL g565 ( .A(n_517), .B(n_462), .C(n_460), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_520), .B(n_466), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_545), .B(n_446), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_548), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_520), .B(n_450), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_518), .B(n_450), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_518), .B(n_475), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_516), .B(n_507), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_512), .B(n_452), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_516), .B(n_475), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_508), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_527), .B(n_474), .C(n_457), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_526), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_507), .B(n_478), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_514), .B(n_494), .C(n_495), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_502), .B(n_484), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_521), .Y(n_582) );
AND4x1_ASAP7_75t_L g583 ( .A(n_501), .B(n_468), .C(n_485), .D(n_469), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_550), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_515), .B(n_453), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_453), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_502), .B(n_505), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_505), .B(n_448), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_519), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_549), .A2(n_469), .B(n_488), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_519), .B(n_448), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_506), .B(n_485), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_509), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_498), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_496), .B(n_480), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_498), .B(n_324), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_506), .B(n_323), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_524), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_544), .B(n_289), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_289), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_523), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_530), .B(n_289), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_276), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_551), .B(n_276), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_553), .B(n_276), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_525), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_559), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_576), .B(n_500), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_582), .B(n_525), .Y(n_610) );
AOI222xp33_ASAP7_75t_L g611 ( .A1(n_577), .A2(n_541), .B1(n_533), .B2(n_532), .C1(n_534), .C2(n_547), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_578), .B(n_511), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_587), .B(n_547), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_594), .B(n_511), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_565), .A2(n_533), .B1(n_532), .B2(n_534), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_567), .B(n_513), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_562), .A2(n_541), .B1(n_537), .B2(n_540), .C1(n_529), .C2(n_552), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_572), .B(n_511), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_572), .B(n_513), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_580), .A2(n_590), .B1(n_581), .B2(n_595), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_563), .A2(n_549), .B(n_546), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_593), .B(n_513), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_594), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_563), .A2(n_542), .B(n_529), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_555), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_563), .A2(n_542), .B(n_554), .Y(n_630) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_568), .Y(n_631) );
AOI332xp33_ASAP7_75t_L g632 ( .A1(n_589), .A2(n_537), .A3(n_531), .B1(n_539), .B2(n_536), .B3(n_542), .C1(n_192), .C2(n_214), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_595), .A2(n_601), .B1(n_579), .B2(n_560), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_591), .B(n_259), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_579), .A2(n_203), .B(n_214), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_591), .A2(n_203), .B1(n_259), .B2(n_271), .Y(n_636) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_566), .A2(n_203), .B(n_259), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_566), .B(n_271), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_599), .B(n_203), .C(n_271), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_569), .B(n_274), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_556), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_585), .B(n_203), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_633), .B(n_586), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_620), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_616), .B(n_583), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_623), .A2(n_561), .A3(n_564), .B(n_573), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_628), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g648 ( .A1(n_623), .A2(n_574), .B(n_570), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_626), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_614), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_611), .A2(n_574), .B1(n_570), .B2(n_571), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_629), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_607), .B(n_586), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_609), .B(n_585), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_609), .A2(n_557), .B1(n_575), .B2(n_588), .C(n_568), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_624), .B(n_605), .C(n_604), .Y(n_656) );
AOI221x1_ASAP7_75t_L g657 ( .A1(n_627), .A2(n_557), .B1(n_575), .B2(n_584), .C(n_602), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_627), .B(n_584), .Y(n_658) );
AOI21xp33_ASAP7_75t_SL g659 ( .A1(n_618), .A2(n_606), .B(n_596), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_641), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_614), .B(n_606), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_621), .B(n_569), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_608), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_610), .B(n_571), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g665 ( .A1(n_612), .A2(n_600), .A3(n_602), .B(n_592), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_655), .B(n_617), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_651), .A2(n_619), .B1(n_613), .B2(n_631), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_648), .A2(n_625), .B(n_631), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g669 ( .A1(n_645), .A2(n_592), .A3(n_637), .B1(n_622), .B2(n_615), .C1(n_642), .C2(n_635), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_644), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_645), .A2(n_630), .B(n_639), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_661), .Y(n_672) );
AOI221xp5_ASAP7_75t_SL g673 ( .A1(n_659), .A2(n_630), .B1(n_636), .B2(n_600), .C(n_638), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_647), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_652), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_660), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_663), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_646), .A2(n_636), .B1(n_597), .B2(n_639), .C(n_632), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_653), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_671), .A2(n_657), .B(n_665), .C(n_649), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_672), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_666), .B(n_643), .Y(n_682) );
INVxp33_ASAP7_75t_L g683 ( .A(n_673), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_668), .A2(n_658), .B(n_661), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g685 ( .A(n_669), .B(n_658), .C(n_656), .Y(n_685) );
OAI22xp33_ASAP7_75t_SL g686 ( .A1(n_672), .A2(n_650), .B1(n_654), .B2(n_664), .Y(n_686) );
OAI222xp33_ASAP7_75t_L g687 ( .A1(n_667), .A2(n_650), .B1(n_662), .B2(n_634), .C1(n_596), .C2(n_640), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_681), .Y(n_688) );
NOR3xp33_ASAP7_75t_SL g689 ( .A(n_685), .B(n_678), .C(n_679), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_682), .B(n_677), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_683), .B(n_680), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_688), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_691), .B(n_686), .C(n_684), .Y(n_693) );
AND5x1_ASAP7_75t_L g694 ( .A(n_689), .B(n_678), .C(n_687), .D(n_670), .E(n_674), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_692), .B(n_690), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_693), .B(n_675), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_695), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_697), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_696), .B(n_694), .Y(n_699) );
OR2x6_ASAP7_75t_L g700 ( .A(n_699), .B(n_676), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_274), .B1(n_603), .B2(n_692), .C(n_693), .Y(n_701) );
endmodule