module fake_jpeg_10967_n_477 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_477);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_477;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_17),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_55),
.B(n_61),
.Y(n_149)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_67),
.Y(n_99)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_82),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_79),
.Y(n_111)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_33),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_16),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_89),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_0),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_96),
.Y(n_151)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_35),
.B(n_0),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_42),
.B1(n_32),
.B2(n_23),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_103),
.A2(n_109),
.B1(n_117),
.B2(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_23),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_46),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_52),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_42),
.B1(n_44),
.B2(n_43),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_123),
.A2(n_122),
.B1(n_112),
.B2(n_133),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_51),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_130),
.B1(n_134),
.B2(n_141),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_89),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_62),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_86),
.A2(n_21),
.B1(n_31),
.B2(n_28),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_50),
.A2(n_38),
.B1(n_31),
.B2(n_28),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_22),
.B1(n_57),
.B2(n_72),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_76),
.A2(n_31),
.B1(n_28),
.B2(n_22),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_94),
.B1(n_19),
.B2(n_5),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_68),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_70),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_198),
.C(n_200),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_103),
.A2(n_69),
.B1(n_93),
.B2(n_90),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_127),
.B(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_175),
.Y(n_211)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_182),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_146),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_123),
.A2(n_22),
.B1(n_57),
.B2(n_85),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_89),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_1),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_21),
.B1(n_84),
.B2(n_77),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_178),
.A2(n_203),
.B(n_15),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_184),
.B1(n_189),
.B2(n_190),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_111),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_183),
.B1(n_188),
.B2(n_192),
.Y(n_236)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_99),
.B(n_100),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_111),
.A2(n_19),
.B1(n_4),
.B2(n_6),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_19),
.B1(n_4),
.B2(n_6),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_101),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_195),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_197),
.Y(n_219)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_106),
.B1(n_120),
.B2(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_112),
.A2(n_19),
.B1(n_7),
.B2(n_10),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_133),
.A2(n_1),
.B1(n_7),
.B2(n_10),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_193),
.A2(n_114),
.B1(n_137),
.B2(n_98),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_119),
.A2(n_1),
.B1(n_10),
.B2(n_11),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_201),
.B1(n_204),
.B2(n_132),
.Y(n_248)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_202),
.Y(n_251)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_125),
.B(n_10),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_11),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_129),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_122),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_205),
.B(n_206),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_129),
.C(n_15),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_228),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_136),
.B(n_102),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_162),
.A2(n_135),
.B1(n_118),
.B2(n_113),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_226),
.B1(n_247),
.B2(n_178),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_128),
.B1(n_102),
.B2(n_136),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_152),
.B(n_175),
.CI(n_154),
.CON(n_228),
.SN(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_152),
.A2(n_142),
.B1(n_113),
.B2(n_137),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_237),
.B1(n_246),
.B2(n_153),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_176),
.A2(n_127),
.B(n_104),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_245),
.Y(n_269)
);

OR2x2_ASAP7_75t_SL g234 ( 
.A(n_198),
.B(n_104),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g291 ( 
.A(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_137),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_238),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_114),
.B1(n_98),
.B2(n_121),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_177),
.A2(n_104),
.B(n_132),
.C(n_121),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_155),
.B(n_132),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_250),
.C(n_198),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_248),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_158),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_156),
.A2(n_165),
.B1(n_166),
.B2(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_121),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_160),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_250),
.C(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_171),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_258),
.B(n_268),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_272),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_165),
.B1(n_190),
.B2(n_179),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_160),
.B1(n_189),
.B2(n_153),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_271),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_229),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_211),
.B(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_208),
.B(n_157),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_270),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_184),
.B1(n_166),
.B2(n_163),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_277),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_219),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_206),
.A2(n_191),
.B(n_161),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_238),
.B(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_174),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_283),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_197),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_208),
.B(n_219),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_288),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_213),
.A2(n_166),
.B1(n_196),
.B2(n_181),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_289),
.B1(n_232),
.B2(n_237),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_199),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_213),
.A2(n_195),
.B1(n_159),
.B2(n_164),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_230),
.A2(n_202),
.B1(n_170),
.B2(n_169),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_207),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_230),
.A2(n_169),
.B1(n_170),
.B2(n_187),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_290),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_294),
.A2(n_305),
.B(n_306),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_296),
.A2(n_300),
.B1(n_313),
.B2(n_261),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_205),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_298),
.C(n_301),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_231),
.B(n_216),
.C(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_221),
.C(n_217),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_244),
.B(n_226),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_281),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_234),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_309),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_236),
.B1(n_221),
.B2(n_229),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_330),
.C(n_286),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_275),
.A2(n_245),
.B(n_224),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

AOI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_267),
.A2(n_210),
.B(n_240),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_273),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_331),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_224),
.C(n_214),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_292),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_287),
.B1(n_260),
.B2(n_283),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_332),
.A2(n_333),
.B1(n_346),
.B2(n_352),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_259),
.B1(n_286),
.B2(n_272),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_252),
.Y(n_336)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_266),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_349),
.C(n_350),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_329),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_361),
.Y(n_364)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_345),
.A2(n_355),
.B1(n_360),
.B2(n_299),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_303),
.A2(n_291),
.B1(n_255),
.B2(n_271),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_274),
.Y(n_347)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_280),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_348),
.B(n_357),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_291),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_304),
.A2(n_286),
.B1(n_279),
.B2(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_313),
.A2(n_253),
.B1(n_240),
.B2(n_243),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_214),
.C(n_239),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_350),
.C(n_344),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_312),
.B(n_243),
.CI(n_227),
.CON(n_357),
.SN(n_357)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_359),
.A2(n_330),
.B1(n_303),
.B2(n_310),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_296),
.A2(n_306),
.B1(n_305),
.B2(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_331),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_348),
.B(n_310),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_374),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_301),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_373),
.A2(n_375),
.B1(n_376),
.B2(n_388),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_336),
.B(n_323),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_360),
.A2(n_307),
.B1(n_318),
.B2(n_294),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_306),
.B(n_312),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_378),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_339),
.B(n_314),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_380),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_384),
.C(n_356),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_323),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_382),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_320),
.C(n_315),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_327),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_324),
.B(n_322),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_387),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_354),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_355),
.B1(n_335),
.B2(n_341),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_332),
.B(n_315),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_351),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_381),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_379),
.Y(n_394)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_394),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_364),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_396),
.B(n_401),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_406),
.C(n_408),
.Y(n_415)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_334),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_388),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_351),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_411),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_365),
.A2(n_338),
.B1(n_335),
.B2(n_333),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_405),
.A2(n_368),
.B1(n_367),
.B2(n_383),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_346),
.C(n_340),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_352),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_409),
.B(n_410),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_357),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_378),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_398),
.Y(n_412)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_SL g414 ( 
.A1(n_390),
.A2(n_386),
.B(n_376),
.C(n_363),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_395),
.A2(n_368),
.B1(n_363),
.B2(n_377),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_400),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_383),
.B1(n_367),
.B2(n_370),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_426),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_420),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_407),
.B(n_374),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_425),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_408),
.A2(n_395),
.B(n_411),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_424),
.A2(n_428),
.B(n_322),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_391),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_404),
.A2(n_389),
.B1(n_377),
.B2(n_369),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_334),
.Y(n_429)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_432),
.Y(n_447)
);

AOI322xp5_ASAP7_75t_SL g432 ( 
.A1(n_419),
.A2(n_410),
.A3(n_409),
.B1(n_403),
.B2(n_392),
.C1(n_299),
.C2(n_406),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_393),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_423),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_420),
.B1(n_369),
.B2(n_394),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_436),
.A2(n_422),
.B1(n_418),
.B2(n_414),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_399),
.C(n_393),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_443),
.C(n_426),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_424),
.B(n_428),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_361),
.C(n_353),
.Y(n_443)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_441),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_445),
.Y(n_459)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_435),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_443),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_446),
.A2(n_442),
.B(n_437),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_449),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_450),
.B(n_454),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_453),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_439),
.A2(n_427),
.B(n_413),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_452),
.A2(n_433),
.B(n_439),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_414),
.C(n_343),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_430),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_SL g456 ( 
.A1(n_455),
.A2(n_437),
.B(n_414),
.C(n_434),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_458),
.C(n_321),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_457),
.A2(n_454),
.B1(n_463),
.B2(n_450),
.Y(n_465)
);

OAI221xp5_ASAP7_75t_L g460 ( 
.A1(n_447),
.A2(n_430),
.B1(n_431),
.B2(n_342),
.C(n_327),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_460),
.A2(n_464),
.B1(n_362),
.B2(n_309),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_466),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_449),
.B(n_444),
.C(n_311),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_469),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_SL g468 ( 
.A(n_461),
.B(n_448),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_468),
.A2(n_459),
.B(n_460),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_321),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_462),
.B(n_466),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_473),
.B(n_474),
.C(n_471),
.Y(n_475)
);

OAI321xp33_ASAP7_75t_L g476 ( 
.A1(n_475),
.A2(n_302),
.A3(n_316),
.B1(n_472),
.B2(n_474),
.C(n_459),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_476),
.B(n_302),
.Y(n_477)
);


endmodule