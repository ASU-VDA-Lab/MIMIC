module fake_jpeg_6478_n_208 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_32),
.B1(n_26),
.B2(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.Y(n_38)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_43),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_14),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_52),
.B1(n_19),
.B2(n_16),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_14),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_63),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_31),
.B(n_29),
.C(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_23),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_54),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_45),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_52),
.B1(n_40),
.B2(n_50),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_82),
.Y(n_104)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_53),
.B1(n_48),
.B2(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_32),
.B1(n_47),
.B2(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_33),
.B1(n_24),
.B2(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_66),
.B(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_101),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_46),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_85),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_71),
.B(n_73),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_88),
.B(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_105),
.B1(n_98),
.B2(n_111),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_100),
.B1(n_75),
.B2(n_95),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_125),
.B(n_100),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_78),
.B(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_75),
.B1(n_79),
.B2(n_69),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_146),
.B1(n_115),
.B2(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_104),
.C(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_142),
.C(n_145),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_93),
.C(n_103),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_97),
.C(n_76),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_102),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_122),
.C(n_126),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_149),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_95),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_14),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_162),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_147),
.B(n_145),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_125),
.B1(n_116),
.B2(n_124),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_163),
.B1(n_142),
.B2(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_154),
.Y(n_171)
);

AOI21x1_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_125),
.B(n_117),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_14),
.B(n_22),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_116),
.C(n_13),
.D(n_12),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_12),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_57),
.B1(n_70),
.B2(n_99),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_138),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_14),
.B(n_22),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_158),
.B1(n_153),
.B2(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_172),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_170),
.B(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_51),
.C(n_45),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_22),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_21),
.B1(n_51),
.B2(n_25),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_51),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_25),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_177),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_184),
.Y(n_189)
);

BUFx12f_ASAP7_75t_SL g182 ( 
.A(n_166),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_153),
.B1(n_25),
.B2(n_22),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_168),
.A3(n_166),
.B1(n_169),
.B2(n_11),
.C1(n_5),
.C2(n_6),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_175),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_8),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_182),
.C(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_189),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_188),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_9),
.B1(n_2),
.B2(n_8),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_9),
.B(n_201),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_194),
.C(n_195),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);


endmodule