module fake_aes_9692_n_678 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_678);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_678;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_38), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_63), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_80), .Y(n_89) );
BUFx5_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_74), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_56), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_83), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_50), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_75), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_84), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_32), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_85), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_6), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_5), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_20), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_78), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_31), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_68), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_81), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_34), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_12), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_45), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_54), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_55), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_69), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_82), .Y(n_120) );
CKINVDCx14_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_44), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g123 ( .A(n_17), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_41), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_17), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
CKINVDCx8_ASAP7_75t_R g128 ( .A(n_95), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_114), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_114), .Y(n_131) );
OR2x6_ASAP7_75t_L g132 ( .A(n_102), .B(n_0), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
OAI22x1_ASAP7_75t_R g134 ( .A1(n_110), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_123), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_94), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_123), .B(n_2), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_93), .B(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_100), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_109), .B(n_3), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_104), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_109), .B(n_4), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_105), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_121), .B(n_7), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_111), .B(n_37), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_106), .B(n_8), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_112), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_135), .B(n_92), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_141), .A2(n_108), .B1(n_121), .B2(n_126), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_143), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_130), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_128), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_153), .Y(n_165) );
BUFx10_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_128), .Y(n_170) );
AO22x2_ASAP7_75t_L g171 ( .A1(n_147), .A2(n_155), .B1(n_141), .B2(n_138), .Y(n_171) );
INVx1_ASAP7_75t_SL g172 ( .A(n_154), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_132), .B(n_125), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_138), .B(n_90), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_141), .B(n_118), .C(n_119), .Y(n_180) );
BUFx10_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx6_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_145), .B(n_101), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_149), .B(n_87), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
BUFx2_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_148), .B(n_89), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_151), .B(n_90), .Y(n_193) );
CKINVDCx6p67_ASAP7_75t_R g194 ( .A(n_132), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_175), .A2(n_132), .B1(n_155), .B2(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_178), .B(n_151), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_168), .B(n_133), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_178), .B(n_149), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_163), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_193), .B(n_133), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_194), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_158), .A2(n_156), .B(n_137), .C(n_144), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_181), .B(n_155), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_181), .B(n_155), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_193), .B(n_137), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g209 ( .A1(n_170), .A2(n_124), .B1(n_110), .B2(n_117), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_158), .B(n_140), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_188), .B(n_140), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_182), .Y(n_212) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_165), .B(n_117), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_180), .A2(n_156), .B(n_144), .C(n_142), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_181), .B(n_142), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_181), .B(n_113), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_182), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_188), .B(n_127), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_186), .B(n_127), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_165), .B(n_98), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_159), .B(n_146), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_175), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_172), .B(n_146), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
NAND2x1_ASAP7_75t_L g226 ( .A(n_175), .B(n_132), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_184), .B(n_116), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_124), .B1(n_122), .B2(n_150), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_165), .B(n_120), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_165), .B(n_122), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_171), .A2(n_150), .B1(n_143), .B2(n_97), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_161), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_191), .B(n_91), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_175), .A2(n_150), .B1(n_143), .B2(n_131), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_175), .B(n_150), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_150), .B(n_143), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_171), .A2(n_150), .B1(n_131), .B2(n_129), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_171), .B(n_131), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_171), .B(n_131), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_194), .B(n_131), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_164), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_167), .B(n_129), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_167), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_179), .B(n_129), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g245 ( .A(n_204), .B(n_157), .C(n_134), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_223), .B(n_176), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_224), .B(n_174), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_196), .B(n_174), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_195), .A2(n_176), .B1(n_174), .B2(n_169), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_200), .B(n_174), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_206), .A2(n_176), .B(n_169), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_228), .B(n_192), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_169), .B(n_177), .C(n_189), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_207), .A2(n_176), .B(n_177), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_222), .A2(n_177), .B(n_168), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_203), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_198), .B(n_192), .Y(n_258) );
NOR2xp67_ASAP7_75t_L g259 ( .A(n_199), .B(n_8), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_205), .A2(n_179), .B(n_189), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_210), .B(n_185), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_232), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_215), .A2(n_168), .B(n_187), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_209), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_219), .A2(n_168), .B(n_187), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_233), .B(n_168), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_205), .A2(n_168), .B(n_185), .Y(n_267) );
AO22x1_ASAP7_75t_L g268 ( .A1(n_203), .A2(n_134), .B1(n_10), .B2(n_11), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_223), .B(n_129), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_220), .A2(n_166), .B(n_173), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_228), .A2(n_129), .B1(n_183), .B2(n_173), .Y(n_271) );
AOI22x1_ASAP7_75t_L g272 ( .A1(n_225), .A2(n_190), .B1(n_173), .B2(n_160), .Y(n_272) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_226), .A2(n_166), .B(n_183), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_225), .A2(n_173), .B(n_160), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_231), .A2(n_183), .B1(n_160), .B2(n_166), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_209), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_211), .B(n_166), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_213), .B(n_9), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_218), .B(n_160), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_241), .B(n_9), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_229), .A2(n_190), .B(n_183), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_227), .B(n_10), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_237), .B(n_190), .Y(n_284) );
OR2x6_ASAP7_75t_SL g285 ( .A(n_199), .B(n_11), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_231), .A2(n_190), .B(n_183), .C(n_14), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_243), .B(n_12), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_213), .A2(n_190), .B1(n_15), .B2(n_16), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_243), .B(n_13), .Y(n_290) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_242), .A2(n_190), .B(n_46), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_201), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_235), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_255), .A2(n_240), .B(n_216), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_248), .A2(n_201), .B(n_202), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_250), .A2(n_202), .B(n_212), .Y(n_297) );
AO31x2_ASAP7_75t_L g298 ( .A1(n_253), .A2(n_239), .A3(n_238), .B(n_214), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_289), .B(n_237), .C(n_230), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_291), .A2(n_273), .B(n_272), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_283), .A2(n_235), .B(n_236), .C(n_230), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_264), .B(n_277), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_290), .Y(n_304) );
BUFx2_ASAP7_75t_R g305 ( .A(n_285), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_275), .A2(n_236), .B(n_244), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
O2A1O1Ixp5_ASAP7_75t_L g308 ( .A1(n_284), .A2(n_221), .B(n_217), .C(n_212), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_221), .B(n_217), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_267), .A2(n_234), .B(n_197), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_265), .A2(n_43), .B(n_79), .Y(n_311) );
AO31x2_ASAP7_75t_L g312 ( .A1(n_253), .A2(n_13), .A3(n_15), .B(n_16), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_257), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_252), .B(n_18), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_268), .A2(n_245), .B(n_259), .C(n_271), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_247), .A2(n_49), .B(n_19), .Y(n_316) );
NOR2xp33_ASAP7_75t_SL g317 ( .A(n_249), .B(n_51), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_247), .A2(n_52), .B(n_21), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_293), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_278), .A2(n_53), .B(n_22), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_287), .B(n_18), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_251), .A2(n_23), .B(n_24), .Y(n_322) );
AO31x2_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_25), .A3(n_26), .B(n_27), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_254), .A2(n_28), .B(n_29), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_245), .B(n_30), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_266), .A2(n_35), .B(n_36), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_261), .B(n_40), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_293), .B(n_42), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_283), .B(n_57), .C(n_58), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_313), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_321), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_321), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g334 ( .A1(n_325), .A2(n_279), .B1(n_284), .B2(n_258), .C1(n_293), .C2(n_260), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
AOI21xp5_ASAP7_75t_SL g337 ( .A1(n_302), .A2(n_274), .B(n_269), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_303), .B(n_262), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
AOI21x1_ASAP7_75t_L g341 ( .A1(n_301), .A2(n_294), .B(n_329), .Y(n_341) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_299), .A2(n_256), .B(n_246), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_330), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_295), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_300), .B(n_292), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_304), .B(n_274), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_311), .A2(n_270), .B(n_263), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_327), .A2(n_269), .B(n_246), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_314), .B(n_274), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_307), .Y(n_351) );
OA21x2_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_280), .B(n_266), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_297), .A2(n_269), .B(n_276), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_298), .B(n_59), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_60), .B(n_61), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_296), .A2(n_62), .B(n_64), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_350), .A2(n_299), .B(n_329), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_359), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_350), .A2(n_318), .B(n_316), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_340), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_359), .A2(n_326), .B(n_324), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_355), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_336), .B(n_298), .Y(n_367) );
OA21x2_ASAP7_75t_L g368 ( .A1(n_354), .A2(n_320), .B(n_310), .Y(n_368) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_337), .B(n_328), .Y(n_369) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_354), .A2(n_312), .B(n_323), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_353), .A2(n_323), .B(n_298), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_341), .B(n_348), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_333), .B(n_315), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_346), .B(n_323), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_346), .B(n_315), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_346), .B(n_317), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_345), .B(n_317), .Y(n_384) );
AOI21x1_ASAP7_75t_L g385 ( .A1(n_341), .A2(n_65), .B(n_66), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_347), .A2(n_67), .B(n_73), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_76), .B(n_86), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_380), .B(n_338), .Y(n_389) );
NAND2x1p5_ASAP7_75t_SL g390 ( .A(n_369), .B(n_345), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_381), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_381), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_382), .B(n_344), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_381), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_380), .B(n_338), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_384), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_382), .B(n_344), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_386), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
NOR2x1_ASAP7_75t_SL g403 ( .A(n_388), .B(n_349), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_382), .B(n_345), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_378), .B(n_331), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_386), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_382), .B(n_334), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_378), .A2(n_335), .B1(n_343), .B2(n_349), .C(n_358), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
INVx4_ASAP7_75t_SL g412 ( .A(n_367), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_372), .B(n_334), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_372), .B(n_351), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_375), .Y(n_415) );
OR2x6_ASAP7_75t_L g416 ( .A(n_384), .B(n_336), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_379), .B(n_342), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_379), .B(n_342), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_363), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_375), .B(n_351), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_375), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_379), .B(n_342), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_376), .B(n_342), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_384), .A2(n_357), .B1(n_352), .B2(n_339), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_376), .B(n_336), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_389), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_417), .B(n_422), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_408), .B(n_367), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_417), .B(n_367), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_418), .B(n_367), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_418), .B(n_367), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_422), .B(n_367), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_399), .B(n_383), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_408), .B(n_371), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_395), .B(n_383), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_391), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_395), .B(n_383), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_389), .B(n_398), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_371), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_398), .B(n_388), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_414), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_414), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_371), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_423), .B(n_371), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_401), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_413), .B(n_386), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_411), .B(n_371), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_421), .B(n_371), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_425), .B(n_377), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_423), .B(n_373), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_419), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_424), .B(n_385), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_425), .B(n_370), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_396), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_396), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_405), .B(n_357), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_416), .B(n_404), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_404), .B(n_373), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_412), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_416), .B(n_373), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_416), .B(n_373), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_397), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_428), .B(n_420), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_428), .B(n_426), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_477), .B(n_412), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_430), .B(n_412), .Y(n_486) );
AND2x2_ASAP7_75t_SL g487 ( .A(n_477), .B(n_424), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_450), .B(n_409), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_429), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_444), .B(n_357), .Y(n_490) );
NOR2xp67_ASAP7_75t_L g491 ( .A(n_477), .B(n_397), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_444), .B(n_416), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_477), .B(n_412), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_429), .B(n_419), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_475), .B(n_416), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_451), .B(n_410), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_430), .B(n_419), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_427), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_475), .B(n_390), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_439), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_438), .B(n_443), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_440), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_438), .B(n_407), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_457), .B(n_410), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_443), .B(n_407), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_442), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_431), .B(n_390), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_455), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_431), .B(n_390), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_474), .B(n_388), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_455), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_441), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_445), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_441), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_432), .B(n_403), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_445), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_448), .B(n_369), .C(n_358), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_447), .B(n_452), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
AND2x2_ASAP7_75t_SL g526 ( .A(n_478), .B(n_402), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_467), .B(n_403), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_449), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_456), .B(n_366), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_456), .B(n_432), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_447), .B(n_370), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_452), .B(n_370), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_454), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_433), .B(n_402), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_449), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_459), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_464), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_433), .B(n_402), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_434), .B(n_363), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_476), .B(n_459), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_507), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_484), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_485), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_524), .B(n_476), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_486), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_541), .B(n_437), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_488), .B(n_437), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_502), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_503), .B(n_465), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_434), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_538), .B(n_465), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_504), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_500), .A2(n_448), .B(n_468), .C(n_478), .Y(n_556) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_515), .B(n_479), .C(n_468), .D(n_369), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_508), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_490), .A2(n_388), .B(n_460), .C(n_462), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_531), .B(n_453), .Y(n_561) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_484), .B(n_479), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_513), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_513), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_498), .B(n_435), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_520), .B(n_435), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_505), .B(n_453), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_510), .B(n_460), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_518), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_497), .B(n_436), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_481), .B(n_462), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_519), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_529), .B(n_483), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_512), .B(n_463), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_539), .B(n_436), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_491), .B(n_480), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_514), .B(n_463), .Y(n_580) );
AOI322xp5_ASAP7_75t_L g581 ( .A1(n_490), .A2(n_458), .A3(n_470), .B1(n_480), .B2(n_472), .C1(n_471), .C2(n_449), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_522), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_525), .B(n_458), .Y(n_583) );
NAND2xp33_ASAP7_75t_L g584 ( .A(n_484), .B(n_464), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_509), .B(n_470), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_516), .B(n_472), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_493), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_489), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_493), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_540), .B(n_469), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_493), .B(n_388), .Y(n_591) );
OR2x6_ASAP7_75t_SL g592 ( .A(n_532), .B(n_471), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_544), .Y(n_593) );
AOI22xp5_ASAP7_75t_SL g594 ( .A1(n_546), .A2(n_489), .B1(n_496), .B2(n_492), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_547), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_542), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_584), .A2(n_492), .B1(n_487), .B2(n_496), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_556), .A2(n_533), .B1(n_523), .B2(n_494), .C(n_534), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_550), .B(n_537), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_581), .B(n_530), .C(n_519), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_577), .B(n_536), .Y(n_602) );
AOI21x1_ASAP7_75t_L g603 ( .A1(n_579), .A2(n_527), .B(n_385), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_551), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_565), .B(n_496), .Y(n_605) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_588), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_592), .A2(n_487), .B1(n_526), .B2(n_494), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_560), .A2(n_388), .B(n_536), .C(n_527), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_587), .B(n_526), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_565), .A2(n_527), .B(n_535), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_580), .B(n_528), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_548), .B(n_528), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_562), .A2(n_535), .B1(n_469), .B2(n_466), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_560), .B(n_517), .C(n_482), .Y(n_615) );
NOR3xp33_ASAP7_75t_SL g616 ( .A(n_562), .B(n_535), .C(n_373), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_543), .A2(n_482), .B1(n_517), .B2(n_473), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_556), .B(n_469), .C(n_466), .D(n_461), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_543), .A2(n_469), .B1(n_466), .B2(n_473), .Y(n_619) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_579), .A2(n_473), .B(n_461), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_558), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_588), .A2(n_387), .B(n_356), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_466), .B1(n_461), .B2(n_370), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_591), .A2(n_373), .B(n_370), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_590), .A2(n_370), .B1(n_363), .B2(n_362), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_573), .A2(n_363), .B1(n_364), .B2(n_362), .C(n_365), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_593), .Y(n_627) );
NAND2xp33_ASAP7_75t_L g628 ( .A(n_607), .B(n_553), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_608), .B(n_557), .C(n_563), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_594), .A2(n_552), .B1(n_567), .B2(n_561), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_597), .A2(n_554), .B1(n_545), .B2(n_563), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_620), .A2(n_564), .B(n_583), .Y(n_632) );
OAI322xp33_ASAP7_75t_SL g633 ( .A1(n_599), .A2(n_568), .A3(n_570), .B1(n_582), .B2(n_569), .C1(n_559), .C2(n_575), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_609), .A2(n_564), .B(n_586), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_614), .A2(n_572), .B1(n_576), .B2(n_566), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_598), .A2(n_585), .B(n_571), .C(n_578), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_596), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_605), .A2(n_574), .B1(n_363), .B2(n_362), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_618), .A2(n_363), .B1(n_362), .B2(n_365), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_606), .A2(n_339), .B(n_362), .C(n_360), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_606), .B(n_360), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_608), .A2(n_387), .B(n_356), .C(n_339), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_616), .B(n_364), .C(n_339), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_600), .B(n_362), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_624), .A2(n_365), .B(n_360), .C(n_368), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_602), .B(n_360), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_615), .A2(n_364), .B1(n_365), .B2(n_360), .C(n_374), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_623), .A2(n_366), .B1(n_377), .B2(n_374), .C(n_387), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_610), .A2(n_385), .B1(n_368), .B2(n_366), .C(n_377), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_617), .A2(n_387), .B(n_356), .C(n_364), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_626), .A2(n_364), .B(n_347), .C(n_377), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_625), .A2(n_364), .B(n_347), .C(n_374), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_622), .B(n_366), .C(n_374), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_612), .A2(n_368), .B1(n_364), .B2(n_352), .C(n_360), .Y(n_654) );
NOR3x1_ASAP7_75t_L g655 ( .A(n_595), .B(n_365), .C(n_368), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_601), .A2(n_364), .B1(n_365), .B2(n_368), .C(n_352), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_604), .A2(n_352), .B1(n_368), .B2(n_611), .C(n_621), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_636), .A2(n_630), .B1(n_631), .B2(n_637), .Y(n_659) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_642), .B(n_629), .C(n_651), .D(n_650), .E(n_639), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_644), .A2(n_634), .B(n_638), .C(n_647), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_628), .B(n_641), .C(n_640), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_635), .B(n_658), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_655), .B(n_652), .C(n_645), .D(n_643), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_659), .B(n_645), .C(n_648), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_663), .B(n_646), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_662), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_661), .B(n_632), .Y(n_668) );
NAND4xp75_ASAP7_75t_L g669 ( .A(n_668), .B(n_660), .C(n_664), .D(n_657), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_667), .B(n_627), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_669), .B(n_665), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_670), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_672), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_671), .B(n_666), .C(n_633), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_674), .A2(n_653), .B(n_649), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_603), .B(n_654), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_676), .B(n_619), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_656), .B1(n_368), .B2(n_352), .Y(n_678) );
endmodule