module real_jpeg_16148_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_0),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_0),
.A2(n_111),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_0),
.A2(n_111),
.B1(n_165),
.B2(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_0),
.A2(n_111),
.B1(n_446),
.B2(n_449),
.Y(n_445)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_2),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_88),
.Y(n_274)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_3),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_3),
.B(n_262),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_3),
.A2(n_171),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_3),
.A2(n_404),
.A3(n_406),
.B1(n_409),
.B2(n_414),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_3),
.A2(n_313),
.B1(n_428),
.B2(n_430),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_3),
.A2(n_108),
.B(n_274),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_161),
.B1(n_165),
.B2(n_170),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_4),
.A2(n_170),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_4),
.A2(n_170),
.B1(n_531),
.B2(n_533),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_5),
.A2(n_31),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_5),
.A2(n_31),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_5),
.A2(n_31),
.B1(n_474),
.B2(n_476),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_6),
.A2(n_291),
.B1(n_293),
.B2(n_295),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_6),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_6),
.A2(n_295),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_6),
.A2(n_295),
.B1(n_365),
.B2(n_389),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_6),
.A2(n_295),
.B1(n_434),
.B2(n_439),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_7),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_8),
.A2(n_210),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_8),
.A2(n_215),
.B1(n_539),
.B2(n_542),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_9),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_9),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_151),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_10),
.A2(n_155),
.B1(n_239),
.B2(n_244),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_10),
.A2(n_155),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_175),
.B1(n_177),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_179),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_13),
.A2(n_86),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_13),
.A2(n_86),
.B1(n_364),
.B2(n_367),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_13),
.A2(n_33),
.B1(n_86),
.B2(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_73),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_14),
.A2(n_73),
.B1(n_418),
.B2(n_419),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_14),
.A2(n_73),
.B1(n_108),
.B2(n_293),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_16),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g164 ( 
.A(n_16),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_517),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_296),
.B(n_515),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_248),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_22),
.B(n_248),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_184),
.Y(n_22)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_23),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_78),
.C(n_114),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_24),
.B(n_79),
.Y(n_250)
);

OAI22x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_37),
.B1(n_66),
.B2(n_67),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_26),
.A2(n_38),
.B1(n_255),
.B2(n_262),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_27),
.Y(n_405)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_28),
.Y(n_429)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_29),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_30),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_30),
.Y(n_272)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_35),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_35),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_36),
.Y(n_432)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_36),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_37),
.A2(n_66),
.B1(n_67),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_37),
.A2(n_66),
.B1(n_427),
.B2(n_433),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_37),
.A2(n_66),
.B1(n_433),
.B2(n_457),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_37),
.A2(n_66),
.B1(n_457),
.B2(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_38),
.A2(n_262),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_47),
.B(n_54),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_39),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_53),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_61),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_62),
.Y(n_327)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_62),
.Y(n_357)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_62),
.Y(n_479)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_66),
.Y(n_262)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_72),
.Y(n_442)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B1(n_107),
.B2(n_113),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_80),
.A2(n_90),
.B1(n_113),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_85),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_90),
.A2(n_107),
.B1(n_113),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_90),
.A2(n_113),
.B1(n_290),
.B2(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_90),
.A2(n_113),
.B1(n_231),
.B2(n_552),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_97),
.B(n_101),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_97),
.A2(n_265),
.B1(n_273),
.B2(n_275),
.Y(n_264)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_100),
.Y(n_269)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_110),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_113),
.B(n_313),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_115),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_159),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_116),
.A2(n_117),
.B1(n_159),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_139),
.B1(n_148),
.B2(n_150),
.Y(n_117)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_118),
.B(n_150),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_118),
.A2(n_148),
.B1(n_324),
.B2(n_328),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_118),
.A2(n_148),
.B1(n_328),
.B2(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_118),
.A2(n_148),
.B1(n_351),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_118),
.A2(n_148),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_127),
.Y(n_119)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_121),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_122),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_126),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B1(n_136),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_131),
.Y(n_408)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_139),
.Y(n_492)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_147),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_149),
.A2(n_187),
.B1(n_188),
.B2(n_195),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_149),
.B(n_313),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_149),
.A2(n_187),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_149),
.A2(n_187),
.B1(n_473),
.B2(n_492),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_157),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_158),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_158),
.Y(n_448)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_158),
.Y(n_544)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_159),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_171),
.B1(n_174),
.B2(n_180),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_160),
.A2(n_171),
.B1(n_280),
.B2(n_287),
.Y(n_279)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_164),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_169),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_205),
.B(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_171),
.A2(n_334),
.B1(n_339),
.B2(n_341),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_171),
.A2(n_363),
.B1(n_388),
.B2(n_394),
.Y(n_393)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_172),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_172),
.A2(n_223),
.B1(n_362),
.B2(n_372),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_175),
.Y(n_418)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_176),
.Y(n_286)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_176),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_180),
.Y(n_416)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_180),
.Y(n_465)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_217),
.B1(n_246),
.B2(n_247),
.Y(n_184)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_185),
.B(n_247),
.C(n_520),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_203),
.B1(n_204),
.B2(n_216),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_186),
.B(n_204),
.Y(n_547)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_194),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g537 ( 
.A(n_195),
.Y(n_537)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_196),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_198),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_202),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_203),
.A2(n_204),
.B1(n_550),
.B2(n_551),
.Y(n_549)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_229),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_218),
.B(n_523),
.C(n_524),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B(n_222),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_220),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_223),
.A2(n_342),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_223),
.A2(n_281),
.B1(n_417),
.B2(n_465),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_226),
.Y(n_394)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_227),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_230),
.Y(n_524)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_237),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_238),
.Y(n_528)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_242),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_249),
.B(n_251),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_253),
.B(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.C(n_288),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_254),
.A2(n_288),
.B1(n_289),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_254),
.Y(n_505)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_255),
.Y(n_494)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_263),
.B(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_279),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_264),
.B(n_279),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_272),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_305),
.A3(n_308),
.B1(n_312),
.B2(n_315),
.Y(n_304)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_499),
.B(n_513),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_484),
.B(n_498),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_452),
.B(n_483),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_399),
.B(n_451),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_359),
.B(n_398),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_332),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_303),
.B(n_332),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_322),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_304),
.A2(n_322),
.B1(n_323),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_313),
.B(n_382),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_313),
.B(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_347),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_333),
.B(n_349),
.C(n_358),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_358),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_375),
.B(n_397),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_373),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_373),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_392),
.B(n_396),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_387),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_395),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_400),
.B(n_401),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_424),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_402),
.B(n_425),
.C(n_444),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_415),
.B1(n_422),
.B2(n_423),
.Y(n_402)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_423),
.Y(n_470)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_415),
.Y(n_423)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_443),
.B2(n_444),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_482),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_482),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_468),
.B2(n_469),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_471),
.C(n_480),
.Y(n_497)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_462),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_463),
.C(n_467),
.Y(n_488)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_480),
.B2(n_481),
.Y(n_469)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_497),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_497),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_488),
.C(n_489),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_495),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_493),
.C(n_495),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_500),
.A2(n_502),
.B(n_509),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_502),
.C(n_514),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.C(n_508),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_503),
.B(n_512),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_508),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_511),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_554),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_519),
.B(n_521),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_546),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_527),
.A2(n_536),
.B(n_545),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_536),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_547),
.A2(n_548),
.B1(n_549),
.B2(n_553),
.Y(n_546)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_547),
.Y(n_553)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);


endmodule