module fake_aes_3442_n_584 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_154, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_584);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_584;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_524;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g156 ( .A(n_7), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_110), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_15), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_69), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_124), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_111), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_118), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_21), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_55), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_11), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_148), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_112), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_40), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_144), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_131), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_114), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_150), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_136), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_14), .Y(n_180) );
BUFx5_ASAP7_75t_L g181 ( .A(n_75), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_67), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_53), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_70), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_29), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_109), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_25), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_54), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_26), .Y(n_190) );
BUFx5_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_126), .B(n_116), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_138), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_120), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_72), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_44), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_128), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_18), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_45), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_33), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_122), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_56), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_139), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_94), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_119), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_133), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_8), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_90), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_91), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_121), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_113), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_58), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_146), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_130), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_48), .Y(n_220) );
NOR2xp67_ASAP7_75t_L g221 ( .A(n_62), .B(n_3), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_100), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_101), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_81), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_98), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_117), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_37), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_106), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_129), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_4), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_104), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_87), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_30), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_3), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_47), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_16), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_123), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_79), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_147), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_107), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_65), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_2), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_59), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_64), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_22), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g246 ( .A(n_88), .B(n_102), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_43), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_103), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_31), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_80), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_93), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_143), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_153), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_35), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_23), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_115), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_199), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_181), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_211), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_182), .B(n_0), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_242), .B(n_0), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_230), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_165), .B(n_1), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_156), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_195), .Y(n_269) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_158), .A2(n_99), .B(n_154), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_189), .B(n_1), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_202), .A2(n_220), .B1(n_194), .B2(n_213), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_160), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_163), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_225), .B(n_2), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_267), .B(n_171), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_269), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_263), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_257), .A2(n_256), .B1(n_255), .B2(n_254), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_260), .B(n_227), .Y(n_283) );
INVxp33_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_275), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_287), .B(n_240), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_285), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_287), .B(n_259), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_284), .B(n_265), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_276), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_280), .A2(n_272), .B1(n_271), .B2(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_278), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_283), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_282), .B(n_261), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_290), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_294), .B(n_157), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_297), .A2(n_281), .B(n_278), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_288), .B(n_279), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_292), .A2(n_266), .B(n_221), .C(n_168), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_295), .B(n_184), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_291), .B(n_159), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_296), .A2(n_270), .B(n_169), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_289), .B(n_196), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_293), .B(n_217), .Y(n_308) );
BUFx10_ASAP7_75t_L g309 ( .A(n_301), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_298), .B(n_167), .Y(n_310) );
OAI21xp5_ASAP7_75t_L g311 ( .A1(n_300), .A2(n_270), .B(n_174), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_307), .Y(n_312) );
BUFx8_ASAP7_75t_SL g313 ( .A(n_308), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_305), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_306), .A2(n_192), .B(n_176), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_299), .B(n_201), .Y(n_316) );
AND2x6_ASAP7_75t_L g317 ( .A(n_303), .B(n_172), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_304), .B(n_246), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_302), .A2(n_212), .B(n_180), .C(n_253), .Y(n_319) );
OAI21xp33_ASAP7_75t_L g320 ( .A1(n_298), .A2(n_252), .B(n_222), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_186), .B(n_183), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_298), .B(n_198), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_306), .A2(n_205), .B(n_200), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_298), .B(n_161), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_315), .A2(n_209), .B(n_208), .Y(n_326) );
OAI21x1_ASAP7_75t_SL g327 ( .A1(n_321), .A2(n_214), .B(n_210), .Y(n_327) );
BUFx10_ASAP7_75t_L g328 ( .A(n_314), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_324), .A2(n_219), .B(n_218), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_311), .A2(n_235), .B(n_231), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_316), .A2(n_237), .B(n_236), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_322), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_318), .B(n_241), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_323), .A2(n_245), .B(n_244), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_320), .B(n_162), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_317), .A2(n_181), .B1(n_191), .B2(n_204), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_325), .A2(n_250), .B(n_248), .Y(n_340) );
BUFx4_ASAP7_75t_SL g341 ( .A(n_313), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_319), .A2(n_251), .B(n_286), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_166), .B(n_164), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_309), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_324), .A2(n_191), .B(n_181), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_324), .A2(n_191), .B(n_181), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_311), .A2(n_191), .B(n_268), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_324), .A2(n_191), .B(n_216), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_322), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_311), .A2(n_268), .B(n_226), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_312), .A2(n_249), .B(n_247), .Y(n_356) );
CKINVDCx11_ASAP7_75t_R g357 ( .A(n_309), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_216), .B(n_226), .Y(n_358) );
AOI21x1_ASAP7_75t_L g359 ( .A1(n_311), .A2(n_226), .B(n_243), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_315), .A2(n_197), .B(n_233), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_355), .A2(n_4), .B(n_5), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_350), .B(n_5), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_358), .A2(n_6), .B(n_9), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_359), .A2(n_239), .B(n_232), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
INVx3_ASAP7_75t_SL g369 ( .A(n_354), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_341), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_351), .B(n_10), .Y(n_371) );
OA21x2_ASAP7_75t_L g372 ( .A1(n_352), .A2(n_229), .B(n_228), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_170), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_332), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_344), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_328), .B(n_224), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_338), .B(n_12), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_331), .B(n_356), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_348), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_330), .B(n_327), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_343), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_334), .B(n_223), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
BUFx5_ASAP7_75t_L g391 ( .A(n_334), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_336), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_342), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_337), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_326), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_360), .B(n_173), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_350), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_333), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_333), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_215), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_355), .A2(n_207), .B(n_206), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_350), .B(n_175), .Y(n_408) );
AOI21x1_ASAP7_75t_L g409 ( .A1(n_359), .A2(n_203), .B(n_193), .Y(n_409) );
AO21x1_ASAP7_75t_L g410 ( .A1(n_348), .A2(n_13), .B(n_17), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_333), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_350), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_333), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_333), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_346), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_415), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_177), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_391), .B(n_178), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_362), .B(n_179), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_401), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_412), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_363), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_397), .B1(n_382), .B2(n_391), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_414), .B(n_185), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_363), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_392), .A2(n_190), .B(n_188), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_364), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_375), .B(n_19), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_364), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_405), .B(n_187), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_414), .B(n_155), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_408), .B(n_20), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_406), .B(n_24), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_406), .B(n_27), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_28), .B1(n_32), .B2(n_34), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_411), .B(n_36), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_371), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_413), .B(n_38), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_413), .B(n_39), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_391), .B(n_41), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_391), .A2(n_42), .B1(n_46), .B2(n_49), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_368), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_368), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_384), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_384), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_390), .B(n_50), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_391), .B(n_51), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_385), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_377), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_392), .A2(n_52), .B(n_57), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_369), .B(n_60), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_388), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_403), .B(n_61), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_388), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_386), .Y(n_464) );
INVxp67_ASAP7_75t_R g465 ( .A(n_371), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_373), .B(n_152), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_378), .B(n_63), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_389), .B(n_66), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_450), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_449), .B(n_379), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_444), .B(n_416), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_429), .B(n_395), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_419), .B(n_393), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_421), .B(n_387), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_422), .B(n_376), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_424), .B(n_370), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_449), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_464), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_439), .B(n_383), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_437), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_456), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_452), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_464), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_461), .A2(n_361), .B(n_410), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_458), .B(n_394), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_454), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_444), .Y(n_494) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_465), .B(n_367), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_460), .B(n_372), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_445), .B(n_367), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_461), .B(n_463), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_417), .B(n_372), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_482), .B(n_457), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_471), .B(n_462), .Y(n_508) );
NOR2x1p5_ASAP7_75t_L g509 ( .A(n_504), .B(n_466), .Y(n_509) );
AOI211xp5_ASAP7_75t_SL g510 ( .A1(n_504), .A2(n_442), .B(n_467), .C(n_468), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_474), .B(n_425), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_476), .B(n_443), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_478), .B(n_463), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_472), .B(n_446), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_483), .B(n_436), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_502), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_494), .B(n_447), .Y(n_517) );
AND2x4_ASAP7_75t_SL g518 ( .A(n_470), .B(n_455), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_484), .B(n_453), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_490), .B(n_453), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_480), .B(n_470), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_498), .B(n_438), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_477), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_479), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_481), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_502), .B(n_459), .Y(n_526) );
NAND4xp25_ASAP7_75t_SL g527 ( .A(n_488), .B(n_426), .C(n_448), .D(n_420), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_469), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_469), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_523), .B(n_489), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_524), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_510), .A2(n_491), .B(n_495), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_525), .B(n_487), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_528), .B(n_493), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_511), .B(n_500), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_508), .B(n_497), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_530), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_513), .B(n_501), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_521), .B(n_505), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_516), .B(n_505), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_530), .B(n_503), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_522), .B(n_492), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_507), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g545 ( .A1(n_512), .A2(n_506), .B(n_428), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_531), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_532), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_533), .A2(n_509), .B1(n_517), .B2(n_518), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_544), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_544), .B(n_529), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_534), .Y(n_551) );
OAI31xp33_ASAP7_75t_L g552 ( .A1(n_537), .A2(n_527), .A3(n_526), .B(n_431), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_535), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_536), .B(n_519), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_539), .B(n_520), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_548), .A2(n_540), .B1(n_543), .B2(n_541), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_552), .A2(n_545), .B1(n_542), .B2(n_538), .C(n_496), .Y(n_557) );
AOI31xp33_ASAP7_75t_L g558 ( .A1(n_549), .A2(n_526), .A3(n_515), .B(n_442), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_546), .A2(n_499), .B(n_418), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_547), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_554), .A2(n_514), .B1(n_428), .B2(n_475), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_557), .A2(n_553), .B1(n_551), .B2(n_555), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_556), .A2(n_550), .B1(n_485), .B2(n_473), .Y(n_563) );
OAI211xp5_ASAP7_75t_SL g564 ( .A1(n_561), .A2(n_559), .B(n_560), .C(n_558), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_556), .A2(n_380), .B1(n_381), .B2(n_433), .Y(n_565) );
NAND3xp33_ASAP7_75t_SL g566 ( .A(n_562), .B(n_398), .C(n_459), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_563), .Y(n_567) );
NOR2xp33_ASAP7_75t_SL g568 ( .A(n_565), .B(n_409), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_567), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_566), .B(n_564), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_569), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_570), .A2(n_568), .B(n_365), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_572), .A2(n_407), .B1(n_71), .B2(n_73), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_571), .B(n_68), .Y(n_574) );
OAI22x1_ASAP7_75t_L g575 ( .A1(n_574), .A2(n_74), .B1(n_76), .B2(n_77), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_573), .Y(n_576) );
NOR2xp67_ASAP7_75t_L g577 ( .A(n_576), .B(n_575), .Y(n_577) );
OAI22x1_ASAP7_75t_SL g578 ( .A1(n_576), .A2(n_78), .B1(n_82), .B2(n_83), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_578), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_577), .A2(n_151), .B(n_85), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_84), .B(n_86), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_581), .B(n_579), .Y(n_582) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_149), .B(n_92), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_89), .B1(n_95), .B2(n_96), .Y(n_584) );
endmodule