module fake_netlist_6_348_n_181 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_181);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_181;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_14),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_53),
.B(n_46),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_21),
.B(n_23),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_45),
.B(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_52),
.B(n_47),
.C(n_49),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_52),
.B(n_2),
.C(n_5),
.Y(n_84)
);

CKINVDCx8_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_18),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_19),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_67),
.B(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_74),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_67),
.B(n_68),
.C(n_63),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_72),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_72),
.B1(n_66),
.B2(n_64),
.C(n_69),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_55),
.Y(n_98)
);

NOR2x1_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_59),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_55),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_71),
.B1(n_87),
.B2(n_86),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_86),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_78),
.B(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

OR2x6_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_93),
.B1(n_95),
.B2(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_93),
.Y(n_115)
);

OAI221xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_97),
.B1(n_91),
.B2(n_90),
.C(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_90),
.B(n_86),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_85),
.B(n_57),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_108),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_116),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_101),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_104),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_104),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_130),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_107),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_124),
.C(n_129),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_129),
.C(n_127),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_140),
.Y(n_146)
);

NOR3x1_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_124),
.C(n_85),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_129),
.B1(n_133),
.B2(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

OAI322xp33_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_82),
.A3(n_76),
.B1(n_11),
.B2(n_7),
.C1(n_8),
.C2(n_54),
.Y(n_150)
);

NOR3x1_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_57),
.C(n_54),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_137),
.B1(n_140),
.B2(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_138),
.B1(n_142),
.B2(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_139),
.B1(n_142),
.B2(n_107),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_132),
.B1(n_107),
.B2(n_71),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_131),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_132),
.B1(n_71),
.B2(n_76),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_82),
.C(n_54),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_12),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_25),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_59),
.B1(n_28),
.B2(n_31),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_71),
.C(n_26),
.Y(n_174)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_71),
.C(n_59),
.D(n_99),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_59),
.B1(n_71),
.B2(n_93),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_173),
.A2(n_165),
.B(n_164),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_168),
.B(n_163),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_169),
.B(n_166),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_172),
.B(n_162),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_177),
.B1(n_176),
.B2(n_178),
.C(n_59),
.Y(n_181)
);


endmodule