module fake_ibex_4_n_1127 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_132, n_174, n_210, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1127);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_132;
input n_174;
input n_210;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1127;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_1100;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_1080;
wire n_583;
wire n_887;
wire n_909;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_449;
wire n_547;
wire n_727;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_497;
wire n_243;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_1001;
wire n_944;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_433;
wire n_299;
wire n_262;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_1057;
wire n_1049;
wire n_763;
wire n_1086;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_397;
wire n_366;
wire n_894;
wire n_803;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_947;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_320;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_890;
wire n_816;
wire n_874;
wire n_912;
wire n_921;
wire n_1058;
wire n_1105;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_1000;
wire n_394;
wire n_984;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1038;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_42),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_82),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_84),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_93),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_65),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_120),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_59),
.Y(n_235)
);

BUFx2_ASAP7_75t_SL g236 ( 
.A(n_147),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_24),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_112),
.B(n_92),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_117),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_67),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_107),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_18),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_66),
.B(n_109),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_51),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_37),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_29),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_34),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_98),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_73),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_91),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_162),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_6),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_46),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_155),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_52),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_174),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_119),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_118),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_27),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_5),
.B(n_197),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_47),
.B(n_165),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_79),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_63),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_122),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_54),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_167),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_22),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_19),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_178),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_64),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_210),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_194),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_25),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_69),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_77),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_37),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_50),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_189),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_60),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_206),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_74),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_121),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_7),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_36),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_70),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_13),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_38),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_97),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_113),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_115),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_17),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_45),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_143),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_145),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_130),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_76),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_42),
.B(n_55),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_96),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_1),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_158),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_140),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_16),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_50),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_128),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_6),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_192),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_47),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_193),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_108),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_149),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_55),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_183),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_14),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_30),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_132),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_176),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_127),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_38),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_181),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_27),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_0),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_80),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_28),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_177),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_101),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_124),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_153),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_204),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_21),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_44),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_105),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_20),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_26),
.B(n_81),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_21),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_102),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_45),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_151),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_34),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_312),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_218),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_218),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_253),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_253),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_284),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_225),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_255),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_332),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_297),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_225),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_219),
.B(n_62),
.Y(n_386)
);

BUFx8_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_257),
.B(n_7),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_301),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_312),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_273),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_311),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_285),
.B(n_11),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_283),
.B(n_12),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_273),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_309),
.B(n_12),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_226),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_226),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_288),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_227),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_288),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_284),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_283),
.B(n_14),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_216),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_217),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_235),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_277),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_235),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_259),
.B(n_296),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_252),
.B(n_16),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_252),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_227),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_304),
.A2(n_106),
.B(n_209),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_328),
.B(n_17),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_304),
.Y(n_419)
);

BUFx8_ASAP7_75t_SL g420 ( 
.A(n_332),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_281),
.B(n_20),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_287),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_221),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_224),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_228),
.A2(n_111),
.B(n_208),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_231),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_232),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_233),
.A2(n_104),
.B(n_205),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_334),
.B(n_23),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_240),
.B(n_241),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_244),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_287),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_245),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_251),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_336),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_343),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_439)
);

OAI22x1_ASAP7_75t_SL g440 ( 
.A1(n_343),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_254),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_220),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_31),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_348),
.B(n_32),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_350),
.B(n_33),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_212),
.B(n_33),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_256),
.A2(n_126),
.B(n_202),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_258),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_350),
.B(n_35),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_260),
.A2(n_125),
.B(n_199),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_263),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_213),
.B(n_35),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_271),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_272),
.A2(n_123),
.B(n_196),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_413),
.B(n_278),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_416),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_222),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_413),
.B(n_279),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_396),
.B(n_292),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_407),
.B(n_289),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_396),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_375),
.B(n_315),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_406),
.B(n_223),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_SL g470 ( 
.A1(n_386),
.A2(n_237),
.B(n_230),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_387),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_386),
.A2(n_294),
.B1(n_292),
.B2(n_324),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_376),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_406),
.B(n_246),
.C(n_242),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

OAI22xp33_ASAP7_75t_L g477 ( 
.A1(n_370),
.A2(n_353),
.B1(n_249),
.B2(n_340),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_375),
.B(n_290),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_408),
.B(n_300),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_405),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_426),
.B(n_303),
.Y(n_486)
);

CKINVDCx6p67_ASAP7_75t_R g487 ( 
.A(n_405),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_423),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_448),
.A2(n_313),
.B(n_307),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_265),
.C(n_250),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_377),
.B(n_229),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_403),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx8_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_443),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_425),
.A2(n_344),
.B1(n_320),
.B2(n_280),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_432),
.B(n_314),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_415),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_387),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_371),
.B(n_286),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_372),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_322),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_383),
.B(n_236),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_370),
.A2(n_392),
.B1(n_394),
.B2(n_439),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_R g513 ( 
.A(n_387),
.B(n_294),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_399),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_372),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_388),
.B(n_331),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

BUFx8_ASAP7_75t_SL g520 ( 
.A(n_420),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_376),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_418),
.B(n_234),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_452),
.B(n_425),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_399),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_410),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_402),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_372),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_386),
.A2(n_338),
.B1(n_324),
.B2(n_299),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_383),
.B(n_326),
.C(n_360),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_404),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_437),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_379),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_379),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_454),
.B(n_323),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_387),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_L g540 ( 
.A1(n_428),
.A2(n_308),
.B(n_293),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_316),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_376),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_446),
.B(n_450),
.C(n_440),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_380),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_400),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_400),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_378),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_429),
.A2(n_435),
.B1(n_449),
.B2(n_436),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_428),
.B(n_327),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_429),
.A2(n_351),
.B1(n_361),
.B2(n_220),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_435),
.B(n_282),
.Y(n_552)
);

INVx8_ASAP7_75t_L g553 ( 
.A(n_450),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_392),
.A2(n_268),
.B1(n_266),
.B2(n_365),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_SL g555 ( 
.A1(n_435),
.A2(n_364),
.B(n_333),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_401),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

BUFx6f_ASAP7_75t_SL g558 ( 
.A(n_373),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_401),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_436),
.B(n_329),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_389),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_436),
.A2(n_342),
.B1(n_367),
.B2(n_220),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_442),
.B(n_282),
.Y(n_563)
);

AO21x2_ASAP7_75t_L g564 ( 
.A1(n_427),
.A2(n_337),
.B(n_335),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_394),
.A2(n_269),
.B1(n_352),
.B2(n_357),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_442),
.B(n_339),
.Y(n_566)
);

OA22x2_ASAP7_75t_L g567 ( 
.A1(n_439),
.A2(n_352),
.B1(n_325),
.B2(n_330),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_380),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_409),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_409),
.Y(n_570)
);

OAI22x1_ASAP7_75t_L g571 ( 
.A1(n_434),
.A2(n_325),
.B1(n_358),
.B2(n_357),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_417),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_395),
.B(n_220),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_442),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_414),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_539),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_538),
.B(n_449),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_557),
.B(n_354),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_461),
.A2(n_444),
.B1(n_445),
.B2(n_421),
.Y(n_580)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_464),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_466),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_513),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_574),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_468),
.A2(n_358),
.B1(n_362),
.B2(n_306),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_385),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_494),
.B(n_373),
.Y(n_587)
);

AO22x1_ASAP7_75t_L g588 ( 
.A1(n_529),
.A2(n_317),
.B1(n_215),
.B2(n_239),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_461),
.B(n_419),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_419),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_463),
.B(n_341),
.Y(n_591)
);

AND2x6_ASAP7_75t_SL g592 ( 
.A(n_510),
.B(n_520),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_468),
.A2(n_424),
.B1(n_274),
.B2(n_275),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_457),
.B(n_381),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_467),
.B(n_522),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_512),
.A2(n_424),
.B(n_382),
.C(n_391),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_458),
.B(n_214),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_497),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_518),
.B(n_384),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_495),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_390),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_463),
.B(n_345),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_480),
.B(n_390),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_480),
.B(n_391),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_502),
.B(n_427),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_501),
.B(n_243),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_472),
.A2(n_363),
.B1(n_342),
.B2(n_298),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_516),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_501),
.B(n_247),
.Y(n_614)
);

NOR2x1_ASAP7_75t_L g615 ( 
.A(n_492),
.B(n_490),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_545),
.Y(n_617)
);

O2A1O1Ixp5_ASAP7_75t_L g618 ( 
.A1(n_535),
.A2(n_359),
.B(n_356),
.C(n_355),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_459),
.B(n_291),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_530),
.B(n_417),
.Y(n_620)
);

AND2x4_ASAP7_75t_SL g621 ( 
.A(n_471),
.B(n_298),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_573),
.B(n_261),
.Y(n_622)
);

OAI22x1_ASAP7_75t_R g623 ( 
.A1(n_471),
.A2(n_368),
.B1(n_347),
.B2(n_264),
.Y(n_623)
);

OAI22xp33_ASAP7_75t_L g624 ( 
.A1(n_510),
.A2(n_363),
.B1(n_342),
.B2(n_367),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_519),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_552),
.B(n_448),
.C(n_451),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_520),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_459),
.B(n_295),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_527),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_510),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_477),
.A2(n_363),
.B1(n_367),
.B2(n_342),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_459),
.B(n_346),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_469),
.B(n_262),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_531),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_572),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_476),
.B(n_267),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_456),
.B(n_270),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_481),
.B(n_276),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_484),
.B(n_448),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_545),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_568),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_534),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_567),
.A2(n_298),
.B1(n_363),
.B2(n_367),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_507),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_565),
.B(n_451),
.C(n_448),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_553),
.B(n_302),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_460),
.B(n_451),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_553),
.A2(n_455),
.B1(n_430),
.B2(n_451),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_550),
.B(n_305),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_553),
.B(n_310),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_567),
.A2(n_319),
.B1(n_366),
.B2(n_248),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_571),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_506),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_550),
.B(n_430),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_540),
.A2(n_455),
.B1(n_238),
.B2(n_41),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_508),
.B(n_68),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_487),
.Y(n_662)
);

INVxp33_ASAP7_75t_SL g663 ( 
.A(n_504),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_71),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_473),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_535),
.B(n_72),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_523),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_477),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_572),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_500),
.B(n_75),
.Y(n_670)
);

BUFx5_ASAP7_75t_L g671 ( 
.A(n_546),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_465),
.B(n_482),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_542),
.B(n_78),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_465),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_486),
.B(n_46),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_555),
.B(n_142),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_542),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_493),
.B(n_49),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_462),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_541),
.B(n_53),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_560),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_493),
.B(n_56),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_537),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_544),
.B(n_58),
.Y(n_686)
);

AOI221xp5_ASAP7_75t_L g687 ( 
.A1(n_554),
.A2(n_211),
.B1(n_83),
.B2(n_85),
.C(n_87),
.Y(n_687)
);

BUFx8_ASAP7_75t_L g688 ( 
.A(n_558),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_556),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_504),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_500),
.B(n_94),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_559),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_649),
.A2(n_572),
.B(n_564),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_594),
.B(n_569),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_671),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_598),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_646),
.A2(n_489),
.B(n_560),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_581),
.B(n_570),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_612),
.B(n_558),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_587),
.A2(n_536),
.B(n_533),
.C(n_575),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_632),
.A2(n_566),
.B(n_576),
.C(n_551),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_601),
.B(n_485),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_578),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_582),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_601),
.B(n_473),
.Y(n_705)
);

OR2x6_ASAP7_75t_SL g706 ( 
.A(n_628),
.B(n_576),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_610),
.B(n_526),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_640),
.A2(n_526),
.B(n_483),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_595),
.B(n_479),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_644),
.A2(n_562),
.B1(n_479),
.B2(n_491),
.Y(n_710)
);

NAND2x1_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_478),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_671),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_636),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_621),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_611),
.A2(n_524),
.B1(n_491),
.B2(n_488),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_599),
.B(n_491),
.Y(n_716)
);

BUFx8_ASAP7_75t_L g717 ( 
.A(n_631),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_688),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_688),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_672),
.A2(n_491),
.B(n_524),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_632),
.A2(n_514),
.B(n_517),
.C(n_525),
.Y(n_721)
);

OR2x6_ASAP7_75t_SL g722 ( 
.A(n_583),
.B(n_99),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_627),
.B(n_524),
.Y(n_723)
);

OAI21xp33_ASAP7_75t_L g724 ( 
.A1(n_580),
.A2(n_525),
.B(n_498),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_650),
.A2(n_620),
.B(n_664),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_585),
.B(n_103),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_597),
.B(n_116),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_606),
.A2(n_607),
.B(n_639),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_647),
.B(n_129),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_596),
.A2(n_511),
.B(n_505),
.C(n_499),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_685),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_655),
.B(n_131),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_656),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_591),
.B(n_604),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_657),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_648),
.B(n_133),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_680),
.A2(n_543),
.B1(n_561),
.B2(n_548),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_636),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_591),
.B(n_134),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_605),
.A2(n_630),
.B(n_613),
.C(n_625),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_579),
.B(n_137),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_669),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_591),
.B(n_138),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_652),
.B(n_148),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_657),
.B(n_665),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_653),
.A2(n_521),
.B1(n_474),
.B2(n_543),
.C(n_169),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_604),
.B(n_150),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_SL g749 ( 
.A(n_687),
.B(n_157),
.C(n_166),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_604),
.B(n_170),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_678),
.A2(n_474),
.B1(n_175),
.B2(n_179),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_667),
.A2(n_172),
.B(n_182),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_684),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_635),
.B(n_643),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_616),
.B(n_195),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_690),
.B(n_191),
.Y(n_756)
);

BUFx2_ASAP7_75t_SL g757 ( 
.A(n_662),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_602),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_619),
.B(n_629),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_577),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_651),
.A2(n_589),
.B(n_590),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_623),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_633),
.B(n_651),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_686),
.B(n_654),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_577),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_586),
.A2(n_589),
.B(n_590),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_675),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_660),
.A2(n_677),
.B(n_586),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_681),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_615),
.A2(n_682),
.B1(n_631),
.B2(n_638),
.Y(n_770)
);

AND2x2_ASAP7_75t_SL g771 ( 
.A(n_663),
.B(n_666),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_685),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_L g773 ( 
.A1(n_593),
.A2(n_614),
.B(n_609),
.Y(n_773)
);

CKINVDCx11_ASAP7_75t_R g774 ( 
.A(n_592),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_624),
.A2(n_637),
.B1(n_634),
.B2(n_584),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_689),
.B(n_692),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_659),
.A2(n_676),
.B1(n_674),
.B2(n_668),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_645),
.B(n_665),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_668),
.A2(n_683),
.B1(n_679),
.B2(n_600),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_645),
.A2(n_642),
.B1(n_641),
.B2(n_617),
.Y(n_780)
);

CKINVDCx6p67_ASAP7_75t_R g781 ( 
.A(n_670),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_661),
.A2(n_666),
.B1(n_673),
.B2(n_691),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_673),
.B(n_466),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_649),
.A2(n_640),
.B(n_658),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_587),
.A2(n_470),
.B(n_596),
.C(n_603),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_662),
.B(n_598),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_649),
.A2(n_640),
.B(n_658),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_588),
.B(n_529),
.C(n_512),
.Y(n_788)
);

O2A1O1Ixp5_ASAP7_75t_L g789 ( 
.A1(n_618),
.A2(n_658),
.B(n_608),
.C(n_535),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_628),
.Y(n_790)
);

NOR2x1_ASAP7_75t_SL g791 ( 
.A(n_757),
.B(n_703),
.Y(n_791)
);

NAND3x1_ASAP7_75t_L g792 ( 
.A(n_788),
.B(n_774),
.C(n_706),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_758),
.B(n_694),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_771),
.A2(n_785),
.B1(n_754),
.B2(n_776),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_769),
.B(n_759),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_735),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_779),
.A2(n_741),
.B1(n_777),
.B2(n_783),
.Y(n_797)
);

AOI221xp5_ASAP7_75t_SL g798 ( 
.A1(n_777),
.A2(n_779),
.B1(n_773),
.B2(n_728),
.C(n_738),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_767),
.B(n_733),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_763),
.B(n_770),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_768),
.B(n_761),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_718),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_768),
.A2(n_725),
.B1(n_782),
.B2(n_745),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_789),
.A2(n_697),
.B(n_766),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_705),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_747),
.B(n_725),
.C(n_715),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_762),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_716),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_699),
.B(n_702),
.Y(n_811)
);

AOI21xp33_ASAP7_75t_L g812 ( 
.A1(n_738),
.A2(n_753),
.B(n_751),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_790),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_708),
.A2(n_743),
.B(n_739),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_786),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_SL g816 ( 
.A(n_722),
.B(n_727),
.C(n_717),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_756),
.B(n_760),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_753),
.A2(n_749),
.B(n_737),
.Y(n_818)
);

BUFx4f_ASAP7_75t_SL g819 ( 
.A(n_717),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_786),
.B(n_696),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_780),
.Y(n_821)
);

BUFx2_ASAP7_75t_SL g822 ( 
.A(n_736),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_765),
.B(n_736),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_721),
.A2(n_742),
.B(n_701),
.C(n_700),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_SL g825 ( 
.A1(n_713),
.A2(n_739),
.B(n_751),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_775),
.B(n_726),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_739),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_764),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_734),
.A2(n_781),
.B1(n_729),
.B2(n_732),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_719),
.B(n_723),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_755),
.A2(n_709),
.B1(n_710),
.B2(n_707),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_695),
.B(n_712),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_752),
.A2(n_720),
.B(n_744),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_724),
.A2(n_730),
.B(n_772),
.C(n_731),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_740),
.A2(n_750),
.B(n_748),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_778),
.B(n_746),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_711),
.A2(n_789),
.B(n_787),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_704),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_725),
.A2(n_697),
.B(n_626),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_747),
.B(n_788),
.C(n_646),
.Y(n_840)
);

NAND2x1p5_ASAP7_75t_L g841 ( 
.A(n_714),
.B(n_598),
.Y(n_841)
);

OA21x2_ASAP7_75t_L g842 ( 
.A1(n_725),
.A2(n_697),
.B(n_626),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_758),
.B(n_466),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_704),
.Y(n_844)
);

AO31x2_ASAP7_75t_L g845 ( 
.A1(n_693),
.A2(n_784),
.A3(n_787),
.B(n_785),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_788),
.A2(n_779),
.B1(n_470),
.B2(n_611),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_718),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_769),
.B(n_581),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_758),
.B(n_466),
.Y(n_849)
);

OA21x2_ASAP7_75t_L g850 ( 
.A1(n_725),
.A2(n_697),
.B(n_626),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_718),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_758),
.B(n_466),
.Y(n_852)
);

AO21x2_ASAP7_75t_L g853 ( 
.A1(n_725),
.A2(n_697),
.B(n_693),
.Y(n_853)
);

NAND3x1_ASAP7_75t_L g854 ( 
.A(n_788),
.B(n_394),
.C(n_530),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_736),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_714),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_714),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_758),
.B(n_703),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_736),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_706),
.Y(n_860)
);

BUFx12f_ASAP7_75t_L g861 ( 
.A(n_718),
.Y(n_861)
);

OA22x2_ASAP7_75t_L g862 ( 
.A1(n_762),
.A2(n_472),
.B1(n_529),
.B2(n_510),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_789),
.A2(n_787),
.B(n_784),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_757),
.B(n_553),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_779),
.A2(n_529),
.B1(n_788),
.B2(n_611),
.Y(n_865)
);

AO32x2_ASAP7_75t_L g866 ( 
.A1(n_779),
.A2(n_777),
.A3(n_738),
.B1(n_753),
.B2(n_611),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_466),
.Y(n_867)
);

OAI22x1_ASAP7_75t_L g868 ( 
.A1(n_762),
.A2(n_472),
.B1(n_434),
.B2(n_422),
.Y(n_868)
);

OA21x2_ASAP7_75t_L g869 ( 
.A1(n_725),
.A2(n_697),
.B(n_626),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_789),
.A2(n_787),
.B(n_784),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_725),
.A2(n_697),
.B(n_693),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_762),
.B(n_457),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_758),
.B(n_466),
.Y(n_873)
);

CKINVDCx8_ASAP7_75t_R g874 ( 
.A(n_718),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_SL g875 ( 
.A1(n_779),
.A2(n_218),
.B(n_374),
.C(n_373),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_714),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_779),
.B(n_470),
.C(n_788),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_758),
.B(n_466),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_718),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_718),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_762),
.B(n_457),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_698),
.B(n_594),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_758),
.B(n_466),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_789),
.A2(n_787),
.B(n_784),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_747),
.B(n_788),
.C(n_646),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_706),
.Y(n_886)
);

AO31x2_ASAP7_75t_L g887 ( 
.A1(n_693),
.A2(n_784),
.A3(n_787),
.B(n_785),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_758),
.B(n_466),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_714),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_704),
.Y(n_890)
);

AOI21xp33_ASAP7_75t_L g891 ( 
.A1(n_777),
.A2(n_738),
.B(n_779),
.Y(n_891)
);

BUFx4f_ASAP7_75t_L g892 ( 
.A(n_762),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_789),
.A2(n_787),
.B(n_784),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_703),
.B(n_758),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_788),
.B(n_513),
.C(n_504),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_706),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_758),
.B(n_466),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_844),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_845),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_793),
.B(n_882),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_843),
.B(n_849),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_819),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_815),
.B(n_802),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_890),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_801),
.B(n_862),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_858),
.B(n_800),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_877),
.A2(n_865),
.B1(n_891),
.B2(n_846),
.Y(n_907)
);

AO21x2_ASAP7_75t_L g908 ( 
.A1(n_891),
.A2(n_806),
.B(n_812),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_864),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_845),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_852),
.B(n_867),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_SL g912 ( 
.A(n_816),
.B(n_846),
.C(n_813),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_873),
.B(n_878),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_798),
.B(n_875),
.C(n_797),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_883),
.B(n_888),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_863),
.A2(n_884),
.B(n_893),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_897),
.B(n_795),
.Y(n_917)
);

BUFx10_ASAP7_75t_L g918 ( 
.A(n_864),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_864),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_870),
.A2(n_833),
.B(n_806),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_872),
.B(n_881),
.Y(n_921)
);

AO21x2_ASAP7_75t_L g922 ( 
.A1(n_812),
.A2(n_840),
.B(n_885),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_840),
.A2(n_885),
.B(n_826),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_799),
.B(n_848),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_887),
.Y(n_925)
);

AO21x1_ASAP7_75t_SL g926 ( 
.A1(n_894),
.A2(n_810),
.B(n_796),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_887),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_791),
.B(n_894),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_837),
.A2(n_835),
.B(n_803),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_803),
.A2(n_814),
.B(n_825),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_802),
.B(n_815),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_854),
.B(n_807),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_860),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_820),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_818),
.A2(n_805),
.B(n_824),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_841),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_855),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_821),
.B(n_811),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_830),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_886),
.B(n_896),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_808),
.A2(n_834),
.B(n_805),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_855),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_866),
.B(n_794),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_828),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_839),
.A2(n_842),
.B(n_869),
.Y(n_945)
);

AOI21x1_ASAP7_75t_L g946 ( 
.A1(n_829),
.A2(n_869),
.B(n_850),
.Y(n_946)
);

AOI21xp33_ASAP7_75t_SL g947 ( 
.A1(n_868),
.A2(n_804),
.B(n_809),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_879),
.B(n_880),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_823),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_817),
.B(n_857),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_829),
.A2(n_836),
.B(n_832),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_855),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_822),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_847),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_856),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_853),
.A2(n_871),
.B(n_831),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_859),
.A2(n_831),
.B(n_871),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_827),
.Y(n_958)
);

OA21x2_ASAP7_75t_L g959 ( 
.A1(n_853),
.A2(n_866),
.B(n_889),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_866),
.A2(n_876),
.B(n_895),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_792),
.A2(n_892),
.B1(n_851),
.B2(n_861),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_892),
.A2(n_851),
.B(n_874),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_858),
.B(n_791),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_858),
.B(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_793),
.B(n_882),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_793),
.B(n_882),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_838),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_864),
.Y(n_968)
);

INVx4_ASAP7_75t_SL g969 ( 
.A(n_928),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_902),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_899),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_907),
.B(n_935),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_902),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_928),
.Y(n_974)
);

INVx11_ASAP7_75t_L g975 ( 
.A(n_948),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_934),
.B(n_965),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_943),
.B(n_907),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_910),
.Y(n_978)
);

INVxp67_ASAP7_75t_SL g979 ( 
.A(n_916),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_910),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_906),
.B(n_900),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_906),
.B(n_900),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_925),
.Y(n_983)
);

AO21x1_ASAP7_75t_SL g984 ( 
.A1(n_926),
.A2(n_958),
.B(n_952),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_927),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_934),
.B(n_966),
.Y(n_986)
);

AO21x2_ASAP7_75t_L g987 ( 
.A1(n_941),
.A2(n_923),
.B(n_914),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_943),
.B(n_908),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_929),
.A2(n_938),
.B(n_905),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_963),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_957),
.B(n_951),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_964),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_898),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_964),
.Y(n_994)
);

NOR2xp67_ASAP7_75t_L g995 ( 
.A(n_912),
.B(n_919),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_929),
.A2(n_905),
.B(n_920),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_904),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_903),
.Y(n_999)
);

OR2x2_ASAP7_75t_SL g1000 ( 
.A(n_962),
.B(n_960),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_967),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_977),
.B(n_959),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_977),
.B(n_922),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_977),
.B(n_922),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_976),
.B(n_959),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_972),
.B(n_908),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_976),
.B(n_932),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_988),
.B(n_945),
.Y(n_1008)
);

CKINVDCx6p67_ASAP7_75t_R g1009 ( 
.A(n_999),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_988),
.B(n_956),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_996),
.B(n_969),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_986),
.B(n_921),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_SL g1013 ( 
.A(n_999),
.B(n_962),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_971),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_969),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_969),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_978),
.B(n_946),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_980),
.B(n_960),
.Y(n_1018)
);

OAI31xp33_ASAP7_75t_L g1019 ( 
.A1(n_999),
.A2(n_917),
.A3(n_901),
.B(n_911),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_980),
.B(n_983),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_983),
.B(n_930),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1002),
.B(n_979),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1003),
.B(n_1004),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1002),
.B(n_979),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1002),
.B(n_1008),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1014),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1014),
.Y(n_1027)
);

NAND2x1_ASAP7_75t_L g1028 ( 
.A(n_1015),
.B(n_990),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_1015),
.B(n_974),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1008),
.B(n_1017),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_1019),
.B(n_995),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1008),
.B(n_985),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1011),
.B(n_991),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1020),
.B(n_989),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_SL g1037 ( 
.A(n_1015),
.B(n_984),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1004),
.B(n_987),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1025),
.B(n_1018),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_1018),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_1030),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1031),
.B(n_1018),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1031),
.B(n_1021),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_1021),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1032),
.A2(n_1019),
.B1(n_982),
.B2(n_981),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1023),
.B(n_1006),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1022),
.B(n_1021),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1026),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1022),
.B(n_1010),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1023),
.B(n_1006),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_1029),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1022),
.B(n_1010),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1026),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1029),
.B(n_1033),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1027),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1033),
.B(n_1010),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_1056),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1051),
.B(n_1036),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1051),
.B(n_1036),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_1054),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_1047),
.B(n_1015),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1048),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1048),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1053),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1039),
.B(n_1024),
.Y(n_1066)
);

AO221x1_ASAP7_75t_L g1067 ( 
.A1(n_1041),
.A2(n_1037),
.B1(n_992),
.B2(n_990),
.C(n_994),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1056),
.B(n_1034),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_1041),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1055),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1039),
.B(n_1024),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1062),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1057),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_1069),
.B(n_1045),
.C(n_1046),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1057),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1061),
.A2(n_1045),
.B(n_995),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1060),
.Y(n_1077)
);

OR3x2_ASAP7_75t_L g1078 ( 
.A(n_1067),
.B(n_975),
.C(n_940),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1058),
.B(n_1046),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1065),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1067),
.A2(n_1050),
.B1(n_1052),
.B2(n_1049),
.Y(n_1081)
);

NOR4xp25_ASAP7_75t_L g1082 ( 
.A(n_1059),
.B(n_997),
.C(n_993),
.D(n_1001),
.Y(n_1082)
);

AOI32xp33_ASAP7_75t_L g1083 ( 
.A1(n_1071),
.A2(n_1044),
.A3(n_1040),
.B1(n_1049),
.B2(n_1052),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1062),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1066),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1083),
.A2(n_1074),
.B1(n_1079),
.B2(n_1082),
.C(n_1077),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_1076),
.A2(n_933),
.B(n_1013),
.Y(n_1087)
);

OAI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_1081),
.A2(n_1061),
.B1(n_1050),
.B2(n_1068),
.C(n_947),
.Y(n_1088)
);

AOI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1078),
.A2(n_1016),
.B(n_961),
.C(n_1013),
.Y(n_1089)
);

AOI322xp5_ASAP7_75t_L g1090 ( 
.A1(n_1079),
.A2(n_1071),
.A3(n_1066),
.B1(n_1042),
.B2(n_1040),
.C1(n_1044),
.C2(n_1043),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1078),
.A2(n_1073),
.B1(n_1075),
.B2(n_1085),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1080),
.A2(n_948),
.B(n_954),
.C(n_919),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1072),
.B(n_1042),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_975),
.B1(n_1009),
.B2(n_1016),
.Y(n_1094)
);

AOI211xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1086),
.A2(n_998),
.B(n_1012),
.C(n_990),
.Y(n_1095)
);

NAND4xp25_ASAP7_75t_SL g1096 ( 
.A(n_1090),
.B(n_1037),
.C(n_1044),
.D(n_1043),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_1088),
.A2(n_1084),
.B1(n_1072),
.B2(n_1070),
.C(n_1065),
.Y(n_1097)
);

AOI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_1092),
.A2(n_1084),
.B1(n_1070),
.B2(n_1038),
.C(n_1064),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1089),
.A2(n_1028),
.B(n_1047),
.C(n_1035),
.Y(n_1099)
);

OAI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_1087),
.A2(n_1038),
.B1(n_948),
.B2(n_1063),
.C(n_1064),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_1093),
.B(n_970),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1095),
.A2(n_1028),
.B(n_1035),
.C(n_973),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_1096),
.B(n_970),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1100),
.B(n_968),
.C(n_909),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_1097),
.B(n_1030),
.C(n_903),
.Y(n_1105)
);

AND4x1_ASAP7_75t_L g1106 ( 
.A(n_1099),
.B(n_970),
.C(n_962),
.D(n_953),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_1098),
.B(n_944),
.C(n_993),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1103),
.B(n_1094),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_1105),
.B(n_1101),
.C(n_950),
.Y(n_1109)
);

NAND5xp2_ASAP7_75t_L g1110 ( 
.A(n_1102),
.B(n_1030),
.C(n_982),
.D(n_981),
.E(n_939),
.Y(n_1110)
);

AOI211xp5_ASAP7_75t_SL g1111 ( 
.A1(n_1104),
.A2(n_998),
.B(n_924),
.C(n_955),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1107),
.B(n_1063),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1106),
.B(n_1007),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1111),
.B(n_1055),
.Y(n_1114)
);

AND3x1_ASAP7_75t_L g1115 ( 
.A(n_1109),
.B(n_998),
.C(n_992),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1110),
.B(n_949),
.C(n_913),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1108),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_L g1118 ( 
.A(n_1113),
.B(n_931),
.Y(n_1118)
);

XNOR2x1_ASAP7_75t_L g1119 ( 
.A(n_1117),
.B(n_1112),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1115),
.B(n_1113),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_1118),
.B1(n_1114),
.B2(n_1116),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1121),
.A2(n_1119),
.B(n_931),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1122),
.A2(n_936),
.B1(n_931),
.B2(n_1016),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_998),
.B(n_915),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_1125),
.B(n_936),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1126),
.A2(n_942),
.B(n_937),
.Y(n_1127)
);


endmodule