module fake_netlist_6_4667_n_1861 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1861);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1861;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_20),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_50),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_143),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_71),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_104),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_109),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g210 ( 
.A(n_126),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_98),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_96),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_94),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_15),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_90),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_18),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_119),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_56),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_112),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_54),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_75),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_38),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_176),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_12),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_47),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_92),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_108),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_138),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_35),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_19),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_64),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_59),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_54),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_86),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_106),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_77),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

INVxp33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_51),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_148),
.Y(n_278)
);

BUFx8_ASAP7_75t_SL g279 ( 
.A(n_118),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_137),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_95),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_125),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_113),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_83),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_159),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_123),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_156),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_107),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_58),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_76),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_183),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_88),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_101),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_161),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_155),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_172),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_8),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_169),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_145),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_61),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_51),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_43),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_182),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_91),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_129),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_19),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_52),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_164),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_166),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_173),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_116),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_55),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_33),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_163),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_150),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_79),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_135),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_67),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_53),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_11),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_8),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_72),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_57),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_144),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_102),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_34),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_24),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_30),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_46),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_99),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_185),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_66),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_7),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_35),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_70),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_84),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_21),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_122),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_187),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_42),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_23),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_58),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_100),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_50),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_32),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_46),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_165),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_45),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_44),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_117),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_82),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_23),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_87),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_186),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_9),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_44),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_254),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_254),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_254),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_291),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_274),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_279),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_274),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_243),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_192),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_280),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_337),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_237),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_193),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_192),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_195),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_204),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_239),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_240),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_248),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_251),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_241),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_326),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_196),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_252),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_255),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_259),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_269),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_270),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_244),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_288),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_292),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_202),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_294),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_265),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_314),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_278),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_216),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_217),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_268),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_196),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_285),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_197),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_287),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_216),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_303),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_267),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_235),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_235),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_249),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_249),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_303),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_321),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_198),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_321),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_328),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_328),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_221),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_221),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_289),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_266),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_266),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_226),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_336),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_336),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_295),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_268),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_299),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_267),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_194),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_307),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_199),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_197),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_228),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_198),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_203),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_214),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_282),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_387),
.B(n_191),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_401),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_391),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_282),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_322),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_400),
.B(n_191),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_376),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_408),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_218),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_322),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_411),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g493 ( 
.A1(n_446),
.A2(n_219),
.B(n_215),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_200),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_447),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_423),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_378),
.A2(n_338),
.B1(n_340),
.B2(n_260),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_415),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_450),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_418),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_198),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_458),
.B(n_224),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_453),
.B(n_267),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_229),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_379),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_232),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_383),
.A2(n_272),
.B1(n_370),
.B2(n_363),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_451),
.A2(n_462),
.B1(n_220),
.B2(n_223),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_394),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_464),
.A2(n_245),
.B(n_233),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_395),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_395),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_429),
.B(n_191),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_460),
.B(n_258),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_432),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_385),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_464),
.B(n_261),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_381),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_381),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_448),
.B(n_352),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_382),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_389),
.B(n_390),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_390),
.B(n_263),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_382),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_384),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_384),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_514),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_468),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_473),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_386),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_480),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_472),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_503),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_510),
.B(n_386),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_525),
.A2(n_283),
.B(n_276),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_470),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_510),
.A2(n_402),
.B1(n_431),
.B2(n_427),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_503),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_541),
.C(n_475),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_474),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_473),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_290),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_473),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_474),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_466),
.B(n_454),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_505),
.B(n_456),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_388),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_466),
.A2(n_431),
.B1(n_402),
.B2(n_461),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_477),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_503),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_475),
.B(n_459),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_482),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_483),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_483),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_503),
.B(n_210),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_514),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_SL g586 ( 
.A(n_508),
.B(n_393),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_505),
.B(n_380),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_484),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_484),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_473),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_525),
.A2(n_296),
.B(n_293),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_486),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_476),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_476),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_483),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_486),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_467),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_479),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_492),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_494),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_532),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_486),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_519),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_519),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_523),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_487),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_506),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_481),
.B(n_392),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_532),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_509),
.B(n_207),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_476),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_516),
.B(n_388),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_503),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_503),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_504),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_526),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_491),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_525),
.A2(n_206),
.B(n_297),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

AND3x2_ASAP7_75t_L g638 ( 
.A(n_516),
.B(n_300),
.C(n_298),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_511),
.A2(n_425),
.B1(n_424),
.B2(n_267),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_499),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_476),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_471),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_517),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_522),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_517),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_491),
.Y(n_648)
);

CKINVDCx6p67_ASAP7_75t_R g649 ( 
.A(n_471),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_527),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_527),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_511),
.B(n_201),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_511),
.B(n_311),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_530),
.B(n_207),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_533),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_511),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_533),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_511),
.B(n_313),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_520),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_485),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_520),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_534),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_520),
.B(n_436),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_531),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_520),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_478),
.A2(n_306),
.B(n_301),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_534),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_316),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_529),
.A2(n_267),
.B1(n_410),
.B2(n_397),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_501),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_488),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_501),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_488),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_529),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_529),
.A2(n_419),
.B1(n_399),
.B2(n_403),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_515),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_488),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_481),
.B(n_207),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_529),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_485),
.Y(n_683)
);

INVxp33_ASAP7_75t_L g684 ( 
.A(n_522),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_436),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_535),
.B(n_318),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_500),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_535),
.B(n_317),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_500),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_521),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_500),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_500),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_485),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_502),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_615),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_635),
.A2(n_493),
.B1(n_535),
.B2(n_329),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_607),
.B(n_535),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_621),
.B(n_528),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_656),
.A2(n_489),
.B1(n_231),
.B2(n_334),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_630),
.B(n_469),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_612),
.B(n_535),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_556),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_656),
.A2(n_281),
.B1(n_312),
.B2(n_286),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_659),
.B(n_469),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_612),
.B(n_536),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_613),
.B(n_536),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_685),
.B(n_521),
.C(n_490),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_613),
.B(n_536),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_614),
.B(n_536),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_670),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_572),
.B(n_200),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_614),
.B(n_537),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_578),
.B(n_537),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_659),
.B(n_324),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_661),
.B(n_335),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_661),
.B(n_205),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_549),
.A2(n_478),
.B(n_540),
.C(n_403),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_636),
.B(n_397),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_648),
.B(n_561),
.Y(n_719)
);

AOI22x1_ASAP7_75t_L g720 ( 
.A1(n_663),
.A2(n_361),
.B1(n_365),
.B2(n_366),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_531),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_556),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_549),
.A2(n_493),
.B1(n_354),
.B2(n_351),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_556),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_561),
.B(n_208),
.Y(n_725)
);

BUFx12f_ASAP7_75t_SL g726 ( 
.A(n_649),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_555),
.A2(n_493),
.B1(n_537),
.B2(n_358),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_676),
.A2(n_540),
.B(n_493),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_676),
.B(n_208),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_555),
.B(n_493),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_648),
.B(n_284),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_618),
.B(n_513),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_619),
.B(n_513),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_619),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_437),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_629),
.Y(n_736)
);

AO221x1_ASAP7_75t_L g737 ( 
.A1(n_609),
.A2(n_441),
.B1(n_437),
.B2(n_438),
.C(n_439),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_682),
.A2(n_209),
.B1(n_355),
.B2(n_357),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_690),
.A2(n_646),
.B1(n_684),
.B2(n_622),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_552),
.B(n_496),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_629),
.B(n_513),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_550),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_631),
.B(n_632),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_631),
.B(n_632),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_553),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_606),
.B(n_209),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_650),
.B(n_513),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_617),
.B(n_305),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_606),
.B(n_211),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_650),
.B(n_513),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_575),
.B(n_438),
.Y(n_751)
);

INVx8_ASAP7_75t_L g752 ( 
.A(n_644),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_553),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_652),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_651),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_651),
.B(n_513),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_655),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_559),
.B(n_439),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_655),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_570),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_657),
.B(n_495),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_657),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_626),
.A2(n_347),
.B1(n_330),
.B2(n_323),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_574),
.B(n_626),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_605),
.B(n_441),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_606),
.B(n_212),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_570),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_606),
.B(n_212),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_662),
.B(n_667),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_662),
.B(n_667),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_681),
.B(n_634),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_636),
.B(n_670),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_670),
.A2(n_213),
.B1(n_222),
.B2(n_225),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_573),
.B(n_213),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_636),
.B(n_222),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_587),
.B(n_444),
.C(n_443),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_571),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_653),
.B(n_225),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_SL g779 ( 
.A(n_620),
.B(n_305),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_658),
.B(n_234),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_663),
.B(n_574),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_638),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_565),
.A2(n_357),
.B1(n_368),
.B2(n_364),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_665),
.B(n_502),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_665),
.B(n_502),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_671),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_623),
.B(n_443),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_640),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_673),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_571),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_678),
.Y(n_791)
);

O2A1O1Ixp5_ASAP7_75t_L g792 ( 
.A1(n_688),
.A2(n_498),
.B(n_507),
.C(n_512),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_665),
.B(n_502),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_664),
.B(n_444),
.Y(n_794)
);

AO221x1_ASAP7_75t_L g795 ( 
.A1(n_678),
.A2(n_445),
.B1(n_271),
.B2(n_398),
.C(n_413),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_665),
.B(n_502),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_234),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_627),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_565),
.B(n_445),
.Y(n_799)
);

BUFx5_ASAP7_75t_L g800 ( 
.A(n_694),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_679),
.B(n_498),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_565),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_679),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_586),
.B(n_319),
.C(n_236),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_610),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_547),
.B(n_236),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_668),
.B(n_319),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_686),
.B(n_496),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_547),
.B(n_325),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_669),
.A2(n_355),
.B1(n_349),
.B2(n_348),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_565),
.A2(n_507),
.B(n_512),
.C(n_542),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_551),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_649),
.B(n_398),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_558),
.B(n_507),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_558),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_562),
.B(n_512),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_677),
.A2(n_404),
.B(n_399),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_639),
.B(n_325),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_563),
.B(n_568),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_563),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_568),
.B(n_246),
.C(n_242),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_576),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_687),
.B(n_502),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_584),
.A2(n_327),
.B1(n_332),
.B2(n_342),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_579),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_583),
.B(n_485),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_583),
.B(n_327),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_588),
.B(n_332),
.Y(n_828)
);

NOR2x1p5_ASAP7_75t_L g829 ( 
.A(n_588),
.B(n_218),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_589),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_589),
.B(n_518),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_557),
.B(n_404),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_687),
.B(n_518),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_689),
.B(n_342),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_689),
.B(n_518),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_691),
.B(n_539),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_691),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_692),
.B(n_253),
.C(n_250),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_692),
.B(n_343),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_584),
.B(n_268),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_580),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_593),
.A2(n_544),
.B(n_543),
.C(n_542),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_584),
.B(n_405),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_554),
.B(n_343),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_557),
.A2(n_330),
.B1(n_223),
.B2(n_227),
.Y(n_845)
);

BUFx5_ASAP7_75t_L g846 ( 
.A(n_694),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_594),
.B(n_599),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_594),
.B(n_599),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_584),
.B(n_405),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_610),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_610),
.B(n_344),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_580),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_719),
.A2(n_584),
.B1(n_628),
.B2(n_554),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_802),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_802),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_730),
.A2(n_728),
.B(n_792),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_697),
.B(n_627),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_781),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_764),
.B(n_407),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_781),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_695),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_710),
.B(n_560),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_710),
.B(n_560),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_710),
.B(n_577),
.Y(n_864)
);

NOR2x2_ASAP7_75t_L g865 ( 
.A(n_700),
.B(n_604),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_710),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_805),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_736),
.B(n_577),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_698),
.B1(n_754),
.B2(n_704),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_765),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_734),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_850),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_R g874 ( 
.A(n_788),
.B(n_666),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_752),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_794),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_755),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_723),
.B(n_546),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_784),
.A2(n_624),
.B(n_545),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_R g880 ( 
.A(n_726),
.B(n_666),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_721),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_704),
.A2(n_731),
.B1(n_771),
.B2(n_843),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_735),
.B(n_731),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_713),
.B(n_546),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_702),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_752),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_757),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_830),
.B(n_672),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_752),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_739),
.B(n_247),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_718),
.B(n_683),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_774),
.A2(n_591),
.B(n_557),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_759),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

NOR3x1_ASAP7_75t_L g895 ( 
.A(n_795),
.B(n_409),
.C(n_407),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_724),
.Y(n_896)
);

AND2x2_ASAP7_75t_SL g897 ( 
.A(n_845),
.B(n_611),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_700),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_762),
.B(n_672),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_786),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_700),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_771),
.A2(n_591),
.B1(n_641),
.B2(n_616),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_789),
.Y(n_903)
);

AND2x4_ASAP7_75t_SL g904 ( 
.A(n_799),
.B(n_305),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_791),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_774),
.B(n_262),
.C(n_256),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_803),
.B(n_812),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_723),
.A2(n_591),
.B1(n_680),
.B2(n_674),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_703),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_739),
.B(n_264),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_815),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_820),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_800),
.B(n_546),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_742),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_717),
.A2(n_604),
.B(n_645),
.C(n_647),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_699),
.Y(n_916)
);

AO22x1_ASAP7_75t_L g917 ( 
.A1(n_797),
.A2(n_331),
.B1(n_220),
.B2(n_230),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_849),
.A2(n_616),
.B1(n_633),
.B2(n_641),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_718),
.Y(n_919)
);

AND2x2_ASAP7_75t_SL g920 ( 
.A(n_845),
.B(n_696),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_751),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_707),
.B(n_409),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_822),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_837),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_745),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_758),
.B(n_740),
.Y(n_926)
);

AND3x1_ASAP7_75t_L g927 ( 
.A(n_804),
.B(n_412),
.C(n_410),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_753),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_799),
.B(n_829),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_837),
.B(n_674),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_798),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_799),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_760),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_847),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_840),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_743),
.B(n_680),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_548),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_763),
.B(n_412),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_782),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_792),
.A2(n_645),
.B(n_633),
.Y(n_940)
);

AND2x6_ASAP7_75t_L g941 ( 
.A(n_798),
.B(n_611),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_769),
.B(n_548),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_798),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_767),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_777),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_770),
.B(n_548),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_848),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_790),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_763),
.B(n_413),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_800),
.B(n_546),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_800),
.B(n_546),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_819),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_806),
.B(n_548),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_727),
.A2(n_581),
.B1(n_582),
.B2(n_597),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_727),
.A2(n_701),
.B(n_811),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_748),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_825),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_841),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_772),
.B(n_683),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_838),
.B(n_683),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_784),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_761),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_787),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_737),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_696),
.A2(n_832),
.B1(n_720),
.B2(n_725),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_806),
.B(n_809),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_808),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_778),
.A2(n_647),
.B1(n_611),
.B2(n_693),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_852),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_775),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_800),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_809),
.B(n_566),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_817),
.A2(n_581),
.B1(n_582),
.B2(n_597),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_801),
.A2(n_362),
.B1(n_371),
.B2(n_370),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_800),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_800),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_785),
.A2(n_545),
.B(n_675),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_714),
.B(n_715),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_714),
.B(n_566),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_846),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_814),
.A2(n_360),
.B1(n_371),
.B2(n_363),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_785),
.B(n_546),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_787),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_821),
.B(n_693),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_715),
.B(n_566),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_846),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_846),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_779),
.B(n_344),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_787),
.Y(n_989)
);

OR2x2_ASAP7_75t_SL g990 ( 
.A(n_797),
.B(n_804),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_746),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_846),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_711),
.A2(n_693),
.B1(n_566),
.B2(n_625),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_816),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_846),
.B(n_567),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_776),
.B(n_567),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_846),
.B(n_567),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_833),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_749),
.B(n_416),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_783),
.B(n_738),
.C(n_766),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_768),
.B(n_273),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_835),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_L g1003 ( 
.A(n_836),
.B(n_567),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_851),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_705),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_706),
.A2(n_275),
.B1(n_323),
.B2(n_331),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_776),
.B(n_590),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_708),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_709),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_793),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_827),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_793),
.A2(n_675),
.B(n_660),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_773),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_716),
.A2(n_729),
.B1(n_807),
.B2(n_780),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_834),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_712),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_732),
.B(n_585),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_595),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_810),
.B(n_416),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_826),
.B(n_595),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_828),
.Y(n_1021)
);

NOR3x1_ASAP7_75t_L g1022 ( 
.A(n_824),
.B(n_417),
.C(n_430),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_733),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_823),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_796),
.A2(n_369),
.B1(n_364),
.B2(n_368),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_741),
.B(n_747),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_750),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_886),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_953),
.A2(n_796),
.B(n_756),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_966),
.B(n_818),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_941),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_SL g1034 ( 
.A(n_989),
.B(n_585),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_890),
.A2(n_844),
.B(n_842),
.C(n_417),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_972),
.A2(n_603),
.B(n_600),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_883),
.B(n_926),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_952),
.B(n_595),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_920),
.A2(n_882),
.B1(n_965),
.B2(n_869),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_919),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_878),
.A2(n_675),
.B(n_660),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_920),
.A2(n_348),
.B1(n_349),
.B2(n_369),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_934),
.B(n_625),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_919),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_947),
.B(n_625),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_873),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_866),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_878),
.A2(n_675),
.B(n_660),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_940),
.A2(n_637),
.B(n_625),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_SL g1050 ( 
.A1(n_892),
.A2(n_430),
.B(n_428),
.C(n_421),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_886),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_857),
.A2(n_660),
.B(n_624),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_876),
.B(n_585),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_924),
.B(n_637),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_989),
.B(n_585),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_860),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_864),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_962),
.B(n_637),
.Y(n_1058)
);

INVx3_ASAP7_75t_SL g1059 ( 
.A(n_898),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_965),
.A2(n_637),
.B1(n_642),
.B2(n_643),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1010),
.A2(n_643),
.B1(n_642),
.B2(n_564),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_856),
.A2(n_600),
.B(n_601),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_921),
.B(n_277),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_873),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_SL g1065 ( 
.A(n_916),
.B(n_275),
.C(n_362),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_860),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_864),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_870),
.B(n_916),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_SL g1069 ( 
.A1(n_908),
.A2(n_419),
.B(n_420),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_R g1070 ( 
.A(n_880),
.B(n_339),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_890),
.A2(n_420),
.B(n_428),
.C(n_421),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_866),
.B(n_545),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_866),
.B(n_624),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_875),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_989),
.B(n_909),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_879),
.A2(n_603),
.B(n_602),
.Y(n_1076)
);

AO32x1_ASAP7_75t_L g1077 ( 
.A1(n_964),
.A2(n_602),
.A3(n_497),
.B1(n_542),
.B2(n_543),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_980),
.B(n_564),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_910),
.A2(n_497),
.B(n_543),
.C(n_539),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_864),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_915),
.A2(n_544),
.B(n_121),
.C(n_188),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_SL g1082 ( 
.A1(n_1027),
.A2(n_302),
.B(n_304),
.C(n_310),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_861),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_859),
.B(n_315),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_961),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_931),
.B(n_564),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_871),
.B(n_347),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1010),
.A2(n_643),
.B1(n_642),
.B2(n_598),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_L g1089 ( 
.A(n_941),
.B(n_971),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_939),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_994),
.B(n_544),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_872),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_995),
.A2(n_643),
.B(n_642),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_941),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_997),
.A2(n_868),
.B(n_977),
.Y(n_1095)
);

AOI22x1_ASAP7_75t_L g1096 ( 
.A1(n_1028),
.A2(n_643),
.B1(n_642),
.B2(n_598),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1000),
.A2(n_514),
.B1(n_359),
.B2(n_592),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_932),
.B(n_80),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_998),
.B(n_1002),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1012),
.A2(n_598),
.B(n_596),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_1013),
.B(n_598),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_998),
.B(n_596),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_937),
.A2(n_598),
.B(n_596),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_922),
.B(n_7),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_858),
.B(n_78),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_942),
.A2(n_596),
.B(n_592),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1002),
.B(n_596),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_867),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_SL g1109 ( 
.A1(n_915),
.A2(n_85),
.B(n_184),
.C(n_179),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_935),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_946),
.A2(n_596),
.B(n_592),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_877),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_991),
.A2(n_592),
.B1(n_569),
.B2(n_564),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_907),
.B(n_887),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_901),
.B(n_585),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_885),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_910),
.A2(n_1001),
.B(n_1021),
.C(n_956),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_889),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1010),
.A2(n_592),
.B1(n_569),
.B2(n_564),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1026),
.A2(n_9),
.B(n_10),
.C(n_13),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_854),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_893),
.B(n_564),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_989),
.B(n_585),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_929),
.B(n_569),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_991),
.B(n_569),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1014),
.A2(n_569),
.B1(n_65),
.B2(n_74),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_978),
.A2(n_955),
.B(n_906),
.C(n_1011),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1003),
.A2(n_569),
.B(n_62),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_885),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_938),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_961),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_999),
.B(n_14),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_970),
.A2(n_16),
.B(n_17),
.C(n_24),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_961),
.A2(n_97),
.B1(n_168),
.B2(n_154),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_900),
.B(n_903),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_901),
.B(n_1015),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_865),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_855),
.B(n_153),
.Y(n_1138)
);

AO32x2_ASAP7_75t_L g1139 ( 
.A1(n_897),
.A2(n_25),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_971),
.A2(n_514),
.B(n_89),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_963),
.Y(n_1141)
);

AOI222xp33_ASAP7_75t_L g1142 ( 
.A1(n_949),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.C1(n_32),
.C2(n_33),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_905),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1019),
.B(n_34),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_911),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1027),
.A2(n_127),
.B(n_151),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_975),
.A2(n_514),
.B(n_124),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_975),
.A2(n_514),
.B(n_132),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_912),
.B(n_39),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_976),
.A2(n_514),
.B(n_133),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_881),
.Y(n_1151)
);

AO32x1_ASAP7_75t_L g1152 ( 
.A1(n_923),
.A2(n_1009),
.A3(n_1016),
.B1(n_1008),
.B2(n_928),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_941),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_881),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_983),
.B(n_40),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1004),
.A2(n_40),
.B(n_42),
.C(n_45),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_881),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1023),
.B(n_48),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_943),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_898),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_897),
.A2(n_984),
.B1(n_891),
.B2(n_996),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_961),
.A2(n_139),
.B1(n_149),
.B2(n_147),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_930),
.B(n_48),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_941),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_891),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_929),
.B(n_136),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_899),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_929),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_983),
.B(n_49),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_874),
.B(n_115),
.Y(n_1170)
);

NAND2xp33_ASAP7_75t_L g1171 ( 
.A(n_874),
.B(n_514),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_996),
.A2(n_1007),
.B1(n_927),
.B2(n_891),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_917),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_986),
.A2(n_120),
.B1(n_141),
.B2(n_142),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_987),
.A2(n_992),
.B(n_936),
.Y(n_1175)
);

AO32x2_ASAP7_75t_L g1176 ( 
.A1(n_1039),
.A2(n_865),
.A3(n_895),
.B1(n_1022),
.B2(n_908),
.Y(n_1176)
);

NOR4xp25_ASAP7_75t_L g1177 ( 
.A(n_1120),
.B(n_974),
.C(n_981),
.D(n_1006),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1095),
.A2(n_884),
.B(n_1020),
.Y(n_1178)
);

CKINVDCx8_ASAP7_75t_R g1179 ( 
.A(n_1029),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_1170),
.A2(n_884),
.B(n_984),
.C(n_960),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1114),
.B(n_1006),
.Y(n_1181)
);

AOI31xp67_ASAP7_75t_L g1182 ( 
.A1(n_1172),
.A2(n_902),
.A3(n_853),
.B(n_968),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1037),
.B(n_981),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1032),
.B(n_974),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1110),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1094),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1068),
.B(n_904),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1151),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1167),
.B(n_1005),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1137),
.B(n_904),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1117),
.B(n_1143),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1127),
.A2(n_954),
.B(n_960),
.Y(n_1192)
);

AO21x2_ASAP7_75t_L g1193 ( 
.A1(n_1036),
.A2(n_918),
.B(n_1017),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1033),
.B(n_943),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1083),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1056),
.B(n_1066),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1051),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1118),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1142),
.B(n_988),
.C(n_880),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_SL g1200 ( 
.A1(n_1126),
.A2(n_944),
.B(n_957),
.C(n_969),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1142),
.A2(n_1007),
.B(n_996),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1035),
.A2(n_1007),
.B(n_984),
.C(n_1018),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_950),
.B(n_913),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1049),
.A2(n_862),
.B(n_863),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1099),
.B(n_888),
.Y(n_1205)
);

BUFx4_ASAP7_75t_SL g1206 ( 
.A(n_1154),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1144),
.B(n_1025),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1092),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1074),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1094),
.B(n_1025),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_SL g1211 ( 
.A1(n_1130),
.A2(n_1017),
.B(n_985),
.C(n_979),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1132),
.B(n_1024),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1090),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1160),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1112),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1059),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1030),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1121),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1031),
.A2(n_960),
.B(n_951),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1137),
.B(n_948),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1050),
.A2(n_954),
.B(n_993),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1175),
.A2(n_951),
.B(n_950),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1052),
.A2(n_913),
.B(n_959),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1135),
.B(n_1024),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1040),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1040),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1056),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1046),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1125),
.B(n_1104),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1101),
.B(n_959),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1093),
.A2(n_973),
.B(n_896),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1128),
.A2(n_973),
.B(n_925),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1113),
.A2(n_959),
.B(n_982),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1163),
.B(n_933),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1082),
.A2(n_896),
.B(n_894),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1063),
.B(n_914),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1056),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1168),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1158),
.B(n_933),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1064),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1173),
.B(n_944),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1172),
.A2(n_969),
.B(n_957),
.C(n_928),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1153),
.B(n_894),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1141),
.B(n_958),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1153),
.Y(n_1245)
);

CKINVDCx11_ASAP7_75t_R g1246 ( 
.A(n_1157),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1149),
.B(n_945),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1116),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1103),
.A2(n_1106),
.B(n_1111),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_SL g1250 ( 
.A(n_1164),
.B(n_49),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1057),
.B(n_55),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1096),
.A2(n_514),
.B(n_1089),
.Y(n_1252)
);

BUFx10_ASAP7_75t_L g1253 ( 
.A(n_1087),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1129),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1061),
.A2(n_1119),
.B(n_1088),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1161),
.A2(n_1091),
.B(n_1060),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1075),
.B(n_1136),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1042),
.B(n_1071),
.C(n_1156),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1065),
.B(n_1155),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1062),
.A2(n_1102),
.B(n_1107),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1108),
.Y(n_1261)
);

AND2x6_ASAP7_75t_L g1262 ( 
.A(n_1085),
.B(n_1131),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1069),
.B(n_1058),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1145),
.A2(n_1164),
.B(n_1174),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1152),
.A2(n_1077),
.A3(n_1122),
.B(n_1038),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1057),
.B(n_1067),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1146),
.A2(n_1078),
.B(n_1062),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1152),
.A2(n_1077),
.A3(n_1043),
.B(n_1045),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1124),
.A2(n_1105),
.B1(n_1097),
.B2(n_1131),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1078),
.A2(n_1073),
.B(n_1072),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1081),
.A2(n_1109),
.B(n_1054),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1152),
.A2(n_1077),
.A3(n_1134),
.B(n_1162),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1072),
.A2(n_1073),
.B(n_1086),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1140),
.A2(n_1150),
.B(n_1148),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1040),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1147),
.A2(n_1047),
.A3(n_1169),
.B(n_1165),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1080),
.B(n_1066),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1171),
.A2(n_1138),
.B(n_1053),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1115),
.A2(n_1123),
.B(n_1055),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1159),
.A2(n_1166),
.B(n_1047),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1168),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1070),
.Y(n_1282)
);

NOR4xp25_ASAP7_75t_L g1283 ( 
.A(n_1139),
.B(n_1085),
.C(n_1131),
.D(n_1098),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1098),
.B(n_1044),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1124),
.B(n_1034),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1124),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1139),
.A2(n_1039),
.B(n_1127),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1139),
.B(n_607),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1041),
.A2(n_878),
.B(n_1048),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1114),
.B(n_607),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1114),
.B(n_607),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1039),
.A2(n_1127),
.B(n_966),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1084),
.B(n_883),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1094),
.A2(n_1164),
.B(n_1153),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1117),
.B(n_698),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1114),
.B(n_607),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1110),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1130),
.A2(n_845),
.B1(n_1039),
.B2(n_966),
.C(n_1120),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1041),
.A2(n_878),
.B(n_1048),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1114),
.B(n_607),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1030),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1083),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1127),
.A2(n_966),
.B(n_1170),
.C(n_1130),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1083),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1114),
.B(n_607),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1039),
.A2(n_1060),
.A3(n_1095),
.B(n_1127),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1114),
.A2(n_966),
.B1(n_920),
.B2(n_882),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1076),
.A2(n_1049),
.B(n_1100),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1114),
.A2(n_966),
.B1(n_920),
.B2(n_882),
.Y(n_1309)
);

AOI221xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1130),
.A2(n_845),
.B1(n_1039),
.B2(n_966),
.C(n_1120),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1032),
.A2(n_966),
.B(n_698),
.C(n_607),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1083),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1117),
.B(n_698),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_SL g1314 ( 
.A(n_1033),
.B(n_1094),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1127),
.A2(n_966),
.B(n_1170),
.C(n_1130),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1191),
.B(n_1184),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1311),
.A2(n_1258),
.B(n_1295),
.C(n_1313),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1229),
.B(n_1220),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1245),
.B(n_1186),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1264),
.A2(n_1250),
.B(n_1278),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1217),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1185),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1293),
.B(n_1244),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1195),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1267),
.A2(n_1223),
.B(n_1204),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1218),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1290),
.A2(n_1296),
.B(n_1291),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1194),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1245),
.B(n_1186),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1300),
.A2(n_1305),
.B1(n_1257),
.B2(n_1181),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1178),
.A2(n_1231),
.B(n_1222),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1287),
.A2(n_1192),
.B(n_1201),
.C(n_1307),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1287),
.A2(n_1255),
.B(n_1221),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1199),
.A2(n_1309),
.B1(n_1183),
.B2(n_1259),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1275),
.Y(n_1335)
);

AOI222xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1185),
.A2(n_1297),
.B1(n_1213),
.B2(n_1208),
.C1(n_1215),
.C2(n_1312),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1240),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1236),
.B(n_1297),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1245),
.B(n_1286),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1302),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1207),
.B(n_1225),
.Y(n_1341)
);

INVx3_ASAP7_75t_SL g1342 ( 
.A(n_1197),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1248),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1304),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1226),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1209),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1177),
.A2(n_1180),
.B(n_1315),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1189),
.B(n_1212),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1219),
.A2(n_1260),
.B(n_1252),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1303),
.A2(n_1298),
.B(n_1310),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1187),
.A2(n_1269),
.B1(n_1284),
.B2(n_1241),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1192),
.A2(n_1201),
.B(n_1298),
.C(n_1233),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1228),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1254),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_SL g1355 ( 
.A(n_1196),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1206),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1274),
.A2(n_1270),
.B(n_1235),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1196),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1274),
.A2(n_1235),
.B(n_1273),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1200),
.A2(n_1263),
.B(n_1221),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1261),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1294),
.B(n_1269),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1263),
.A2(n_1242),
.B(n_1202),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1198),
.B(n_1239),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1253),
.A2(n_1234),
.B1(n_1247),
.B2(n_1256),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1227),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1282),
.B(n_1230),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1214),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1245),
.B(n_1277),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1203),
.A2(n_1224),
.B(n_1279),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1251),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1256),
.A2(n_1205),
.B1(n_1190),
.B2(n_1246),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1211),
.A2(n_1182),
.B(n_1280),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1262),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1210),
.A2(n_1285),
.B1(n_1188),
.B2(n_1314),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1243),
.B(n_1266),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1306),
.A2(n_1272),
.A3(n_1271),
.B(n_1265),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1286),
.A2(n_1281),
.B1(n_1238),
.B2(n_1216),
.Y(n_1378)
);

INVx8_ASAP7_75t_L g1379 ( 
.A(n_1262),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1262),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1227),
.B(n_1237),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1193),
.A2(n_1306),
.B(n_1268),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1237),
.A2(n_1176),
.B1(n_1301),
.B2(n_1283),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1176),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1283),
.A2(n_1272),
.B1(n_1276),
.B2(n_1179),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1276),
.A2(n_1265),
.B(n_1272),
.Y(n_1386)
);

AOI21xp33_ASAP7_75t_L g1387 ( 
.A1(n_1191),
.A2(n_966),
.B(n_1184),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1287),
.A2(n_1249),
.B(n_1292),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_SL g1389 ( 
.A(n_1179),
.B(n_1151),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1199),
.A2(n_920),
.B1(n_1142),
.B2(n_1184),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1245),
.B(n_1033),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1218),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1218),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1287),
.A2(n_1249),
.B(n_1292),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1229),
.B(n_1220),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1287),
.A2(n_1249),
.B(n_1292),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1195),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1199),
.A2(n_920),
.B1(n_1142),
.B2(n_1184),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1308),
.A2(n_1299),
.B(n_1289),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1184),
.A2(n_966),
.B1(n_1199),
.B2(n_1201),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1216),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1184),
.A2(n_966),
.B1(n_1199),
.B2(n_1201),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1184),
.A2(n_966),
.B1(n_1199),
.B2(n_1201),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1191),
.A2(n_966),
.B1(n_1291),
.B2(n_1290),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1264),
.A2(n_1250),
.B(n_1278),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1191),
.A2(n_748),
.B1(n_779),
.B2(n_920),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1255),
.A2(n_1039),
.A3(n_1249),
.B(n_1288),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1191),
.B(n_1184),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1287),
.A2(n_1249),
.B(n_1292),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1255),
.A2(n_1039),
.A3(n_1249),
.B(n_1288),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1195),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1191),
.A2(n_966),
.B1(n_1291),
.B2(n_1290),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1293),
.B(n_1244),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_SL g1414 ( 
.A1(n_1264),
.A2(n_1250),
.B(n_1278),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1196),
.B(n_1245),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1195),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_SL g1417 ( 
.A(n_1191),
.B(n_779),
.C(n_748),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1264),
.A2(n_1250),
.B(n_1278),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1191),
.B(n_1184),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1191),
.A2(n_966),
.B1(n_1291),
.B2(n_1290),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1191),
.A2(n_748),
.B1(n_779),
.B2(n_920),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1191),
.B(n_1184),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1308),
.A2(n_1299),
.B(n_1289),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1195),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1293),
.B(n_1244),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1195),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1195),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1196),
.B(n_1245),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1308),
.A2(n_1299),
.B(n_1289),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1195),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1293),
.B(n_1244),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1293),
.B(n_1244),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1195),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1377),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1404),
.B(n_1412),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_1390),
.B2(n_1398),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1390),
.A2(n_1398),
.B1(n_1422),
.B2(n_1408),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1362),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1316),
.B(n_1408),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1337),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1343),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1316),
.A2(n_1419),
.B1(n_1422),
.B2(n_1334),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1391),
.A2(n_1417),
.B(n_1330),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1419),
.A2(n_1334),
.B1(n_1367),
.B2(n_1378),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1323),
.B(n_1413),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1335),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1347),
.A2(n_1360),
.B(n_1373),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1425),
.B(n_1431),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1432),
.B(n_1341),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1387),
.A2(n_1420),
.B(n_1317),
.C(n_1402),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1338),
.B(n_1367),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1392),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1400),
.A2(n_1403),
.B(n_1402),
.C(n_1351),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1364),
.B(n_1318),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1322),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1378),
.A2(n_1332),
.B1(n_1372),
.B2(n_1352),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1415),
.B(n_1428),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1332),
.A2(n_1372),
.B1(n_1352),
.B2(n_1375),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1392),
.B(n_1393),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1400),
.A2(n_1403),
.B(n_1327),
.C(n_1371),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1393),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1350),
.A2(n_1360),
.B(n_1383),
.C(n_1365),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1348),
.B(n_1326),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1335),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1340),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1344),
.B(n_1397),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1366),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1366),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1365),
.A2(n_1418),
.B1(n_1405),
.B2(n_1414),
.C(n_1320),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1411),
.A2(n_1433),
.B(n_1426),
.C(n_1416),
.Y(n_1470)
);

NOR2xp67_ASAP7_75t_L g1471 ( 
.A(n_1353),
.B(n_1354),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1383),
.A2(n_1385),
.B(n_1379),
.C(n_1384),
.Y(n_1472)
);

AOI21x1_ASAP7_75t_SL g1473 ( 
.A1(n_1369),
.A2(n_1336),
.B(n_1333),
.Y(n_1473)
);

OAI31xp33_ASAP7_75t_L g1474 ( 
.A1(n_1368),
.A2(n_1346),
.A3(n_1321),
.B(n_1345),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_SL g1475 ( 
.A(n_1362),
.B(n_1374),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1362),
.A2(n_1385),
.B1(n_1430),
.B2(n_1427),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1342),
.Y(n_1477)
);

AOI21x1_ASAP7_75t_SL g1478 ( 
.A1(n_1333),
.A2(n_1388),
.B(n_1394),
.Y(n_1478)
);

AOI211xp5_ASAP7_75t_L g1479 ( 
.A1(n_1342),
.A2(n_1389),
.B(n_1424),
.C(n_1321),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1361),
.B(n_1328),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1401),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1374),
.A2(n_1355),
.B1(n_1339),
.B2(n_1380),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1381),
.B(n_1339),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1379),
.A2(n_1363),
.B(n_1359),
.C(n_1357),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1388),
.B(n_1394),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1396),
.B(n_1409),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1355),
.A2(n_1363),
.B1(n_1391),
.B2(n_1319),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1396),
.B(n_1409),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1359),
.A2(n_1382),
.B(n_1399),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1319),
.A2(n_1329),
.B1(n_1401),
.B2(n_1356),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1370),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1386),
.B(n_1377),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1377),
.B(n_1376),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1376),
.Y(n_1498)
);

O2A1O1Ixp5_ASAP7_75t_L g1499 ( 
.A1(n_1331),
.A2(n_1349),
.B(n_1325),
.C(n_1429),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1423),
.B(n_1358),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1318),
.B(n_1395),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1323),
.B(n_1413),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1323),
.B(n_1413),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1401),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1323),
.B(n_1413),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1417),
.A2(n_1311),
.B(n_966),
.C(n_1258),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1404),
.B(n_1412),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1324),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1347),
.A2(n_1360),
.B(n_1373),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_916),
.B2(n_1191),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_916),
.B2(n_1191),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_916),
.B2(n_1191),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1316),
.B(n_1408),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_916),
.B2(n_1191),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1335),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1417),
.A2(n_1311),
.B(n_966),
.C(n_1258),
.Y(n_1516)
);

BUFx12f_ASAP7_75t_L g1517 ( 
.A(n_1401),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1401),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1347),
.A2(n_1360),
.B(n_1373),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1417),
.A2(n_1311),
.B(n_966),
.C(n_1258),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1323),
.B(n_1413),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1417),
.A2(n_1311),
.B(n_966),
.C(n_1258),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1406),
.A2(n_1421),
.B1(n_916),
.B2(n_1191),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1404),
.B(n_1412),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_R g1525 ( 
.A(n_1517),
.B(n_1477),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1500),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1500),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1435),
.B(n_1507),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1441),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1495),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_SL g1531 ( 
.A(n_1464),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1524),
.B(n_1439),
.Y(n_1532)
);

INVxp33_ASAP7_75t_L g1533 ( 
.A(n_1451),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1453),
.B(n_1487),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1446),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1482),
.B(n_1485),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1439),
.B(n_1513),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1442),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1488),
.B(n_1492),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1489),
.B(n_1486),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1461),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1498),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1443),
.B(n_1491),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1447),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1452),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1434),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1459),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1490),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_SL g1550 ( 
.A(n_1438),
.B(n_1458),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1515),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1447),
.B(n_1509),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1497),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1447),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1509),
.B(n_1519),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1465),
.B(n_1452),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1470),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1499),
.A2(n_1462),
.B(n_1496),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1501),
.B(n_1454),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1450),
.B(n_1437),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1466),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1506),
.A2(n_1522),
.B(n_1520),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1460),
.B(n_1471),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1476),
.B(n_1456),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1484),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1472),
.A2(n_1436),
.B(n_1516),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1449),
.B(n_1505),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1444),
.A2(n_1523),
.B1(n_1514),
.B2(n_1512),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1493),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1479),
.B(n_1474),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1549),
.B(n_1463),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1493),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1571),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1571),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1545),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1545),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1529),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1478),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1553),
.B(n_1455),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1529),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1536),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1537),
.B(n_1440),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1556),
.B(n_1469),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1547),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1554),
.Y(n_1587)
);

AOI222xp33_ASAP7_75t_L g1588 ( 
.A1(n_1561),
.A2(n_1511),
.B1(n_1510),
.B2(n_1448),
.C1(n_1503),
.C2(n_1521),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1543),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1527),
.B(n_1475),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1445),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1547),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1541),
.B(n_1548),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1559),
.B(n_1502),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1570),
.A2(n_1473),
.B(n_1494),
.C(n_1483),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1586),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1588),
.A2(n_1570),
.B1(n_1539),
.B2(n_1561),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1596),
.A2(n_1568),
.B1(n_1550),
.B2(n_1539),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1592),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1596),
.A2(n_1572),
.B1(n_1564),
.B2(n_1585),
.C(n_1528),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1592),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1594),
.B(n_1530),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1581),
.A2(n_1566),
.B1(n_1534),
.B2(n_1528),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1594),
.B(n_1530),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1588),
.A2(n_1568),
.B1(n_1566),
.B2(n_1564),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1575),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1593),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1575),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1581),
.Y(n_1615)
);

NOR4xp25_ASAP7_75t_SL g1616 ( 
.A(n_1589),
.B(n_1558),
.C(n_1550),
.D(n_1567),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1581),
.A2(n_1566),
.B1(n_1534),
.B2(n_1532),
.Y(n_1618)
);

BUFx10_ASAP7_75t_L g1619 ( 
.A(n_1595),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_R g1620 ( 
.A(n_1573),
.B(n_1481),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1579),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1624)
);

OAI33xp33_ASAP7_75t_L g1625 ( 
.A1(n_1593),
.A2(n_1532),
.A3(n_1557),
.B1(n_1538),
.B2(n_1558),
.B3(n_1565),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1585),
.A2(n_1565),
.B1(n_1568),
.B2(n_1533),
.C(n_1560),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1585),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1580),
.B(n_1566),
.C(n_1534),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1582),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1566),
.C(n_1534),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1590),
.A2(n_1568),
.B1(n_1534),
.B2(n_1544),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1544),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1574),
.B(n_1526),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1595),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1590),
.A2(n_1544),
.B1(n_1531),
.B2(n_1457),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1578),
.A2(n_1542),
.B1(n_1562),
.B2(n_1546),
.C(n_1557),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1582),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1583),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1574),
.B(n_1526),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1584),
.B(n_1525),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1584),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1569),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1634),
.B(n_1587),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1598),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

CKINVDCx14_ASAP7_75t_R g1646 ( 
.A(n_1620),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1598),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1613),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1617),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1612),
.B(n_1578),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1623),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1610),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1623),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1629),
.Y(n_1656)
);

NOR2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1628),
.B(n_1535),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1606),
.B(n_1574),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1629),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1637),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1599),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1604),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1599),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1601),
.B(n_1603),
.Y(n_1665)
);

INVx4_ASAP7_75t_SL g1666 ( 
.A(n_1611),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1632),
.A2(n_1563),
.B(n_1555),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1601),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1603),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1622),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1605),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1649),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1642),
.B(n_1626),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1666),
.B(n_1650),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1660),
.B(n_1627),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1624),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1649),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1627),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1663),
.B(n_1636),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1666),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1666),
.B(n_1606),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1666),
.B(n_1650),
.Y(n_1688)
);

NOR2xp67_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1630),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1608),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1665),
.Y(n_1691)
);

NAND2x1_ASAP7_75t_L g1692 ( 
.A(n_1643),
.B(n_1611),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1608),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1653),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1669),
.B(n_1602),
.C(n_1618),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1650),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1650),
.B(n_1633),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1652),
.B(n_1633),
.Y(n_1699)
);

BUFx2_ASAP7_75t_SL g1700 ( 
.A(n_1652),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1652),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1652),
.B(n_1639),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1655),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.B(n_1639),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1659),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1651),
.B(n_1641),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1659),
.Y(n_1708)
);

AND3x2_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1640),
.C(n_1638),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1665),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_SL g1711 ( 
.A(n_1651),
.B(n_1616),
.C(n_1631),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1662),
.B(n_1607),
.C(n_1635),
.D(n_1615),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

OAI31xp33_ASAP7_75t_L g1714 ( 
.A1(n_1657),
.A2(n_1615),
.A3(n_1597),
.B(n_1580),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1646),
.B(n_1504),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1658),
.B(n_1619),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_SL g1718 ( 
.A(n_1700),
.B(n_1535),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1706),
.Y(n_1719)
);

NAND4xp25_ASAP7_75t_L g1720 ( 
.A(n_1684),
.B(n_1662),
.C(n_1673),
.D(n_1664),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1713),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1687),
.B(n_1658),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.B(n_1643),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1706),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1678),
.B(n_1664),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1676),
.B(n_1646),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1708),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1709),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1708),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1674),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1716),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1693),
.B(n_1643),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1713),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1674),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1689),
.B(n_1668),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1679),
.B(n_1673),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1680),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1713),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1678),
.B(n_1683),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1680),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1686),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1683),
.B(n_1668),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1686),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1689),
.B(n_1569),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1694),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1677),
.B(n_1667),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1712),
.B(n_1504),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_1668),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1675),
.B(n_1643),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1677),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1737),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1739),
.B(n_1715),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1731),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1730),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1731),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1719),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1754),
.B(n_1685),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1754),
.B(n_1688),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1742),
.B(n_1691),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1721),
.Y(n_1764)
);

AOI21xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1727),
.A2(n_1695),
.B(n_1714),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1733),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1721),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1743),
.B(n_1710),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1703),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1722),
.B(n_1675),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1725),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1753),
.B(n_1682),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1753),
.B(n_1682),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1750),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1735),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1740),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1723),
.B(n_1685),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1741),
.B(n_1697),
.Y(n_1780)
);

OAI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1758),
.A2(n_1720),
.B(n_1738),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_R g1782 ( 
.A1(n_1765),
.A2(n_1752),
.B(n_1741),
.C(n_1726),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1766),
.B(n_1728),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1758),
.A2(n_1751),
.B1(n_1700),
.B2(n_1746),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1761),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1766),
.B(n_1752),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1762),
.B(n_1778),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1762),
.B(n_1740),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1755),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1765),
.B(n_1728),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1755),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1780),
.A2(n_1711),
.B1(n_1692),
.B2(n_1750),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1767),
.A2(n_1724),
.B(n_1723),
.Y(n_1793)
);

OAI32xp33_ASAP7_75t_L g1794 ( 
.A1(n_1780),
.A2(n_1749),
.A3(n_1778),
.B1(n_1756),
.B2(n_1763),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1769),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1767),
.B(n_1724),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1763),
.A2(n_1770),
.B1(n_1768),
.B2(n_1764),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1770),
.A2(n_1748),
.B(n_1747),
.C(n_1732),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_L g1799 ( 
.A(n_1774),
.B(n_1701),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1769),
.B(n_1525),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1785),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1786),
.B(n_1777),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1789),
.B(n_1768),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1797),
.B(n_1761),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1787),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1790),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1783),
.B(n_1774),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1788),
.B(n_1776),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1791),
.B(n_1776),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1797),
.B(n_1795),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1799),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1782),
.B1(n_1794),
.B2(n_1792),
.C(n_1781),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1807),
.B(n_1784),
.C(n_1800),
.D(n_1798),
.Y(n_1814)
);

OAI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1804),
.A2(n_1793),
.B1(n_1692),
.B2(n_1749),
.Y(n_1815)
);

NOR3xp33_ASAP7_75t_SL g1816 ( 
.A(n_1802),
.B(n_1771),
.C(n_1760),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1812),
.A2(n_1784),
.B1(n_1775),
.B2(n_1779),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_R g1818 ( 
.A(n_1803),
.B(n_1518),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1812),
.A2(n_1718),
.B(n_1771),
.C(n_1776),
.Y(n_1819)
);

OAI322xp33_ASAP7_75t_L g1820 ( 
.A1(n_1806),
.A2(n_1760),
.A3(n_1773),
.B1(n_1757),
.B2(n_1759),
.C1(n_1736),
.C2(n_1732),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1805),
.A2(n_1801),
.B1(n_1809),
.B2(n_1810),
.C(n_1773),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1808),
.A2(n_1761),
.B(n_1736),
.Y(n_1822)
);

NOR3x1_ASAP7_75t_L g1823 ( 
.A(n_1811),
.B(n_1759),
.C(n_1757),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1811),
.A2(n_1761),
.B(n_1779),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1813),
.A2(n_1816),
.B(n_1817),
.Y(n_1825)
);

OAI21xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1814),
.A2(n_1772),
.B(n_1734),
.Y(n_1826)
);

INVx5_ASAP7_75t_L g1827 ( 
.A(n_1823),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1824),
.A2(n_1822),
.B(n_1819),
.Y(n_1828)
);

INVxp67_ASAP7_75t_SL g1829 ( 
.A(n_1815),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1821),
.A2(n_1718),
.B1(n_1749),
.B2(n_1772),
.C(n_1729),
.Y(n_1830)
);

NAND5xp2_ASAP7_75t_L g1831 ( 
.A(n_1818),
.B(n_1734),
.C(n_1702),
.D(n_1698),
.E(n_1699),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1827),
.B(n_1744),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1828),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1827),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1829),
.B(n_1744),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1825),
.B(n_1698),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1831),
.B(n_1726),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1826),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1834),
.B(n_1830),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1833),
.A2(n_1820),
.B1(n_1625),
.B2(n_1705),
.C(n_1703),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1832),
.Y(n_1841)
);

NOR3xp33_ASAP7_75t_L g1842 ( 
.A(n_1838),
.B(n_1705),
.C(n_1702),
.Y(n_1842)
);

NAND2x1p5_ASAP7_75t_L g1843 ( 
.A(n_1836),
.B(n_1699),
.Y(n_1843)
);

NAND2xp33_ASAP7_75t_R g1844 ( 
.A(n_1835),
.B(n_1837),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1841),
.B(n_1717),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1843),
.A2(n_1839),
.B1(n_1844),
.B2(n_1842),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1840),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1846),
.B(n_1704),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1848),
.B(n_1845),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1847),
.B1(n_1696),
.B2(n_1681),
.Y(n_1850)
);

AO22x2_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1696),
.B1(n_1681),
.B2(n_1656),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1850),
.A2(n_1535),
.B1(n_1656),
.B2(n_1643),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1851),
.A2(n_1717),
.B(n_1647),
.Y(n_1853)
);

CKINVDCx20_ASAP7_75t_R g1854 ( 
.A(n_1852),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1853),
.B(n_1644),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1855),
.A2(n_1659),
.B1(n_1645),
.B2(n_1648),
.C(n_1661),
.Y(n_1856)
);

XNOR2xp5_ASAP7_75t_L g1857 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1647),
.B(n_1644),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1654),
.B1(n_1672),
.B2(n_1671),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1647),
.B1(n_1672),
.B2(n_1671),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1468),
.B(n_1467),
.C(n_1551),
.Y(n_1861)
);


endmodule