module fake_jpeg_9709_n_296 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_23),
.B1(n_21),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_67),
.B1(n_30),
.B2(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_17),
.C(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_34),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_17),
.C(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_24),
.B(n_31),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_63),
.B(n_18),
.C(n_20),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_31),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_65),
.B1(n_48),
.B2(n_60),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_75),
.B(n_69),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_93),
.B1(n_94),
.B2(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_92),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_25),
.B1(n_26),
.B2(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_28),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_26),
.B1(n_27),
.B2(n_42),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_100),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_92),
.B1(n_56),
.B2(n_59),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_119),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_55),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_114),
.C(n_116),
.Y(n_142)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_112),
.B1(n_117),
.B2(n_76),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_111),
.B1(n_54),
.B2(n_91),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_73),
.B1(n_91),
.B2(n_80),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_89),
.C(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_61),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_75),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_107),
.C(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_102),
.B1(n_117),
.B2(n_119),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_84),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_75),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_139),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_85),
.B1(n_66),
.B2(n_57),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_145),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_60),
.B1(n_64),
.B2(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_54),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_103),
.B(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_84),
.B1(n_68),
.B2(n_22),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_77),
.B1(n_91),
.B2(n_49),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_149),
.B(n_156),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_95),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_77),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_49),
.B(n_42),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_143),
.B(n_137),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_42),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_0),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_118),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_168),
.B(n_130),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_68),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_169),
.B(n_22),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_142),
.C(n_120),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_80),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_0),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_131),
.B(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_182),
.C(n_185),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_187),
.B1(n_195),
.B2(n_153),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_160),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_142),
.C(n_121),
.Y(n_182)
);

OA21x2_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_131),
.B(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_170),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_132),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_134),
.B1(n_133),
.B2(n_128),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_165),
.B1(n_169),
.B2(n_153),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_129),
.B1(n_127),
.B2(n_130),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_152),
.C(n_150),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_194),
.C(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_161),
.B(n_148),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_161),
.B(n_158),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_164),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_127),
.C(n_68),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_155),
.B1(n_156),
.B2(n_154),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_194),
.B1(n_177),
.B2(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_204),
.C(n_210),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_213),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_156),
.C(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_212),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_188),
.C(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_154),
.C(n_162),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_158),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_188),
.C(n_181),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_146),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_168),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_153),
.B1(n_127),
.B2(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_175),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_231),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_184),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_227),
.Y(n_247)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_235),
.C(n_202),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_179),
.B(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_173),
.C(n_179),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_173),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_201),
.B1(n_197),
.B2(n_198),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_204),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_244),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_227),
.B1(n_225),
.B2(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_210),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_242),
.C(n_248),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_230),
.B(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_246),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_215),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_213),
.C(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_1),
.C(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_1),
.Y(n_263)
);

XOR2x1_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_220),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_218),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_219),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_263),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_221),
.B1(n_245),
.B2(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_234),
.B1(n_232),
.B2(n_222),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_260),
.B1(n_242),
.B2(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_225),
.B(n_11),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_8),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_12),
.B(n_16),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_7),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_252),
.C(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_256),
.B(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_12),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_5),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_280),
.B(n_13),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_5),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_5),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_283),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_266),
.B(n_264),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_264),
.B(n_277),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_13),
.B(n_16),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_279),
.C(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_285),
.B(n_3),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_291),
.B(n_3),
.Y(n_294)
);

AOI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_1),
.A3(n_4),
.B1(n_292),
.B2(n_293),
.C(n_285),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_1),
.Y(n_296)
);


endmodule