module fake_jpeg_23266_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_3),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_17),
.B(n_18),
.Y(n_20)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_15),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_25),
.B1(n_8),
.B2(n_6),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_13),
.B(n_5),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_19),
.C(n_20),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_25),
.C(n_21),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_17),
.B1(n_11),
.B2(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_26),
.Y(n_31)
);

AOI221xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_29),
.B1(n_12),
.B2(n_1),
.C(n_0),
.Y(n_32)
);

AOI21x1_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_12),
.B(n_0),
.Y(n_33)
);


endmodule