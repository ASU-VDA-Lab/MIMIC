module fake_ariane_770_n_1633 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1633);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1633;

wire n_913;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_43),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_88),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_43),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_26),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_0),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_34),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_20),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_102),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_40),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_27),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_32),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_30),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_56),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_50),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_37),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_31),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_82),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_89),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_90),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_54),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_64),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_37),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_87),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_66),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_91),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_42),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_84),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_24),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_36),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_28),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_32),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_94),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_63),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_48),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_107),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_27),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_10),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_17),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_6),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_49),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_59),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_70),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_78),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_69),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_52),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_62),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_97),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_31),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_50),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_99),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_48),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_35),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_73),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_79),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_19),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_45),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_13),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_111),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_144),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_40),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_57),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_129),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_67),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_16),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_77),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_80),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_58),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_133),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_42),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_92),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_33),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_11),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_143),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_108),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_22),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_85),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_146),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_161),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_147),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_169),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_190),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_175),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_164),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_190),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_230),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_150),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_167),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_167),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_153),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_172),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_155),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_158),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_165),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_158),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_163),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_168),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_169),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_163),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_163),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_158),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_177),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_192),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_183),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_171),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_206),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_192),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_184),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_194),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_194),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_228),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_197),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_179),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_197),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_349),
.Y(n_355)
);

NAND2x1p5_ASAP7_75t_L g356 ( 
.A(n_285),
.B(n_198),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g359 ( 
.A(n_349),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_287),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_335),
.B1(n_344),
.B2(n_342),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_292),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_R g368 ( 
.A(n_303),
.B(n_186),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_293),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_285),
.B(n_231),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_314),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_294),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_286),
.B(n_261),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_286),
.B(n_193),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_295),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_288),
.B(n_179),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_288),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_289),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_289),
.Y(n_392)
);

AND3x2_ASAP7_75t_L g393 ( 
.A(n_318),
.B(n_176),
.C(n_148),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_291),
.B(n_203),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_291),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_296),
.A2(n_298),
.B(n_297),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_296),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_297),
.B(n_203),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_298),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_300),
.B(n_160),
.Y(n_403)
);

NAND2xp33_ASAP7_75t_L g404 ( 
.A(n_300),
.B(n_198),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_304),
.B(n_247),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_304),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_307),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_307),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_308),
.A2(n_218),
.B(n_195),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_309),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_301),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_310),
.B(n_171),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_310),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_350),
.B(n_229),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_320),
.B(n_234),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_397),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_377),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_377),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_323),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_395),
.B(n_305),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_306),
.Y(n_438)
);

CKINVDCx6p67_ASAP7_75t_R g439 ( 
.A(n_395),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_356),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_352),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_380),
.B(n_396),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_334),
.Y(n_452)
);

BUFx6f_ASAP7_75t_SL g453 ( 
.A(n_414),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_343),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_198),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_378),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_391),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_400),
.B(n_311),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_395),
.B(n_346),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_400),
.B(n_329),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_368),
.A2(n_269),
.B1(n_211),
.B2(n_248),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_369),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_313),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g477 ( 
.A(n_360),
.B(n_302),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_381),
.B(n_313),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_355),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

BUFx4f_ASAP7_75t_L g483 ( 
.A(n_356),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g485 ( 
.A(n_356),
.B(n_315),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_370),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_370),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_382),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_382),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_382),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_359),
.Y(n_494)
);

NOR2x1p5_ASAP7_75t_L g495 ( 
.A(n_366),
.B(n_341),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_409),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_405),
.B(n_315),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_359),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_372),
.A2(n_290),
.B1(n_330),
.B2(n_326),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_381),
.B(n_319),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_417),
.B(n_319),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_410),
.A2(n_322),
.B1(n_326),
.B2(n_325),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_417),
.B(n_322),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_389),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_383),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_389),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_389),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_374),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_374),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_374),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_413),
.B(n_341),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_410),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_374),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_368),
.A2(n_250),
.B1(n_243),
.B2(n_238),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_400),
.B(n_324),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_411),
.B(n_198),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_407),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_413),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_400),
.B(n_324),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_416),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_354),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_354),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_416),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_374),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_410),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_359),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_379),
.B(n_414),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_357),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_357),
.Y(n_547)
);

AND3x1_ASAP7_75t_L g548 ( 
.A(n_379),
.B(n_205),
.C(n_200),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_358),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_358),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_361),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_390),
.B(n_325),
.Y(n_552)
);

AND3x2_ASAP7_75t_L g553 ( 
.A(n_414),
.B(n_205),
.C(n_200),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_361),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_390),
.B(n_345),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_364),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_364),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_367),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_535),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_455),
.B(n_398),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_438),
.B(n_398),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_447),
.B(n_431),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_455),
.B(n_401),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_495),
.B(n_414),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_483),
.B(n_401),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_495),
.B(n_414),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_433),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_419),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_451),
.B(n_408),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_483),
.B(n_408),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_418),
.A2(n_404),
.B1(n_412),
.B2(n_399),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_514),
.B(n_362),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_504),
.B(n_412),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_537),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_362),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_510),
.B(n_394),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_473),
.B(n_394),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_399),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_465),
.B(n_393),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_448),
.B(n_359),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_393),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_468),
.A2(n_262),
.B1(n_283),
.B2(n_275),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_479),
.B(n_359),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_448),
.B(n_404),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_467),
.B(n_367),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_371),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_483),
.B(n_195),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_485),
.A2(n_373),
.B(n_371),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_463),
.B(n_373),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_463),
.B(n_482),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_483),
.B(n_218),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_462),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_439),
.B(n_345),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_439),
.A2(n_262),
.B1(n_275),
.B2(n_280),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_471),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_463),
.B(n_376),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_463),
.B(n_376),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_499),
.B(n_471),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_482),
.B(n_384),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_499),
.B(n_210),
.C(n_209),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_482),
.B(n_384),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_441),
.B(n_219),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_441),
.A2(n_199),
.B1(n_196),
.B2(n_208),
.Y(n_610)
);

AOI221xp5_ASAP7_75t_L g611 ( 
.A1(n_548),
.A2(n_258),
.B1(n_220),
.B2(n_227),
.C(n_210),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_212),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_SL g613 ( 
.A(n_482),
.B(n_209),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_525),
.Y(n_614)
);

INVx8_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_452),
.B(n_387),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_462),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_419),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_509),
.B(n_217),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_422),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_422),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_466),
.B(n_347),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_464),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_469),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_422),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_525),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_426),
.B(n_434),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_434),
.B(n_388),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_469),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_424),
.B(n_388),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_552),
.B(n_281),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_432),
.B(n_347),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_418),
.A2(n_280),
.B1(n_283),
.B2(n_258),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_480),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_509),
.B(n_219),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_509),
.B(n_235),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_480),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_509),
.B(n_222),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_531),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_474),
.B(n_475),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_420),
.B(n_235),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_421),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_420),
.A2(n_274),
.B(n_220),
.C(n_227),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_502),
.B(n_223),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_421),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_528),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_474),
.B(n_348),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_475),
.B(n_348),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_477),
.B(n_539),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_421),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_453),
.B(n_201),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_476),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_423),
.B(n_251),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_423),
.A2(n_239),
.B1(n_244),
.B2(n_278),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_476),
.B(n_351),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_478),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_478),
.B(n_351),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_481),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_494),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_534),
.B(n_353),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_550),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_538),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_481),
.B(n_353),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_501),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_484),
.B(n_188),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_224),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_555),
.B(n_226),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_507),
.B(n_157),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_428),
.A2(n_278),
.B(n_239),
.C(n_274),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_519),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_488),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_488),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_497),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_497),
.A2(n_251),
.B(n_259),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_533),
.B(n_236),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_428),
.B(n_259),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_430),
.B(n_149),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_498),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_498),
.B(n_188),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_501),
.B(n_241),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_430),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_450),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_506),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_450),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_517),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_517),
.B(n_244),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_521),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_521),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_550),
.B(n_242),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_501),
.B(n_201),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_523),
.B(n_256),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_524),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_524),
.B(n_270),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_550),
.B(n_270),
.C(n_273),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_546),
.B(n_255),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_546),
.B(n_263),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_435),
.A2(n_207),
.B(n_152),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_547),
.A2(n_213),
.B1(n_156),
.B2(n_162),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_547),
.B(n_268),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_446),
.B(n_151),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_519),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_425),
.B(n_271),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_446),
.B(n_166),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_519),
.B(n_170),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_446),
.B(n_173),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_549),
.B(n_276),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_553),
.B(n_157),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_425),
.B(n_201),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_549),
.B(n_174),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_542),
.B(n_2),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_425),
.B(n_267),
.C(n_266),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_559),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_672),
.A2(n_558),
.B1(n_557),
.B2(n_554),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_563),
.B(n_542),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_664),
.B(n_157),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_563),
.B(n_542),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_561),
.B(n_446),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_526),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_615),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_713),
.A2(n_650),
.B1(n_648),
.B2(n_588),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_565),
.B(n_526),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_R g727 ( 
.A(n_621),
.B(n_526),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_567),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_SL g729 ( 
.A(n_583),
.B(n_607),
.C(n_605),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_602),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_569),
.B(n_568),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_615),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_571),
.B(n_580),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_583),
.B(n_429),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_567),
.B(n_526),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_615),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_653),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_584),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_R g741 ( 
.A(n_576),
.B(n_536),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_674),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_646),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_579),
.B(n_429),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_585),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_642),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_581),
.B(n_582),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_573),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_599),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_617),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_623),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_573),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_666),
.B(n_551),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_715),
.B(n_446),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_625),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_654),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_626),
.Y(n_759)
);

OR2x2_ASAP7_75t_SL g760 ( 
.A(n_601),
.B(n_520),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_536),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_590),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_619),
.A2(n_445),
.B1(n_429),
.B2(n_440),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_631),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_686),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_693),
.A2(n_558),
.B(n_557),
.C(n_554),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_656),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_574),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_660),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_662),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_688),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_685),
.B(n_536),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_685),
.B(n_541),
.Y(n_773)
);

BUFx8_ASAP7_75t_SL g774 ( 
.A(n_634),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_601),
.B(n_446),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_628),
.Y(n_776)
);

NOR2x2_ASAP7_75t_L g777 ( 
.A(n_634),
.B(n_558),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_587),
.B(n_634),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_577),
.B(n_541),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_647),
.A2(n_673),
.B(n_560),
.C(n_564),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_573),
.Y(n_781)
);

NOR2x1p5_ASAP7_75t_L g782 ( 
.A(n_712),
.B(n_551),
.Y(n_782)
);

AO221x2_ASAP7_75t_L g783 ( 
.A1(n_588),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.C(n_12),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_597),
.A2(n_460),
.B(n_456),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_665),
.B(n_541),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_665),
.B(n_541),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_675),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_702),
.B(n_544),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_641),
.B(n_445),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_684),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_690),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_586),
.B(n_511),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_SL g793 ( 
.A(n_671),
.B(n_215),
.C(n_178),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_676),
.B(n_544),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_589),
.A2(n_460),
.B1(n_436),
.B2(n_437),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_573),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_544),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_682),
.Y(n_798)
);

BUFx4f_ASAP7_75t_L g799 ( 
.A(n_684),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_644),
.A2(n_544),
.B(n_456),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_612),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_687),
.B(n_489),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_655),
.B(n_694),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_648),
.A2(n_658),
.B1(n_635),
.B2(n_612),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_689),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_562),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_684),
.Y(n_807)
);

AND2x6_ASAP7_75t_SL g808 ( 
.A(n_670),
.B(n_436),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_570),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_611),
.B(n_489),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_610),
.B(n_511),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_624),
.B(n_520),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_699),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_691),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_658),
.A2(n_427),
.B1(n_508),
.B2(n_491),
.Y(n_815)
);

AND2x2_ASAP7_75t_SL g816 ( 
.A(n_635),
.B(n_520),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_637),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_693),
.A2(n_444),
.B1(n_437),
.B2(n_442),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_692),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_696),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_633),
.B(n_591),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_684),
.A2(n_458),
.B1(n_530),
.B2(n_508),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_616),
.B(n_489),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_637),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_651),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_700),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_703),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_618),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_663),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_663),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_663),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_704),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_670),
.A2(n_449),
.B1(n_442),
.B2(n_443),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_679),
.B(n_511),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_679),
.B(n_490),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_711),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_575),
.B(n_490),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_659),
.B(n_491),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_668),
.B(n_663),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_661),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_668),
.B(n_522),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_667),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_620),
.Y(n_845)
);

NOR2x2_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_522),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_622),
.Y(n_847)
);

INVx8_ASAP7_75t_L g848 ( 
.A(n_684),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_707),
.B(n_491),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_707),
.A2(n_443),
.B1(n_444),
.B2(n_449),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_695),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_592),
.B(n_492),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_697),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_681),
.A2(n_505),
.B(n_492),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_627),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_596),
.B(n_493),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_706),
.B(n_566),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_636),
.A2(n_180),
.B1(n_265),
.B2(n_264),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_566),
.B(n_513),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_640),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_572),
.B(n_513),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_R g862 ( 
.A(n_714),
.B(n_513),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_643),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_572),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_603),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_669),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_709),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_629),
.B(n_518),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_604),
.B(n_493),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_683),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_632),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_609),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_716),
.B(n_513),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_606),
.B(n_496),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_608),
.B(n_496),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_630),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_647),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_678),
.A2(n_540),
.B(n_527),
.C(n_496),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_645),
.B(n_505),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_593),
.B(n_515),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_705),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_717),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_838),
.B(n_593),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_733),
.A2(n_673),
.B(n_638),
.C(n_639),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_730),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_724),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_733),
.B(n_748),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_748),
.B(n_613),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_803),
.B(n_458),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_734),
.A2(n_598),
.B(n_639),
.C(n_638),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_744),
.B(n_598),
.Y(n_891)
);

O2A1O1Ixp5_ASAP7_75t_SL g892 ( 
.A1(n_722),
.A2(n_710),
.B(n_708),
.C(n_705),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_723),
.A2(n_708),
.B(n_710),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_731),
.B(n_515),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_821),
.A2(n_540),
.B(n_594),
.C(n_701),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_723),
.A2(n_657),
.B(n_645),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_724),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_730),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_738),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_729),
.B(n_540),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_828),
.B(n_515),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_779),
.A2(n_680),
.B(n_518),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_772),
.A2(n_516),
.B(n_512),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_762),
.B(n_450),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_729),
.B(n_454),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_724),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_732),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_804),
.A2(n_454),
.B(n_487),
.C(n_486),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_848),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_720),
.B(n_457),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_827),
.B(n_461),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_SL g912 ( 
.A(n_799),
.B(n_458),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_801),
.B(n_182),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_827),
.B(n_461),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_773),
.A2(n_470),
.B(n_486),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_762),
.A2(n_470),
.B(n_472),
.C(n_233),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_773),
.A2(n_470),
.B(n_472),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_874),
.A2(n_221),
.B(n_187),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_800),
.A2(n_530),
.B(n_458),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_834),
.B(n_185),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_871),
.B(n_530),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_874),
.A2(n_246),
.B(n_191),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_746),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_739),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_834),
.B(n_189),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_801),
.B(n_202),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_755),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_760),
.A2(n_214),
.B1(n_216),
.B2(n_232),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_728),
.B(n_732),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_875),
.A2(n_260),
.B(n_254),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_825),
.B(n_530),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_858),
.B(n_249),
.C(n_252),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_783),
.B(n_530),
.C(n_458),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_768),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_741),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_875),
.A2(n_800),
.B(n_856),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_805),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_732),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_737),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_736),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_826),
.B(n_458),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_842),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_780),
.A2(n_857),
.B(n_853),
.C(n_851),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_844),
.A2(n_813),
.B(n_836),
.C(n_814),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_856),
.A2(n_76),
.B(n_139),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_739),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_727),
.B(n_21),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_776),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_774),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_810),
.B(n_23),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_SL g951 ( 
.A(n_740),
.B(n_23),
.C(n_25),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_869),
.A2(n_81),
.B(n_135),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_869),
.A2(n_74),
.B(n_134),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_749),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_745),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_726),
.B(n_33),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_726),
.B(n_735),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_820),
.A2(n_34),
.B(n_38),
.C(n_39),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_747),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_SL g960 ( 
.A(n_793),
.B(n_39),
.C(n_41),
.Y(n_960)
);

INVx8_ASAP7_75t_L g961 ( 
.A(n_848),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_778),
.B(n_41),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_794),
.A2(n_103),
.B(n_131),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_793),
.B(n_44),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_750),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_877),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_791),
.B(n_47),
.Y(n_967)
);

AND2x2_ASAP7_75t_SL g968 ( 
.A(n_799),
.B(n_47),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_819),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_754),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_782),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_735),
.B(n_51),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_783),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_768),
.B(n_65),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_728),
.B(n_83),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_865),
.B(n_100),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_743),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_749),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_780),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_751),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_752),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_737),
.B(n_115),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_757),
.B(n_120),
.C(n_122),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_854),
.A2(n_124),
.B(n_142),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_749),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_766),
.A2(n_787),
.B(n_769),
.C(n_767),
.Y(n_986)
);

AOI222xp33_ASAP7_75t_L g987 ( 
.A1(n_759),
.A2(n_798),
.B1(n_770),
.B2(n_764),
.C1(n_775),
.C2(n_816),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_811),
.A2(n_837),
.B(n_795),
.C(n_835),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_876),
.B(n_761),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_792),
.A2(n_719),
.B(n_721),
.C(n_866),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_753),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_876),
.B(n_761),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_758),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_841),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_872),
.B(n_808),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_789),
.A2(n_873),
.B(n_797),
.C(n_794),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_870),
.A2(n_880),
.B(n_861),
.C(n_859),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_823),
.B(n_852),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_765),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_823),
.B(n_852),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_841),
.Y(n_1001)
);

NOR2xp67_ASAP7_75t_SL g1002 ( 
.A(n_754),
.B(n_807),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_872),
.A2(n_881),
.B(n_849),
.C(n_818),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_771),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_742),
.B(n_830),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_797),
.A2(n_788),
.B(n_840),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_756),
.A2(n_790),
.B1(n_864),
.B2(n_812),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_867),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_784),
.A2(n_786),
.B(n_785),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_806),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_984),
.A2(n_784),
.B(n_879),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_718),
.B1(n_802),
.B2(n_850),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_887),
.B(n_788),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_SL g1014 ( 
.A1(n_888),
.A2(n_785),
.B(n_786),
.Y(n_1014)
);

NAND3x1_ASAP7_75t_L g1015 ( 
.A(n_995),
.B(n_777),
.C(n_846),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_1009),
.A2(n_879),
.B(n_839),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_899),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_885),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_893),
.A2(n_840),
.A3(n_878),
.B(n_802),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_949),
.Y(n_1020)
);

NOR4xp25_ASAP7_75t_L g1021 ( 
.A(n_966),
.B(n_845),
.C(n_847),
.D(n_815),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_929),
.B(n_754),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_934),
.B(n_830),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_L g1024 ( 
.A(n_973),
.B(n_864),
.C(n_809),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_950),
.A2(n_822),
.B1(n_848),
.B2(n_763),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_962),
.B(n_806),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_864),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_937),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_988),
.A2(n_812),
.B(n_822),
.C(n_832),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_896),
.A2(n_901),
.B(n_998),
.Y(n_1030)
);

AOI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_966),
.A2(n_843),
.B1(n_862),
.B2(n_860),
.C(n_855),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_SL g1032 ( 
.A1(n_968),
.A2(n_860),
.B(n_832),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_892),
.A2(n_781),
.B(n_833),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_903),
.A2(n_781),
.B(n_833),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_888),
.B(n_796),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_943),
.A2(n_997),
.B(n_884),
.Y(n_1036)
);

AO22x2_ASAP7_75t_L g1037 ( 
.A1(n_928),
.A2(n_831),
.B1(n_817),
.B2(n_829),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_898),
.B(n_831),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_920),
.B(n_855),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_969),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1000),
.A2(n_996),
.B(n_890),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1000),
.A2(n_817),
.B(n_829),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_987),
.B(n_863),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_940),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_987),
.B(n_863),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1003),
.B(n_863),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_924),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_911),
.B(n_868),
.Y(n_1048)
);

NOR2xp67_ASAP7_75t_SL g1049 ( 
.A(n_946),
.B(n_796),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_915),
.A2(n_868),
.B(n_796),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_SL g1051 ( 
.A1(n_975),
.A2(n_824),
.B(n_868),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_914),
.B(n_868),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_1005),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1001),
.B(n_824),
.Y(n_1054)
);

OA22x2_ASAP7_75t_L g1055 ( 
.A1(n_1007),
.A2(n_928),
.B1(n_883),
.B2(n_971),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1010),
.B(n_994),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1001),
.B(n_955),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_919),
.A2(n_895),
.B(n_917),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_919),
.A2(n_963),
.B(n_986),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_959),
.B(n_965),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_945),
.A2(n_952),
.B(n_953),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_990),
.A2(n_976),
.B(n_905),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_980),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_R g1064 ( 
.A(n_948),
.B(n_1008),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_916),
.A2(n_908),
.A3(n_979),
.B(n_976),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_981),
.B(n_904),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_974),
.B(n_889),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_929),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_951),
.A2(n_900),
.B1(n_967),
.B2(n_933),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_926),
.A2(n_972),
.B(n_913),
.C(n_947),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_923),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_921),
.A2(n_931),
.A3(n_941),
.B(n_1004),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_SL g1073 ( 
.A(n_932),
.B(n_927),
.C(n_942),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_886),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_910),
.B(n_935),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_935),
.B(n_982),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_912),
.A2(n_944),
.B(n_889),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_977),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1002),
.A2(n_989),
.B(n_992),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_991),
.B(n_993),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_909),
.B(n_982),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_999),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_964),
.A2(n_894),
.B(n_925),
.C(n_930),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_918),
.A2(n_922),
.B(n_983),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_939),
.A2(n_897),
.B(n_938),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_939),
.A2(n_897),
.B(n_938),
.Y(n_1086)
);

INVx3_ASAP7_75t_SL g1087 ( 
.A(n_886),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_958),
.A2(n_957),
.B(n_956),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_SL g1089 ( 
.A1(n_960),
.A2(n_909),
.B(n_961),
.C(n_970),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_SL g1090 ( 
.A(n_961),
.B(n_907),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_954),
.B(n_978),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_906),
.B(n_978),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_985),
.A2(n_961),
.B(n_906),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_887),
.A2(n_723),
.B(n_733),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_887),
.B(n_733),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_893),
.A2(n_936),
.B(n_891),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_887),
.A2(n_723),
.B(n_733),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_899),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_887),
.A2(n_723),
.B(n_733),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_984),
.A2(n_1009),
.B(n_902),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_887),
.B(n_733),
.Y(n_1101)
);

OAI22x1_ASAP7_75t_L g1102 ( 
.A1(n_973),
.A2(n_528),
.B1(n_995),
.B2(n_416),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_934),
.B(n_664),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_887),
.A2(n_723),
.B(n_733),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_887),
.A2(n_723),
.B(n_733),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_924),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_899),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_984),
.A2(n_1009),
.B(n_902),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_934),
.B(n_664),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_563),
.B(n_561),
.C(n_733),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_887),
.B(n_733),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_968),
.A2(n_576),
.B1(n_532),
.B2(n_514),
.Y(n_1112)
);

OA21x2_ASAP7_75t_L g1113 ( 
.A1(n_1009),
.A2(n_936),
.B(n_893),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_893),
.A2(n_854),
.A3(n_936),
.B(n_896),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_936),
.A2(n_723),
.B(n_1006),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_887),
.B(n_733),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_899),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_936),
.A2(n_723),
.B(n_1006),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_887),
.B(n_733),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_984),
.A2(n_1009),
.B(n_902),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_961),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_936),
.A2(n_723),
.B(n_1006),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_887),
.B(n_733),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_984),
.A2(n_1009),
.B(n_902),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_887),
.B(n_733),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_893),
.A2(n_1009),
.B(n_936),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_882),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_984),
.A2(n_1009),
.B(n_902),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_887),
.A2(n_733),
.B1(n_804),
.B2(n_713),
.Y(n_1129)
);

AND2x2_ASAP7_75t_SL g1130 ( 
.A(n_968),
.B(n_803),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_924),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_887),
.A2(n_733),
.B1(n_804),
.B2(n_713),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1124),
.A2(n_1128),
.B(n_1096),
.Y(n_1134)
);

CKINVDCx16_ASAP7_75t_R g1135 ( 
.A(n_1064),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1011),
.A2(n_1058),
.B(n_1014),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1126),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1020),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_1071),
.Y(n_1139)
);

INVx6_ASAP7_75t_L g1140 ( 
.A(n_1121),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1058),
.A2(n_1061),
.B(n_1050),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1017),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1115),
.A2(n_1122),
.B(n_1118),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1098),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1115),
.A2(n_1122),
.B(n_1118),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_1073),
.B(n_1110),
.C(n_1024),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1056),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1036),
.A2(n_1059),
.B(n_1062),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1044),
.Y(n_1153)
);

AO32x2_ASAP7_75t_L g1154 ( 
.A1(n_1069),
.A2(n_1132),
.A3(n_1129),
.B1(n_1012),
.B2(n_1025),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1016),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_R g1157 ( 
.A(n_1043),
.B(n_1045),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1041),
.A2(n_1104),
.B(n_1094),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1026),
.B(n_1103),
.Y(n_1159)
);

INVx4_ASAP7_75t_SL g1160 ( 
.A(n_1076),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_1119),
.A2(n_1125),
.B(n_1123),
.C(n_1129),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1063),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1119),
.B(n_1123),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1081),
.B(n_1049),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1047),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1053),
.B(n_1107),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1127),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1125),
.B(n_1023),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1097),
.A2(n_1105),
.A3(n_1099),
.B(n_1025),
.Y(n_1169)
);

INVx5_ASAP7_75t_SL g1170 ( 
.A(n_1022),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1109),
.B(n_1075),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1075),
.B(n_1117),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1078),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1033),
.A2(n_1034),
.B(n_1030),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1082),
.Y(n_1175)
);

OAI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1112),
.A2(n_1070),
.B1(n_1036),
.B2(n_1031),
.C(n_1069),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1080),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1130),
.B(n_1038),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

OAI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1031),
.A2(n_1084),
.B1(n_1083),
.B2(n_1021),
.C(n_1039),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1087),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1046),
.A2(n_1029),
.A3(n_1052),
.B(n_1048),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1057),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1048),
.A2(n_1052),
.B(n_1046),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1042),
.A2(n_1113),
.B(n_1077),
.Y(n_1185)
);

BUFx2_ASAP7_75t_R g1186 ( 
.A(n_1043),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1013),
.A2(n_1067),
.B(n_1126),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1045),
.A2(n_1027),
.B(n_1066),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1057),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1028),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1085),
.A2(n_1086),
.B(n_1079),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1040),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1088),
.A2(n_1018),
.B(n_1032),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1121),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1066),
.A2(n_1051),
.B(n_1089),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1093),
.A2(n_1055),
.B(n_1091),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1076),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1037),
.A2(n_1054),
.B(n_1091),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1106),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1068),
.B(n_1076),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1092),
.A2(n_1074),
.B(n_1076),
.C(n_1131),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1114),
.A2(n_1015),
.B(n_1019),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1114),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1114),
.A2(n_1019),
.B(n_1072),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_SL g1205 ( 
.A(n_1076),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1019),
.A2(n_1065),
.B(n_1037),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1090),
.A2(n_973),
.B1(n_966),
.B2(n_1129),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1065),
.A2(n_1102),
.B1(n_783),
.B2(n_804),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1047),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_1113),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1095),
.B(n_887),
.Y(n_1211)
);

OAI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1112),
.A2(n_1110),
.B(n_973),
.C(n_725),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1016),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1016),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1059),
.A2(n_1118),
.B(n_1115),
.Y(n_1217)
);

NAND3x1_ASAP7_75t_L g1218 ( 
.A(n_1112),
.B(n_973),
.C(n_995),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1219)
);

NAND2x1_ASAP7_75t_L g1220 ( 
.A(n_1076),
.B(n_1051),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1115),
.A2(n_1122),
.B(n_1118),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1129),
.A2(n_1132),
.B1(n_1110),
.B2(n_966),
.C(n_601),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1017),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1115),
.A2(n_854),
.A3(n_1122),
.B(n_1118),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1016),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1129),
.A2(n_1132),
.B1(n_1110),
.B2(n_966),
.C(n_601),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1076),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1115),
.A2(n_1122),
.B(n_1118),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1060),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1110),
.A2(n_733),
.B1(n_1112),
.B2(n_725),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1102),
.A2(n_783),
.B1(n_804),
.B2(n_725),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1026),
.B(n_1103),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1102),
.A2(n_783),
.B1(n_804),
.B2(n_725),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1110),
.A2(n_1132),
.B(n_1129),
.C(n_973),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1060),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1060),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1110),
.A2(n_1132),
.B(n_1129),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1100),
.A2(n_1120),
.B(n_1108),
.Y(n_1244)
);

OAI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1129),
.A2(n_973),
.B1(n_966),
.B2(n_1132),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1026),
.B(n_1103),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1129),
.A2(n_1132),
.B1(n_1110),
.B2(n_966),
.C(n_601),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1135),
.A2(n_1139),
.B1(n_1181),
.B2(n_1176),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1212),
.A2(n_1236),
.B1(n_1232),
.B2(n_1231),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1171),
.B(n_1168),
.Y(n_1250)
);

AOI221x1_ASAP7_75t_SL g1251 ( 
.A1(n_1245),
.A2(n_1207),
.B1(n_1211),
.B2(n_1172),
.C(n_1152),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1137),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1200),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1178),
.B(n_1159),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1145),
.B(n_1152),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1160),
.B(n_1228),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1223),
.A2(n_1227),
.B(n_1247),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1209),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1235),
.B(n_1246),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1148),
.B(n_1142),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1147),
.A2(n_1212),
.B(n_1237),
.C(n_1207),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1224),
.B(n_1145),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1209),
.Y(n_1263)
);

O2A1O1Ixp5_ASAP7_75t_L g1264 ( 
.A1(n_1245),
.A2(n_1243),
.B(n_1237),
.C(n_1193),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1160),
.B(n_1228),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1138),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1156),
.B(n_1211),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1181),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1199),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1217),
.A2(n_1146),
.B(n_1143),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1227),
.B2(n_1223),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1144),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1156),
.B(n_1150),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1165),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1247),
.A2(n_1218),
.B1(n_1208),
.B2(n_1147),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1200),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1203),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1217),
.B(n_1161),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_L g1279 ( 
.A(n_1164),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1162),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1140),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_SL g1283 ( 
.A1(n_1163),
.A2(n_1221),
.B1(n_1219),
.B2(n_1167),
.C(n_1230),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1238),
.B(n_1241),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1183),
.B(n_1189),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1158),
.A2(n_1206),
.B(n_1141),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1208),
.A2(n_1180),
.B1(n_1186),
.B2(n_1164),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1160),
.B(n_1228),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1220),
.B(n_1197),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1185),
.A2(n_1136),
.B(n_1134),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1194),
.A2(n_1149),
.B1(n_1151),
.B2(n_1187),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1173),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1161),
.B(n_1195),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1154),
.B(n_1170),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1149),
.A2(n_1205),
.B1(n_1170),
.B2(n_1198),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1170),
.B(n_1184),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1210),
.A2(n_1184),
.B1(n_1226),
.B2(n_1155),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1210),
.A2(n_1216),
.B1(n_1155),
.B2(n_1214),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1175),
.A2(n_1188),
.B1(n_1201),
.B2(n_1226),
.C(n_1214),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1190),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1204),
.A2(n_1133),
.B(n_1244),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1182),
.B(n_1202),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1182),
.B(n_1169),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1192),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1196),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1222),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1229),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1201),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1157),
.A2(n_1191),
.B(n_1233),
.C(n_1213),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1157),
.A2(n_1239),
.B(n_1215),
.C(n_1242),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1174),
.B(n_1234),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1225),
.A2(n_1231),
.B(n_1110),
.C(n_1147),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1240),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1225),
.A2(n_1110),
.B(n_1031),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1145),
.B(n_1152),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1160),
.B(n_1228),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1223),
.A2(n_1110),
.B(n_1031),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1223),
.A2(n_1110),
.B(n_1031),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1178),
.B(n_1159),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1158),
.A2(n_1217),
.B(n_1207),
.Y(n_1322)
);

O2A1O1Ixp5_ASAP7_75t_L g1323 ( 
.A1(n_1212),
.A2(n_1245),
.B(n_1243),
.C(n_1207),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1178),
.B(n_1159),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1223),
.A2(n_1110),
.B(n_1031),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1145),
.B(n_1152),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1181),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_1217),
.B(n_1207),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1145),
.B(n_1152),
.Y(n_1329)
);

BUFx2_ASAP7_75t_SL g1330 ( 
.A(n_1310),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1313),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1294),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1252),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1323),
.A2(n_1261),
.B(n_1257),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1298),
.B(n_1304),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1292),
.B(n_1305),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1308),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1252),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1278),
.A2(n_1328),
.B(n_1322),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1313),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1262),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1277),
.B(n_1250),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1281),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1280),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1286),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1306),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1255),
.B(n_1317),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1310),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1285),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1271),
.A2(n_1249),
.B1(n_1275),
.B2(n_1288),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1283),
.B(n_1284),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1264),
.A2(n_1311),
.B(n_1312),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1259),
.B(n_1329),
.Y(n_1353)
);

AOI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1251),
.A2(n_1325),
.B1(n_1320),
.B2(n_1319),
.C(n_1314),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1296),
.B(n_1254),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1321),
.B(n_1324),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1311),
.A2(n_1312),
.B(n_1301),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1326),
.B(n_1273),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1267),
.B(n_1295),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1302),
.B(n_1307),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1293),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1295),
.B(n_1309),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1248),
.A2(n_1253),
.B1(n_1276),
.B2(n_1318),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1316),
.A2(n_1279),
.B(n_1297),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1309),
.A2(n_1299),
.B(n_1300),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1303),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1315),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1313),
.A2(n_1265),
.B(n_1256),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1303),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1260),
.B(n_1287),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1291),
.A2(n_1270),
.B(n_1287),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1287),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1256),
.B(n_1289),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1270),
.B(n_1291),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1368),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1362),
.B(n_1359),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1362),
.B(n_1270),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1333),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1332),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1366),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1359),
.B(n_1290),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1342),
.B(n_1336),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1370),
.B(n_1340),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1332),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1338),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1340),
.B(n_1327),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1348),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1345),
.B(n_1258),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1331),
.B(n_1289),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1342),
.B(n_1268),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1339),
.B(n_1318),
.Y(n_1391)
);

CKINVDCx14_ASAP7_75t_R g1392 ( 
.A(n_1356),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1339),
.B(n_1318),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1339),
.B(n_1265),
.Y(n_1394)
);

NOR2x1_ASAP7_75t_L g1395 ( 
.A(n_1361),
.B(n_1282),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1339),
.B(n_1265),
.Y(n_1396)
);

OAI31xp33_ASAP7_75t_L g1397 ( 
.A1(n_1350),
.A2(n_1334),
.A3(n_1354),
.B(n_1351),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1339),
.B(n_1282),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1373),
.B(n_1253),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1345),
.B(n_1263),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1341),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1397),
.B(n_1354),
.C(n_1350),
.Y(n_1402)
);

OAI31xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1395),
.A2(n_1394),
.A3(n_1396),
.B(n_1393),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1397),
.B(n_1334),
.C(n_1364),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1377),
.A2(n_1369),
.B(n_1365),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1399),
.B(n_1373),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1379),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1376),
.B(n_1351),
.C(n_1377),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1401),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1392),
.B(n_1358),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1401),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1392),
.A2(n_1330),
.B1(n_1361),
.B2(n_1363),
.Y(n_1413)
);

NAND4xp25_ASAP7_75t_L g1414 ( 
.A(n_1397),
.B(n_1347),
.C(n_1374),
.D(n_1367),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1375),
.A2(n_1337),
.B1(n_1346),
.B2(n_1349),
.C(n_1343),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1399),
.B(n_1373),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1383),
.B(n_1344),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1381),
.A2(n_1330),
.B1(n_1364),
.B2(n_1348),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1375),
.A2(n_1337),
.B1(n_1357),
.B2(n_1352),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1375),
.A2(n_1357),
.B1(n_1352),
.B2(n_1336),
.C(n_1360),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_SL g1421 ( 
.A(n_1399),
.B(n_1387),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1389),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1386),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1384),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1375),
.A2(n_1357),
.B1(n_1352),
.B2(n_1335),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_R g1426 ( 
.A(n_1390),
.B(n_1266),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1381),
.A2(n_1335),
.B1(n_1357),
.B2(n_1352),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1380),
.A2(n_1369),
.B(n_1365),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1382),
.B(n_1353),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1387),
.B(n_1348),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1378),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1384),
.Y(n_1432)
);

AOI31xp33_ASAP7_75t_L g1433 ( 
.A1(n_1395),
.A2(n_1356),
.A3(n_1355),
.B(n_1353),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1378),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1422),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1407),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1428),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1430),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1414),
.B(n_1431),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1403),
.B(n_1383),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_SL g1441 ( 
.A(n_1402),
.B(n_1398),
.C(n_1390),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1430),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1422),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1405),
.A2(n_1365),
.B(n_1371),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1383),
.Y(n_1445)
);

INVx4_ASAP7_75t_SL g1446 ( 
.A(n_1406),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1425),
.A2(n_1372),
.B(n_1374),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1424),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1424),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1432),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1434),
.Y(n_1451)
);

NOR3xp33_ASAP7_75t_L g1452 ( 
.A(n_1404),
.B(n_1400),
.C(n_1388),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1434),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1410),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1410),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1421),
.B(n_1391),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1412),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1421),
.B(n_1391),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1450),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1450),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1444),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1458),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1441),
.A2(n_1419),
.B1(n_1420),
.B2(n_1427),
.C(n_1408),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1448),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1452),
.B(n_1409),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1457),
.B(n_1433),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1452),
.B(n_1415),
.Y(n_1469)
);

OAI31xp33_ASAP7_75t_L g1470 ( 
.A1(n_1439),
.A2(n_1418),
.A3(n_1413),
.B(n_1398),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1441),
.A2(n_1411),
.B(n_1396),
.C(n_1394),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1457),
.B(n_1412),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1448),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1382),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1448),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1444),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1406),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1458),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1436),
.Y(n_1481)
);

AND2x2_ASAP7_75t_SL g1482 ( 
.A(n_1438),
.B(n_1352),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1438),
.B(n_1406),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1444),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1440),
.B(n_1456),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1442),
.B(n_1416),
.Y(n_1488)
);

NOR3xp33_ASAP7_75t_L g1489 ( 
.A(n_1454),
.B(n_1388),
.C(n_1400),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1457),
.A2(n_1405),
.B(n_1357),
.C(n_1398),
.Y(n_1491)
);

AND2x2_ASAP7_75t_SL g1492 ( 
.A(n_1442),
.B(n_1387),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1447),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1454),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1456),
.B(n_1459),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1455),
.B(n_1417),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1451),
.B(n_1385),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1451),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1483),
.B(n_1451),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1464),
.A2(n_1447),
.B1(n_1444),
.B2(n_1437),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1460),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1483),
.B(n_1453),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1494),
.B(n_1480),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1442),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1494),
.B(n_1453),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1494),
.B(n_1453),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1469),
.C(n_1468),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1482),
.B(n_1459),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1466),
.A2(n_1443),
.B(n_1445),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_R g1511 ( 
.A(n_1463),
.B(n_1266),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1463),
.B(n_1446),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1472),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1460),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1467),
.B(n_1447),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1467),
.B(n_1475),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1449),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1473),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1445),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1461),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1461),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1478),
.B(n_1443),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1481),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1481),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.B(n_1449),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1499),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1492),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1465),
.B(n_1447),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1435),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1465),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1517),
.B(n_1493),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1487),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1520),
.B(n_1497),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1504),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1501),
.A2(n_1471),
.B1(n_1493),
.B2(n_1487),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1508),
.A2(n_1493),
.B1(n_1447),
.B2(n_1470),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.B(n_1505),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1512),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1526),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1505),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1530),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1513),
.A2(n_1462),
.B(n_1477),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1526),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1516),
.A2(n_1493),
.B1(n_1479),
.B2(n_1484),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_SL g1553 ( 
.A(n_1510),
.B(n_1470),
.C(n_1496),
.Y(n_1553)
);

INVx3_ASAP7_75t_SL g1554 ( 
.A(n_1512),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1527),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1512),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1533),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1479),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1544),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

OAI21xp33_ASAP7_75t_L g1561 ( 
.A1(n_1539),
.A2(n_1509),
.B(n_1524),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1541),
.B(n_1524),
.Y(n_1562)
);

OAI32xp33_ASAP7_75t_L g1563 ( 
.A1(n_1538),
.A2(n_1531),
.A3(n_1500),
.B1(n_1503),
.B2(n_1519),
.Y(n_1563)
);

OAI222xp33_ASAP7_75t_L g1564 ( 
.A1(n_1545),
.A2(n_1519),
.B1(n_1515),
.B2(n_1523),
.C1(n_1503),
.C2(n_1500),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1553),
.A2(n_1477),
.B1(n_1462),
.B2(n_1486),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1556),
.B(n_1521),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1550),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1550),
.Y(n_1568)
);

OAI31xp33_ASAP7_75t_L g1569 ( 
.A1(n_1551),
.A2(n_1486),
.A3(n_1485),
.B(n_1521),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1555),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1555),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1545),
.A2(n_1476),
.B(n_1474),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1537),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1542),
.B(n_1502),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1557),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_L g1578 ( 
.A(n_1566),
.B(n_1554),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1562),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1566),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1562),
.B(n_1556),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1576),
.B(n_1546),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1559),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1564),
.B(n_1541),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1542),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1572),
.B(n_1540),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1564),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_SL g1589 ( 
.A(n_1584),
.B(n_1569),
.C(n_1561),
.Y(n_1589)
);

AND4x1_ASAP7_75t_L g1590 ( 
.A(n_1584),
.B(n_1536),
.C(n_1547),
.D(n_1574),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1588),
.A2(n_1563),
.B(n_1573),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1588),
.A2(n_1565),
.B(n_1558),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1581),
.B(n_1543),
.Y(n_1595)
);

NAND2xp33_ASAP7_75t_R g1596 ( 
.A(n_1587),
.B(n_1558),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1578),
.A2(n_1558),
.B(n_1560),
.Y(n_1597)
);

NAND4xp25_ASAP7_75t_L g1598 ( 
.A(n_1582),
.B(n_1543),
.C(n_1558),
.D(n_1571),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1585),
.A2(n_1549),
.B(n_1532),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1593),
.A2(n_1580),
.B(n_1586),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1591),
.A2(n_1583),
.B1(n_1554),
.B2(n_1568),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1598),
.B(n_1567),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1592),
.A2(n_1543),
.B1(n_1534),
.B2(n_1549),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1594),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1603),
.B(n_1590),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1604),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1601),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1600),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1602),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1604),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1609),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1608),
.A2(n_1589),
.B(n_1597),
.C(n_1599),
.Y(n_1612)
);

AOI21xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1608),
.A2(n_1596),
.B(n_1595),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1610),
.A2(n_1548),
.B1(n_1570),
.B2(n_1534),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1606),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1611),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1615),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1614),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_L g1619 ( 
.A(n_1616),
.B(n_1613),
.C(n_1612),
.Y(n_1619)
);

OAI32xp33_ASAP7_75t_L g1620 ( 
.A1(n_1619),
.A2(n_1617),
.A3(n_1605),
.B1(n_1607),
.B2(n_1618),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1620),
.B(n_1515),
.Y(n_1621)
);

NAND2x1_ASAP7_75t_SL g1622 ( 
.A(n_1621),
.B(n_1532),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1622),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1623),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1623),
.A2(n_1269),
.B1(n_1272),
.B2(n_1274),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1624),
.A2(n_1625),
.B1(n_1548),
.B2(n_1485),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1624),
.B(n_1548),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1627),
.A2(n_1269),
.B1(n_1272),
.B2(n_1525),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1626),
.A2(n_1523),
.B1(n_1522),
.B2(n_1527),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1628),
.A2(n_1528),
.B1(n_1474),
.B2(n_1476),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1629),
.A2(n_1528),
.B1(n_1525),
.B2(n_1490),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1630),
.A2(n_1479),
.B1(n_1484),
.B2(n_1488),
.C(n_1490),
.Y(n_1632)
);

AOI211xp5_ASAP7_75t_L g1633 ( 
.A1(n_1632),
.A2(n_1631),
.B(n_1488),
.C(n_1484),
.Y(n_1633)
);


endmodule