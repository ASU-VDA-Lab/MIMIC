module fake_aes_8276_n_272 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_272, n_955);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_272;
output n_955;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_937;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_822;
wire n_706;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_948;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_58), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_110), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_64), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_56), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_43), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_31), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_16), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_50), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_28), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_25), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_55), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_111), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_87), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_70), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_76), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_93), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_3), .Y(n_133) );
NOR2xp67_ASAP7_75t_L g134 ( .A(n_77), .B(n_21), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_54), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_65), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_75), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_52), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_44), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_60), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_101), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_4), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_106), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_66), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_12), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_8), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_72), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_68), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_7), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_84), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_104), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_48), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_8), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_39), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_145), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
BUFx12f_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx5_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_153), .B(n_0), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_124), .A2(n_45), .B(n_108), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_145), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_148), .A2(n_154), .B(n_119), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
CKINVDCx11_ASAP7_75t_R g174 ( .A(n_142), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_118), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_146), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_172), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_172), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_171), .B(n_116), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_175), .B(n_135), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_170), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_177), .A2(n_133), .B1(n_112), .B2(n_134), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_172), .B(n_125), .C(n_126), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_173), .B(n_113), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_173), .B(n_113), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_158), .B(n_115), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_164), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_164), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_163), .B(n_115), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_176), .B(n_117), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_176), .B(n_117), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
INVx5_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_170), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_170), .B(n_120), .Y(n_214) );
INVxp33_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_158), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_157), .B(n_160), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
BUFx10_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_168), .B(n_140), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_220), .B(n_120), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_223), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_225), .Y(n_231) );
NOR3xp33_ASAP7_75t_L g232 ( .A(n_191), .B(n_177), .C(n_156), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_185), .B(n_129), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_225), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_185), .B(n_129), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_225), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_194), .B(n_168), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_225), .B(n_132), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_195), .B(n_132), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_207), .B(n_136), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_208), .B(n_136), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
BUFx10_ASAP7_75t_L g244 ( .A(n_197), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_183), .B(n_169), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_206), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g247 ( .A(n_209), .B(n_138), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_211), .B(n_169), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_206), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_211), .A2(n_167), .B1(n_156), .B2(n_143), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_214), .B(n_138), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_179), .B(n_141), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_206), .B(n_141), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_206), .B(n_143), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_200), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_212), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_193), .B(n_150), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_193), .A2(n_167), .B1(n_150), .B2(n_152), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_200), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_193), .B(n_151), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_202), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_193), .B(n_151), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_192), .A2(n_166), .B(n_144), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_202), .B(n_152), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_203), .B(n_166), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_203), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_205), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_212), .B(n_127), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_226), .A2(n_130), .B1(n_131), .B2(n_140), .Y(n_270) );
BUFx8_ASAP7_75t_L g271 ( .A(n_215), .Y(n_271) );
UNKNOWN g272 ( );
INVx2_ASAP7_75t_SL g273 ( .A(n_205), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_179), .B(n_147), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g275 ( .A(n_227), .B(n_114), .C(n_137), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_180), .B(n_5), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_212), .B(n_161), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_186), .A2(n_162), .B1(n_165), .B2(n_9), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_227), .B(n_165), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_186), .B(n_6), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_189), .B(n_165), .Y(n_282) );
INVx8_ASAP7_75t_L g283 ( .A(n_228), .Y(n_283) );
BUFx6f_ASAP7_75t_SL g284 ( .A(n_227), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_189), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_227), .B(n_228), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_228), .B(n_165), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_228), .B(n_165), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_216), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_217), .B(n_165), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_217), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_217), .Y(n_292) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_216), .B(n_7), .C(n_9), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_236), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_248), .B(n_218), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_265), .B(n_218), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_246), .A2(n_219), .B(n_221), .C(n_224), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_287), .A2(n_224), .B(n_221), .Y(n_299) );
AO21x1_ASAP7_75t_L g300 ( .A1(n_275), .A2(n_219), .B(n_182), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_288), .A2(n_224), .B(n_221), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_293), .A2(n_218), .B(n_213), .C(n_199), .Y(n_302) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_286), .A2(n_213), .B(n_182), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_278), .A2(n_213), .B(n_182), .Y(n_304) );
OAI321xp33_ASAP7_75t_L g305 ( .A1(n_251), .A2(n_196), .A3(n_184), .B1(n_187), .B2(n_188), .C(n_190), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_230), .B(n_10), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_236), .Y(n_308) );
AO32x1_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_196), .A3(n_184), .B1(n_187), .B2(n_188), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_233), .B(n_10), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_293), .A2(n_184), .B(n_187), .C(n_188), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_249), .A2(n_190), .B(n_196), .C(n_199), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_236), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_235), .B(n_11), .Y(n_314) );
BUFx4f_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_259), .B(n_11), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_256), .B(n_12), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_281), .A2(n_199), .B1(n_190), .B2(n_210), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_249), .A2(n_13), .B(n_14), .C(n_15), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_234), .B(n_210), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_234), .B(n_210), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_231), .B(n_210), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_278), .A2(n_210), .B(n_204), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_243), .A2(n_210), .B1(n_14), .B2(n_16), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_250), .A2(n_210), .B(n_204), .C(n_201), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_267), .B(n_13), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_243), .B(n_17), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_242), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_238), .B(n_204), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_264), .A2(n_204), .B(n_201), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_232), .A2(n_204), .B1(n_201), .B2(n_198), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_286), .A2(n_204), .B(n_201), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_201), .B(n_198), .Y(n_334) );
AOI21x1_ASAP7_75t_L g335 ( .A1(n_266), .A2(n_274), .B(n_290), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_229), .B(n_201), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_232), .A2(n_198), .B1(n_181), .B2(n_19), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_263), .B(n_198), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_280), .A2(n_198), .B(n_181), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_260), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_245), .B(n_17), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_244), .B(n_18), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_245), .B(n_18), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_251), .A2(n_198), .B1(n_181), .B2(n_21), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_263), .B(n_19), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_280), .A2(n_181), .B(n_67), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_331), .A2(n_276), .B(n_279), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_319), .A2(n_237), .B(n_268), .C(n_262), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_304), .A2(n_283), .B(n_253), .Y(n_349) );
AOI221x1_ASAP7_75t_L g350 ( .A1(n_325), .A2(n_275), .B1(n_285), .B2(n_254), .C(n_237), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_315), .B(n_270), .Y(n_351) );
AOI21xp5_ASAP7_75t_SL g352 ( .A1(n_318), .A2(n_284), .B(n_277), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_295), .B(n_255), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_315), .B(n_247), .Y(n_354) );
AO31x2_ASAP7_75t_L g355 ( .A1(n_300), .A2(n_277), .A3(n_257), .B(n_289), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_302), .A2(n_252), .B(n_240), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_307), .A2(n_284), .B1(n_261), .B2(n_258), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_307), .B(n_239), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_303), .A2(n_282), .B(n_292), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g361 ( .A(n_337), .B(n_279), .C(n_271), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g362 ( .A1(n_328), .A2(n_241), .B(n_269), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_292), .B(n_283), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_339), .A2(n_283), .B(n_291), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_295), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_319), .A2(n_181), .B(n_244), .C(n_20), .Y(n_366) );
OAI21x1_ASAP7_75t_SL g367 ( .A1(n_308), .A2(n_20), .B(n_22), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_296), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_310), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_314), .Y(n_372) );
BUFx8_ASAP7_75t_L g373 ( .A(n_294), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_333), .A2(n_181), .B(n_23), .Y(n_374) );
NOR2xp33_ASAP7_75t_SL g375 ( .A(n_308), .B(n_22), .Y(n_375) );
NAND2xp33_ASAP7_75t_L g376 ( .A(n_306), .B(n_24), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_334), .A2(n_26), .B(n_27), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_316), .B(n_29), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_302), .A2(n_30), .B(n_32), .C(n_33), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_369), .Y(n_381) );
CKINVDCx14_ASAP7_75t_R g382 ( .A(n_370), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_373), .Y(n_383) );
AO21x1_ASAP7_75t_L g384 ( .A1(n_376), .A2(n_311), .B(n_345), .Y(n_384) );
AOI221x1_ASAP7_75t_SL g385 ( .A1(n_368), .A2(n_342), .B1(n_343), .B2(n_341), .C(n_317), .Y(n_385) );
CKINVDCx6p67_ASAP7_75t_R g386 ( .A(n_365), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_364), .A2(n_332), .B(n_337), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_311), .B(n_332), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_360), .A2(n_309), .B(n_338), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_348), .A2(n_298), .A3(n_346), .B(n_326), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_375), .B(n_313), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_361), .A2(n_344), .B1(n_327), .B2(n_313), .Y(n_395) );
INVx6_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
CKINVDCx11_ASAP7_75t_R g397 ( .A(n_353), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_347), .A2(n_312), .B(n_305), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_312), .B(n_336), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_374), .A2(n_299), .B(n_301), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_353), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_374), .A2(n_330), .B(n_324), .Y(n_404) );
AO21x2_ASAP7_75t_L g405 ( .A1(n_379), .A2(n_297), .B(n_309), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_358), .B(n_306), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_351), .A2(n_329), .B1(n_323), .B2(n_321), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_309), .B(n_320), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_363), .A2(n_34), .B(n_35), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_391), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_390), .A2(n_347), .B(n_377), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_380), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_391), .B(n_355), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_401), .B(n_354), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_391), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_391), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_402), .B(n_355), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_408), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_408), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_385), .A2(n_366), .B1(n_357), .B2(n_362), .C(n_356), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_409), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_409), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_389), .B(n_355), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_379), .B(n_366), .Y(n_435) );
INVx8_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_385), .B(n_355), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_380), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_389), .B(n_377), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_380), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_380), .B(n_359), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_388), .B(n_378), .Y(n_450) );
OAI21x1_ASAP7_75t_L g451 ( .A1(n_390), .A2(n_349), .B(n_352), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_386), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_396), .B(n_376), .Y(n_453) );
AO22x1_ASAP7_75t_L g454 ( .A1(n_388), .A2(n_367), .B1(n_350), .B2(n_38), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_423), .B(n_398), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_423), .B(n_388), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_396), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_410), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_452), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_452), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_452), .B(n_382), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_412), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_405), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_452), .B(n_383), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_452), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_439), .B(n_392), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_421), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_418), .B(n_392), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_418), .B(n_392), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_383), .B(n_392), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_456), .B(n_383), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_424), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_432), .B(n_405), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_456), .B(n_397), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_432), .B(n_405), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_411), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_417), .B(n_405), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_428), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_456), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_417), .B(n_393), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_417), .B(n_444), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_411), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_414), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_436), .B(n_403), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_416), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_419), .B(n_394), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_436), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
INVx3_ASAP7_75t_SL g505 ( .A(n_436), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_420), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_436), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_419), .B(n_404), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_411), .B(n_393), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_437), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_444), .B(n_393), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_414), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_436), .Y(n_514) );
INVx5_ASAP7_75t_L g515 ( .A(n_419), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_448), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_450), .A2(n_395), .B1(n_407), .B2(n_384), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_455), .B(n_393), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_415), .B(n_393), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_446), .B(n_404), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_415), .B(n_393), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_455), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_414), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_443), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_420), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_415), .B(n_384), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_433), .B(n_404), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_450), .B(n_400), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_443), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_445), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_427), .B(n_400), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_446), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_493), .B(n_447), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_488), .B(n_445), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_491), .B(n_453), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_493), .B(n_447), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_534), .B(n_446), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_492), .B(n_449), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_496), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_461), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_449), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_494), .B(n_449), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_494), .B(n_447), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_478), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_505), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_487), .B(n_442), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_534), .B(n_420), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_521), .B(n_425), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_487), .B(n_441), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_471), .B(n_441), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_460), .B(n_453), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_462), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_471), .B(n_441), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_465), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_458), .B(n_442), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_505), .A2(n_427), .B1(n_453), .B2(n_429), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_458), .B(n_442), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_482), .B(n_425), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_482), .B(n_425), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_468), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_466), .B(n_435), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_470), .B(n_435), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_474), .B(n_454), .C(n_431), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_475), .B(n_435), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_485), .B(n_426), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_498), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_485), .B(n_426), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_464), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_513), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_484), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_457), .B(n_426), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_468), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_528), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_476), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_477), .B(n_435), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_457), .B(n_434), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_504), .B(n_435), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_459), .B(n_434), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_459), .B(n_434), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_521), .B(n_451), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_512), .B(n_440), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_521), .B(n_451), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_440), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_520), .B(n_440), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_503), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_520), .B(n_438), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_510), .B(n_511), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_517), .B(n_454), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_522), .B(n_438), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_525), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_522), .B(n_438), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_464), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_515), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_474), .B(n_431), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_527), .B(n_430), .Y(n_604) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_515), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_531), .B(n_430), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_489), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_527), .B(n_429), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_472), .B(n_451), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_469), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_518), .B(n_413), .C(n_400), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_497), .Y(n_613) );
NOR2xp67_ASAP7_75t_L g614 ( .A(n_501), .B(n_36), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_480), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_495), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_524), .B(n_413), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_515), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_516), .B(n_413), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_509), .B(n_37), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_509), .B(n_40), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_500), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_500), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_506), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_532), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_524), .B(n_41), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_519), .B(n_42), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_516), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_507), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_530), .B(n_46), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_529), .B(n_47), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_463), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_463), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_507), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_467), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_501), .B(n_49), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_506), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_526), .B(n_51), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_467), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_582), .B(n_529), .Y(n_640) );
AND3x1_ASAP7_75t_L g641 ( .A(n_581), .B(n_483), .C(n_479), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_575), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_535), .B(n_486), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_575), .B(n_515), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_583), .B(n_533), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_599), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_604), .B(n_608), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_559), .Y(n_648) );
BUFx2_ASAP7_75t_L g649 ( .A(n_601), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_535), .B(n_526), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_561), .Y(n_651) );
NOR2xp33_ASAP7_75t_SL g652 ( .A(n_605), .B(n_501), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_604), .B(n_508), .Y(n_653) );
NAND2x1_ASAP7_75t_L g654 ( .A(n_581), .B(n_514), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_538), .B(n_486), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_577), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_601), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_538), .B(n_486), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_540), .B(n_486), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_567), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_581), .B(n_508), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_605), .Y(n_662) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_551), .B(n_514), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_608), .B(n_473), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_558), .B(n_486), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_542), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_540), .B(n_502), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_544), .B(n_502), .Y(n_668) );
NAND2x1_ASAP7_75t_SL g669 ( .A(n_618), .B(n_514), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_618), .B(n_508), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_567), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_544), .B(n_502), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_579), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_545), .Y(n_674) );
NAND2x1_ASAP7_75t_L g675 ( .A(n_618), .B(n_499), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_548), .Y(n_676) );
OR2x6_ASAP7_75t_L g677 ( .A(n_605), .B(n_490), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_569), .B(n_490), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_615), .B(n_53), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_571), .B(n_59), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_549), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_585), .B(n_61), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_546), .B(n_62), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_556), .B(n_63), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_546), .B(n_69), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_547), .B(n_71), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_547), .B(n_73), .Y(n_687) );
NAND2x1_ASAP7_75t_L g688 ( .A(n_605), .B(n_74), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_556), .B(n_78), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_560), .B(n_79), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_560), .B(n_80), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_552), .B(n_81), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_550), .B(n_82), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_539), .B(n_83), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_557), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_598), .B(n_85), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_565), .B(n_86), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_595), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_552), .B(n_88), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_565), .B(n_566), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_555), .B(n_89), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_555), .B(n_90), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_541), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_566), .B(n_92), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_562), .B(n_95), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_572), .B(n_96), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_541), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_572), .B(n_98), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_574), .B(n_99), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_579), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_543), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_593), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_543), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_574), .B(n_100), .Y(n_714) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_614), .B(n_102), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_611), .B(n_103), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_562), .B(n_105), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_568), .B(n_107), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_109), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_573), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_576), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_564), .B(n_580), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_625), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_616), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_589), .B(n_591), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g726 ( .A(n_605), .B(n_602), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_607), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_603), .B(n_578), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_589), .B(n_591), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_606), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_539), .B(n_602), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_607), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_578), .B(n_584), .Y(n_733) );
OA211x2_ASAP7_75t_L g734 ( .A1(n_628), .A2(n_570), .B(n_626), .C(n_596), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_537), .B(n_594), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_613), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_536), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_610), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_586), .B(n_587), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_586), .B(n_587), .Y(n_740) );
AND2x4_ASAP7_75t_SL g741 ( .A(n_539), .B(n_621), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_610), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_584), .B(n_600), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_619), .B(n_554), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_592), .B(n_600), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_592), .B(n_594), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_597), .B(n_624), .Y(n_747) );
OR2x6_ASAP7_75t_L g748 ( .A(n_654), .B(n_636), .Y(n_748) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_675), .B(n_629), .Y(n_749) );
OR2x2_ASAP7_75t_L g750 ( .A(n_745), .B(n_597), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_645), .B(n_623), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_649), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_745), .B(n_609), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_645), .B(n_624), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_646), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_657), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_725), .B(n_554), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_731), .B(n_588), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_648), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_729), .B(n_554), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_743), .B(n_617), .Y(n_761) );
AOI32xp33_ASAP7_75t_L g762 ( .A1(n_641), .A2(n_634), .A3(n_563), .B1(n_621), .B2(n_620), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_746), .B(n_588), .Y(n_763) );
OR2x2_ASAP7_75t_L g764 ( .A(n_743), .B(n_637), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_737), .B(n_553), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_730), .B(n_637), .Y(n_766) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_694), .B(n_620), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_700), .B(n_623), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_733), .B(n_622), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_739), .B(n_588), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_651), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_731), .B(n_590), .Y(n_772) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_642), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_698), .B(n_622), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_723), .B(n_553), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_722), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_656), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_740), .B(n_590), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_667), .B(n_590), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_724), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_736), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_644), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_668), .B(n_619), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_720), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_741), .A2(n_631), .B1(n_636), .B2(n_619), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_650), .Y(n_786) );
NAND3xp33_ASAP7_75t_SL g787 ( .A(n_652), .B(n_636), .C(n_631), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_672), .B(n_553), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_666), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_733), .B(n_633), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_643), .B(n_632), .Y(n_791) );
NOR2x1p5_ASAP7_75t_L g792 ( .A(n_688), .B(n_612), .Y(n_792) );
AND2x2_ASAP7_75t_SL g793 ( .A(n_641), .B(n_630), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_728), .B(n_639), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_647), .B(n_635), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_647), .B(n_627), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_734), .A2(n_630), .B1(n_638), .B2(n_721), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_728), .B(n_638), .Y(n_798) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_662), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_674), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_655), .B(n_659), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_735), .B(n_747), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_712), .B(n_744), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_747), .B(n_653), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_676), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_712), .B(n_744), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_658), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_681), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_695), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_703), .B(n_713), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_653), .B(n_640), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_664), .B(n_678), .Y(n_812) );
BUFx3_ASAP7_75t_L g813 ( .A(n_663), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_644), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_661), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_661), .B(n_670), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_707), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_711), .Y(n_818) );
NOR2x1_ASAP7_75t_L g819 ( .A(n_677), .B(n_662), .Y(n_819) );
OR2x2_ASAP7_75t_L g820 ( .A(n_678), .B(n_665), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_738), .B(n_742), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_669), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_670), .B(n_727), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_660), .B(n_710), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_671), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_673), .Y(n_826) );
AOI21xp33_ASAP7_75t_L g827 ( .A1(n_679), .A2(n_718), .B(n_680), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_732), .B(n_677), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_693), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_677), .B(n_686), .Y(n_830) );
NOR2x1_ASAP7_75t_L g831 ( .A(n_694), .B(n_715), .Y(n_831) );
NAND3x1_ASAP7_75t_L g832 ( .A(n_652), .B(n_687), .C(n_685), .Y(n_832) );
NOR2xp33_ASAP7_75t_SL g833 ( .A(n_822), .B(n_726), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_L g834 ( .A1(n_784), .A2(n_718), .B(n_716), .C(n_682), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_774), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_774), .Y(n_836) );
INVx2_ASAP7_75t_SL g837 ( .A(n_813), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_766), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_766), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_794), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_793), .A2(n_726), .B(n_701), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_749), .A2(n_690), .B(n_692), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_787), .A2(n_734), .B1(n_683), .B2(n_702), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g844 ( .A1(n_749), .A2(n_684), .B(n_717), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_794), .Y(n_845) );
INVx2_ASAP7_75t_SL g846 ( .A(n_803), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_751), .B(n_680), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_810), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_806), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_810), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_762), .A2(n_682), .B1(n_696), .B2(n_691), .C(n_689), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_816), .B(n_699), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_824), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_773), .Y(n_854) );
OAI21xp33_ASAP7_75t_L g855 ( .A1(n_797), .A2(n_706), .B(n_714), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_753), .B(n_708), .Y(n_856) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_827), .B(n_697), .C(n_704), .D(n_709), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_785), .A2(n_693), .B1(n_705), .B2(n_719), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_751), .B(n_754), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_821), .Y(n_860) );
INVx2_ASAP7_75t_SL g861 ( .A(n_757), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_785), .A2(n_832), .B1(n_829), .B2(n_776), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_821), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_820), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_795), .Y(n_865) );
OR2x2_ASAP7_75t_L g866 ( .A(n_761), .B(n_802), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_764), .Y(n_867) );
AOI21xp33_ASAP7_75t_L g868 ( .A1(n_831), .A2(n_781), .B(n_827), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_790), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_769), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_755), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_759), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_754), .B(n_818), .Y(n_873) );
INVx1_ASAP7_75t_SL g874 ( .A(n_822), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_748), .A2(n_831), .B(n_819), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_771), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_817), .B(n_780), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_777), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_825), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_804), .B(n_811), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_789), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_823), .A2(n_798), .B1(n_772), .B2(n_758), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_763), .B(n_770), .Y(n_883) );
OAI322xp33_ASAP7_75t_L g884 ( .A1(n_862), .A2(n_796), .A3(n_812), .B1(n_775), .B2(n_765), .C1(n_750), .C2(n_752), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_848), .B(n_809), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_850), .B(n_800), .Y(n_886) );
OAI21xp33_ASAP7_75t_L g887 ( .A1(n_868), .A2(n_775), .B(n_756), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_859), .B(n_768), .Y(n_888) );
O2A1O1Ixp33_ASAP7_75t_SL g889 ( .A1(n_837), .A2(n_815), .B(n_782), .C(n_814), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_873), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_860), .B(n_808), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_874), .B(n_815), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_854), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_859), .B(n_786), .Y(n_894) );
AND2x2_ASAP7_75t_SL g895 ( .A(n_833), .B(n_758), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_873), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_849), .B(n_778), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_864), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_841), .A2(n_767), .B1(n_748), .B2(n_814), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_840), .B(n_805), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g901 ( .A1(n_841), .A2(n_868), .B1(n_875), .B2(n_851), .C(n_855), .Y(n_901) );
INVx2_ASAP7_75t_SL g902 ( .A(n_846), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g903 ( .A1(n_843), .A2(n_748), .B1(n_782), .B2(n_819), .Y(n_903) );
INVxp67_ASAP7_75t_L g904 ( .A(n_877), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_842), .A2(n_799), .B(n_772), .Y(n_905) );
INVx2_ASAP7_75t_SL g906 ( .A(n_861), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_863), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_877), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_835), .Y(n_909) );
OAI21xp33_ASAP7_75t_L g910 ( .A1(n_882), .A2(n_791), .B(n_828), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g911 ( .A1(n_842), .A2(n_807), .B1(n_830), .B2(n_826), .C(n_779), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g912 ( .A(n_901), .B(n_834), .C(n_857), .Y(n_912) );
NOR4xp25_ASAP7_75t_SL g913 ( .A(n_889), .B(n_845), .C(n_881), .D(n_872), .Y(n_913) );
OAI221xp5_ASAP7_75t_L g914 ( .A1(n_899), .A2(n_844), .B1(n_858), .B2(n_847), .C(n_839), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_899), .A2(n_844), .B(n_847), .Y(n_915) );
AOI211xp5_ASAP7_75t_SL g916 ( .A1(n_903), .A2(n_865), .B(n_869), .C(n_856), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_884), .B(n_876), .C(n_871), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_904), .B(n_838), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_893), .A2(n_836), .B1(n_878), .B2(n_880), .C(n_853), .Y(n_919) );
NAND3x1_ASAP7_75t_L g920 ( .A(n_892), .B(n_883), .C(n_852), .Y(n_920) );
NAND3xp33_ASAP7_75t_SL g921 ( .A(n_905), .B(n_866), .C(n_879), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_895), .B(n_867), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g923 ( .A1(n_887), .A2(n_760), .B(n_870), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_902), .B(n_801), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_898), .B(n_783), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_885), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_918), .Y(n_927) );
AOI211xp5_ASAP7_75t_L g928 ( .A1(n_912), .A2(n_911), .B(n_910), .C(n_906), .Y(n_928) );
NOR3xp33_ASAP7_75t_L g929 ( .A(n_914), .B(n_908), .C(n_896), .Y(n_929) );
NOR4xp25_ASAP7_75t_L g930 ( .A(n_921), .B(n_890), .C(n_907), .D(n_909), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_922), .B(n_897), .Y(n_931) );
NAND4xp25_ASAP7_75t_L g932 ( .A(n_916), .B(n_900), .C(n_885), .D(n_886), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_923), .B(n_888), .Y(n_933) );
NAND2xp33_ASAP7_75t_SL g934 ( .A(n_913), .B(n_920), .Y(n_934) );
AOI211xp5_ASAP7_75t_SL g935 ( .A1(n_928), .A2(n_915), .B(n_917), .C(n_919), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_927), .Y(n_936) );
NOR4xp25_ASAP7_75t_SL g937 ( .A(n_934), .B(n_926), .C(n_916), .D(n_924), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_929), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_929), .B(n_925), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_936), .Y(n_940) );
INVx1_ASAP7_75t_SL g941 ( .A(n_938), .Y(n_941) );
INVxp67_ASAP7_75t_SL g942 ( .A(n_938), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_940), .B(n_935), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_941), .B(n_932), .Y(n_944) );
NAND2xp5_ASAP7_75t_SL g945 ( .A(n_943), .B(n_941), .Y(n_945) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_944), .B(n_942), .Y(n_946) );
INVx3_ASAP7_75t_SL g947 ( .A(n_945), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_946), .Y(n_948) );
NOR4xp75_ASAP7_75t_L g949 ( .A(n_947), .B(n_939), .C(n_937), .D(n_933), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_948), .A2(n_930), .B(n_931), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_949), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_951), .Y(n_952) );
AOI21xp33_ASAP7_75t_L g953 ( .A1(n_952), .A2(n_950), .B(n_886), .Y(n_953) );
OR2x6_ASAP7_75t_L g954 ( .A(n_953), .B(n_894), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_954), .A2(n_891), .B1(n_788), .B2(n_792), .Y(n_955) );
endmodule