module fake_ibex_66_n_5642 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_961, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_5642);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_5642;

wire n_4557;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_968;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_5591;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_5033;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_4757;
wire n_5254;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_5099;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_5157;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5472;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_5403;
wire n_985;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_4682;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_4733;
wire n_5368;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_4412;
wire n_4266;
wire n_5605;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_5506;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_4926;
wire n_5043;
wire n_4688;
wire n_5097;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5221;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4997;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3788;
wire n_3448;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_5294;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5514;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_5193;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_5153;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_5096;
wire n_3712;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_5217;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_3296;
wire n_2671;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_5450;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_5208;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_5245;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_5184;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_5464;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4975;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_3802;
wire n_5343;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_3097;
wire n_2906;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_2564;
wire n_5110;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_4604;
wire n_5123;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_1003;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_2224;
wire n_5526;
wire n_2233;
wire n_2499;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_5435;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_1523;
wire n_1086;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_994;
wire n_5136;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_5634;
wire n_3028;
wire n_3228;
wire n_5079;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_1839;
wire n_5160;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_5313;
wire n_2108;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_2315;
wire n_3623;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5223;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_1105;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_5293;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_5248;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5533;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_5412;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_5479;
wire n_5598;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_5211;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_5279;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_5613;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_5331;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5077;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5105;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_5481;
wire n_5187;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_5485;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5091;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_5306;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_5409;
wire n_2581;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5118;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_2491;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_4147;
wire n_3992;
wire n_4811;
wire n_5093;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_4544;
wire n_4595;
wire n_4418;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_1791;
wire n_5301;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_5507;
wire n_1164;
wire n_3749;
wire n_5470;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_4978;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g968 ( 
.A(n_89),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_684),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_179),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_526),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_777),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_733),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_338),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_745),
.B(n_332),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_158),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_711),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_232),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_357),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_449),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_881),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_131),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_375),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_843),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_685),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_586),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_529),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_136),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_847),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_711),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_559),
.Y(n_991)
);

BUFx10_ASAP7_75t_L g992 ( 
.A(n_936),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_189),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_857),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_912),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_739),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_568),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_622),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_97),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_133),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_365),
.Y(n_1001)
);

BUFx8_ASAP7_75t_SL g1002 ( 
.A(n_940),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_787),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_241),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_386),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_186),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_938),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_98),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_900),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_396),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_939),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_354),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_427),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_13),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_822),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_318),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_439),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_815),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_218),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_319),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_360),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_864),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_899),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_482),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_934),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_913),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_768),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_853),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_906),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_308),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_930),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_277),
.Y(n_1032)
);

BUFx10_ASAP7_75t_L g1033 ( 
.A(n_608),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_301),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_220),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_808),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_287),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_814),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_763),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_330),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_612),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_784),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_956),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_688),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_620),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_619),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_492),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_828),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_850),
.Y(n_1049)
);

BUFx2_ASAP7_75t_R g1050 ( 
.A(n_834),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_769),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_100),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_373),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_209),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_896),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_477),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_336),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_561),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_19),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_430),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_493),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_159),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_540),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_151),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_276),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_331),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_919),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_202),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_592),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_870),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_160),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_347),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_448),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_613),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_861),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_493),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_21),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_392),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_876),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_512),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_326),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_929),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_840),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_95),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_805),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_358),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_791),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_690),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_95),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_143),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_118),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_955),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_64),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_301),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_763),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_159),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_435),
.Y(n_1097)
);

CKINVDCx14_ASAP7_75t_R g1098 ( 
.A(n_911),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_577),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_887),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_490),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_824),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_415),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_136),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_272),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_716),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_28),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_861),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_425),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_411),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_667),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_665),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_868),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_687),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_80),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_863),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_4),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_713),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_230),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_841),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_827),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_195),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_874),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_17),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_227),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_126),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_39),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_897),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_600),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_965),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_261),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_232),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_349),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_57),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_716),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_773),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_875),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_300),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_813),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_419),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_920),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_671),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_305),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_48),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_816),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_745),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_4),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_846),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_162),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_817),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_472),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_145),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_910),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_942),
.Y(n_1154)
);

CKINVDCx14_ASAP7_75t_R g1155 ( 
.A(n_873),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_139),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_537),
.Y(n_1157)
);

BUFx10_ASAP7_75t_L g1158 ( 
.A(n_534),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_578),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_817),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_346),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_298),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_343),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_928),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_740),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_8),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_756),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_663),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_546),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_638),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_806),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_663),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_850),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_829),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_874),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_872),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_921),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_392),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_895),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_199),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_764),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_867),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_394),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_245),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_140),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_534),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_186),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_929),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_615),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_860),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_607),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_81),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_640),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_328),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_835),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_852),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_950),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_778),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_488),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_450),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_576),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_966),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_730),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_231),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_290),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_136),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_922),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_115),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_597),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_221),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_142),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_931),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_127),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_462),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_441),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_775),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_877),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_820),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_377),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_242),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_364),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_925),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_794),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_673),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_880),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_156),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_923),
.Y(n_1227)
);

BUFx5_ASAP7_75t_L g1228 ( 
.A(n_933),
.Y(n_1228)
);

BUFx5_ASAP7_75t_L g1229 ( 
.A(n_321),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_885),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_467),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_893),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_413),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_864),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_72),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_275),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_230),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_24),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_915),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_108),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_644),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_325),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_706),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_652),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_935),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_315),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_424),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_441),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_442),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_286),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_237),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_322),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_155),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_190),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_396),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_278),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_314),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_841),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_803),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_649),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_923),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_253),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_600),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_818),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_236),
.Y(n_1265)
);

CKINVDCx16_ASAP7_75t_R g1266 ( 
.A(n_856),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_714),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_572),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_844),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_744),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_836),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_19),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_804),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_317),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_800),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_405),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_557),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_589),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_520),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_865),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_649),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_241),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_781),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_878),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_34),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_908),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_914),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_927),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_471),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_42),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_887),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_143),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_907),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_336),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_758),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_57),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_890),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_545),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_106),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_505),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_700),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_585),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_958),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_299),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_903),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_886),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_773),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_267),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_918),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_838),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_465),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_926),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_384),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_706),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_98),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_902),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_805),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_75),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_917),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_739),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_638),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_220),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_758),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_94),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_163),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_140),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_661),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_30),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_14),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_514),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_298),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_418),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_832),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_108),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_78),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_835),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_546),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_325),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_670),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_845),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_839),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_552),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_160),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_221),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_32),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_274),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_256),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_92),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_813),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_671),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_6),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_830),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_812),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_319),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_66),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_541),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_809),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_668),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_862),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_603),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_264),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_858),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_477),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_807),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_515),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_496),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_516),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_453),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_683),
.Y(n_1369)
);

CKINVDCx16_ASAP7_75t_R g1370 ( 
.A(n_434),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_800),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_46),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_718),
.Y(n_1373)
);

CKINVDCx14_ASAP7_75t_R g1374 ( 
.A(n_551),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_727),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_455),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_798),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_582),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_155),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_631),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_891),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_790),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_833),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_871),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_447),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_886),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_527),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_845),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_97),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_210),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_562),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_884),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_883),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_271),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_654),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_519),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_522),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_494),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_912),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_854),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_606),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_310),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_635),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_295),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_963),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_361),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_473),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_129),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_30),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_119),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_346),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_937),
.Y(n_1412)
);

INVxp33_ASAP7_75t_L g1413 ( 
.A(n_532),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_126),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_412),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_892),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_811),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_859),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_919),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_592),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_705),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_553),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_11),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_466),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_888),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_482),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_675),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_950),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_965),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_66),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_65),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_690),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_942),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_793),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_244),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_162),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_755),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_642),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_578),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_826),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_119),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_574),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_171),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_869),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_707),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_416),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_391),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_94),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_222),
.Y(n_1449)
);

BUFx2_ASAP7_75t_SL g1450 ( 
.A(n_589),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_692),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_894),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_138),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_132),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_680),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_295),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_163),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_400),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_751),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_566),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_448),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_275),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_960),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_684),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_413),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_130),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_898),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_879),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_868),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_614),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_576),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_832),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_803),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_367),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_837),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_629),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_849),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_767),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_634),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_88),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_823),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_412),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_831),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_157),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_265),
.Y(n_1485)
);

CKINVDCx14_ASAP7_75t_R g1486 ( 
.A(n_208),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_910),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_702),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_378),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_809),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_622),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_906),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_866),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_932),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_86),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_252),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_567),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_513),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_515),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_385),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_476),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_688),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_427),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_133),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_787),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_83),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_246),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_885),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_901),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_836),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_54),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_606),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_39),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_30),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_461),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_291),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_819),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_675),
.Y(n_1518)
);

CKINVDCx16_ASAP7_75t_R g1519 ( 
.A(n_777),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_917),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_660),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_905),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_909),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_521),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_464),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_810),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_741),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_582),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_623),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_729),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_821),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_78),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_251),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_916),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_904),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_492),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_855),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_6),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_289),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_79),
.Y(n_1540)
);

CKINVDCx16_ASAP7_75t_R g1541 ( 
.A(n_882),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_517),
.Y(n_1542)
);

BUFx10_ASAP7_75t_L g1543 ( 
.A(n_842),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_889),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_960),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_373),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_788),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_625),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_16),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_924),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_323),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_494),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_78),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_254),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_495),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_825),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_823),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_898),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_235),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_384),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_422),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_342),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_669),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_48),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_712),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_848),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_588),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_125),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_662),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_665),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_198),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_399),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_58),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_736),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_620),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_212),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_851),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_458),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_90),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_530),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1345),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1313),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1313),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_999),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1413),
.B(n_0),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1345),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1144),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1098),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1423),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1098),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1568),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1573),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_968),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1008),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1059),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1084),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1089),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1091),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1423),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1155),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1117),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1124),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1155),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1134),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1185),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1240),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1285),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1315),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1324),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1334),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1351),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1486),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1052),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1052),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1409),
.Y(n_1616)
);

CKINVDCx16_ASAP7_75t_R g1617 ( 
.A(n_1022),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1414),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1448),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1156),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1506),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1065),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1486),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1374),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1538),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1211),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1211),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1023),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1296),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1504),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1504),
.Y(n_1631)
);

INVxp33_ASAP7_75t_SL g1632 ( 
.A(n_1145),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1576),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1002),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1576),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_998),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_998),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1045),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1045),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_982),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_988),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1080),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1080),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1100),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1100),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1118),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1552),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1118),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1196),
.Y(n_1649)
);

INVxp33_ASAP7_75t_L g1650 ( 
.A(n_1031),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1064),
.B(n_0),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_L g1652 ( 
.A(n_1020),
.B(n_0),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1196),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1204),
.Y(n_1654)
);

INVxp33_ASAP7_75t_SL g1655 ( 
.A(n_1000),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1204),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1389),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1511),
.Y(n_1658)
);

INVxp33_ASAP7_75t_SL g1659 ( 
.A(n_1014),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1298),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1298),
.Y(n_1661)
);

INVxp33_ASAP7_75t_SL g1662 ( 
.A(n_1077),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1093),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1346),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1346),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1553),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1479),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1266),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1479),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1502),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1348),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1502),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1023),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1023),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1534),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1534),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1104),
.Y(n_1677)
);

CKINVDCx14_ASAP7_75t_R g1678 ( 
.A(n_1342),
.Y(n_1678)
);

BUFx2_ASAP7_75t_SL g1679 ( 
.A(n_1023),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1569),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1023),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1367),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1569),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_972),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_972),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1567),
.Y(n_1686)
);

BUFx10_ASAP7_75t_L g1687 ( 
.A(n_1054),
.Y(n_1687)
);

BUFx10_ASAP7_75t_L g1688 ( 
.A(n_1055),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1023),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_994),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1120),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1107),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_994),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_997),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_997),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1025),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1025),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1027),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1027),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1135),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1228),
.Y(n_1701)
);

INVxp33_ASAP7_75t_SL g1702 ( 
.A(n_1115),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1135),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1228),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1175),
.Y(n_1705)
);

INVxp33_ASAP7_75t_SL g1706 ( 
.A(n_1126),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1175),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1243),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1243),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1348),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1260),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1357),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1678),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1701),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1650),
.B(n_1478),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1655),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1687),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1604),
.B(n_1119),
.Y(n_1718)
);

BUFx12f_ASAP7_75t_L g1719 ( 
.A(n_1634),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1581),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1712),
.B(n_1248),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1640),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1641),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1584),
.B(n_1006),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1704),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1691),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1691),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1712),
.B(n_1370),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1659),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1632),
.A2(n_1127),
.B1(n_1166),
.B2(n_1147),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1587),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1589),
.B(n_1048),
.Y(n_1732)
);

AND2x6_ASAP7_75t_L g1733 ( 
.A(n_1651),
.B(n_1348),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1581),
.Y(n_1734)
);

AND2x6_ASAP7_75t_L g1735 ( 
.A(n_1592),
.B(n_1348),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1662),
.A2(n_1206),
.B1(n_1208),
.B2(n_1192),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1586),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1628),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1593),
.B(n_1308),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1590),
.B(n_1213),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1702),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1663),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1687),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1688),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1673),
.A2(n_1287),
.B(n_1260),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1677),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1691),
.Y(n_1747)
);

INVx5_ASAP7_75t_L g1748 ( 
.A(n_1688),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1674),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1600),
.B(n_1235),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1614),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1706),
.B(n_1424),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1622),
.B(n_1519),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1681),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1615),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1689),
.Y(n_1756)
);

CKINVDCx11_ASAP7_75t_R g1757 ( 
.A(n_1596),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1594),
.A2(n_1307),
.B(n_1287),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1582),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1626),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1583),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1595),
.A2(n_1402),
.B(n_1307),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1627),
.Y(n_1763)
);

AND2x2_ASAP7_75t_SL g1764 ( 
.A(n_1617),
.B(n_1541),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1630),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1692),
.A2(n_1272),
.B1(n_1290),
.B2(n_1238),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1588),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1647),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1633),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1624),
.B(n_1299),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1636),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1631),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1638),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1680),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1639),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_L g1776 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1591),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1601),
.A2(n_1623),
.B1(n_1613),
.B2(n_1602),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1642),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1643),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1644),
.Y(n_1781)
);

INVx5_ASAP7_75t_L g1782 ( 
.A(n_1679),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1620),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1645),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1599),
.B(n_1228),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1683),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1684),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1635),
.B(n_1318),
.Y(n_1788)
);

INVxp33_ASAP7_75t_SL g1789 ( 
.A(n_1585),
.Y(n_1789)
);

INVx6_ASAP7_75t_L g1790 ( 
.A(n_1652),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1685),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1637),
.B(n_1653),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1665),
.B(n_1326),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1646),
.Y(n_1794)
);

INVxp67_ASAP7_75t_SL g1795 ( 
.A(n_1669),
.Y(n_1795)
);

INVx4_ASAP7_75t_L g1796 ( 
.A(n_1603),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1605),
.B(n_1328),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1690),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1648),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1649),
.B(n_1406),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1654),
.B(n_1422),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1606),
.B(n_1228),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1656),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1693),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1660),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1661),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1629),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1664),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1667),
.Y(n_1809)
);

OAI21x1_ASAP7_75t_L g1810 ( 
.A1(n_1607),
.A2(n_1520),
.B(n_1402),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1670),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1608),
.A2(n_1610),
.B(n_1609),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1672),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1675),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1676),
.B(n_1555),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1611),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1694),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1695),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1657),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1612),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1616),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1618),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1619),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1621),
.B(n_1329),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1696),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1625),
.Y(n_1826)
);

INVx6_ASAP7_75t_L g1827 ( 
.A(n_1697),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1698),
.B(n_1562),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1699),
.B(n_1700),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1703),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1658),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1666),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1705),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1707),
.B(n_1513),
.Y(n_1834)
);

BUFx8_ASAP7_75t_L g1835 ( 
.A(n_1708),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1709),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1711),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1671),
.B(n_1335),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_L g1839 ( 
.A(n_1668),
.B(n_1228),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1671),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1710),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1710),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1682),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1686),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1701),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1691),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1604),
.B(n_1520),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1581),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1581),
.Y(n_1849)
);

AOI22x1_ASAP7_75t_SL g1850 ( 
.A1(n_1596),
.A2(n_983),
.B1(n_984),
.B2(n_979),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1604),
.B(n_1355),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1701),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1701),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1632),
.A2(n_1408),
.B1(n_1410),
.B2(n_1372),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1701),
.Y(n_1855)
);

INVx5_ASAP7_75t_L g1856 ( 
.A(n_1687),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1604),
.B(n_1523),
.Y(n_1857)
);

AND2x6_ASAP7_75t_L g1858 ( 
.A(n_1651),
.B(n_1120),
.Y(n_1858)
);

OA21x2_ASAP7_75t_L g1859 ( 
.A1(n_1628),
.A2(n_1548),
.B(n_1523),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1628),
.A2(n_1559),
.B(n_1548),
.Y(n_1860)
);

BUFx12f_ASAP7_75t_L g1861 ( 
.A(n_1634),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1701),
.Y(n_1862)
);

AND2x2_ASAP7_75t_SL g1863 ( 
.A(n_1617),
.B(n_1559),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1691),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1581),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1701),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1604),
.B(n_1428),
.Y(n_1867)
);

INVx4_ASAP7_75t_L g1868 ( 
.A(n_1604),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1655),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1604),
.B(n_969),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1581),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1604),
.B(n_1430),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1691),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1687),
.Y(n_1874)
);

BUFx12f_ASAP7_75t_L g1875 ( 
.A(n_1634),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1604),
.B(n_971),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1701),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1712),
.A2(n_1441),
.B1(n_1453),
.B2(n_1431),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1701),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1701),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1678),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1701),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1604),
.Y(n_1883)
);

OA22x2_ASAP7_75t_SL g1884 ( 
.A1(n_1596),
.A2(n_1050),
.B1(n_1009),
.B2(n_1049),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1604),
.B(n_977),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1701),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1650),
.B(n_1466),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1655),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1701),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1650),
.B(n_1480),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1701),
.Y(n_1891)
);

AND2x6_ASAP7_75t_L g1892 ( 
.A(n_1651),
.B(n_1120),
.Y(n_1892)
);

AND2x6_ASAP7_75t_L g1893 ( 
.A(n_1651),
.B(n_1120),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1581),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1655),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1701),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1701),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1650),
.B(n_1495),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1581),
.B(n_1514),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1581),
.Y(n_1900)
);

AOI22x1_ASAP7_75t_SL g1901 ( 
.A1(n_1596),
.A2(n_1073),
.B1(n_1075),
.B2(n_989),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1691),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1691),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1632),
.A2(n_1540),
.B1(n_1549),
.B2(n_1532),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1581),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1581),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1581),
.Y(n_1907)
);

OA21x2_ASAP7_75t_L g1908 ( 
.A1(n_1628),
.A2(n_1004),
.B(n_986),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1701),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1701),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1701),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1687),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1701),
.Y(n_1913)
);

INVx5_ASAP7_75t_L g1914 ( 
.A(n_1687),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1701),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1678),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1581),
.Y(n_1917)
);

AND2x6_ASAP7_75t_L g1918 ( 
.A(n_1651),
.B(n_1165),
.Y(n_1918)
);

INVxp33_ASAP7_75t_SL g1919 ( 
.A(n_1640),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1604),
.B(n_1010),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1687),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1701),
.Y(n_1922)
);

INVx5_ASAP7_75t_L g1923 ( 
.A(n_1687),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1701),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1701),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1628),
.A2(n_1013),
.B(n_1011),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1604),
.B(n_1028),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1678),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1581),
.B(n_1579),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1581),
.B(n_1454),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1581),
.B(n_970),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1691),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1691),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1701),
.Y(n_1934)
);

OA21x2_ASAP7_75t_L g1935 ( 
.A1(n_1628),
.A2(n_1034),
.B(n_1029),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1701),
.Y(n_1936)
);

INVxp33_ASAP7_75t_SL g1937 ( 
.A(n_1640),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1812),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1842),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1812),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1745),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1821),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1859),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1824),
.B(n_1040),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1731),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1860),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1840),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1760),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_L g1949 ( 
.A1(n_1758),
.A2(n_1047),
.B(n_1042),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1758),
.A2(n_1056),
.B(n_1053),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1760),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1774),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1810),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1782),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1751),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1755),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1748),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1757),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1827),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1771),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1773),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1829),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1783),
.A2(n_1198),
.B1(n_1200),
.B2(n_1088),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1829),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1782),
.B(n_1165),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1774),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1810),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1761),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1717),
.B(n_973),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1775),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1784),
.Y(n_1971)
);

BUFx8_ASAP7_75t_L g1972 ( 
.A(n_1807),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1786),
.Y(n_1973)
);

OA21x2_ASAP7_75t_L g1974 ( 
.A1(n_1926),
.A2(n_1061),
.B(n_1057),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1796),
.B(n_1228),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1762),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1794),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1786),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1816),
.B(n_1165),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1787),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1799),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1803),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1805),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1806),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1787),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1811),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1791),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1824),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1791),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1830),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1768),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1833),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1763),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1765),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1713),
.B(n_1207),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1926),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1772),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1744),
.B(n_974),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1816),
.B(n_1229),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1899),
.B(n_1229),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1798),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1887),
.B(n_1890),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1789),
.A2(n_980),
.B1(n_981),
.B2(n_978),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1798),
.Y(n_2004)
);

INVx3_ASAP7_75t_L g2005 ( 
.A(n_1804),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1716),
.B(n_985),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1898),
.B(n_992),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1804),
.Y(n_2008)
);

OR2x6_ASAP7_75t_L g2009 ( 
.A(n_1719),
.B(n_1239),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1818),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1818),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1825),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1825),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1748),
.B(n_1856),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1874),
.B(n_987),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1836),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1836),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1769),
.Y(n_2018)
);

BUFx6f_ASAP7_75t_L g2019 ( 
.A(n_1743),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1779),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1841),
.Y(n_2021)
);

BUFx8_ASAP7_75t_L g2022 ( 
.A(n_1832),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1881),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1817),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1808),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1813),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1837),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1814),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1930),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1856),
.Y(n_2030)
);

BUFx12f_ASAP7_75t_L g2031 ( 
.A(n_1835),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1759),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1737),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1834),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1780),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1715),
.B(n_992),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1908),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1929),
.B(n_1229),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1781),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1916),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1809),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1928),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1753),
.B(n_1033),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1935),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1838),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1795),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_1883),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1776),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1753),
.B(n_1033),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1792),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1722),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1914),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1720),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_1723),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1734),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1728),
.B(n_1051),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1848),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1778),
.B(n_1870),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1914),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1754),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1849),
.B(n_1229),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1865),
.B(n_1229),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1871),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1894),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_1923),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1729),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1754),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1900),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_1741),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1905),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1868),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1820),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1906),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1876),
.B(n_1165),
.Y(n_2074)
);

AOI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1878),
.A2(n_991),
.B1(n_993),
.B2(n_990),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1907),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1917),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1869),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1740),
.B(n_1229),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1923),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1822),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1823),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1851),
.B(n_1051),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1750),
.B(n_995),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1742),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1826),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1746),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1828),
.Y(n_2088)
);

NAND2xp33_ASAP7_75t_L g2089 ( 
.A(n_1733),
.B(n_1270),
.Y(n_2089)
);

INVx6_ASAP7_75t_L g2090 ( 
.A(n_1861),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1800),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1912),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1738),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1888),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1801),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1815),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1749),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1797),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1756),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1785),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1895),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1735),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1735),
.Y(n_2103)
);

AND2x6_ASAP7_75t_L g2104 ( 
.A(n_1851),
.B(n_1872),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1802),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1788),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1793),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1885),
.B(n_1270),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1931),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1921),
.B(n_1062),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1714),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1847),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1857),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1721),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1724),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1725),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1732),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1920),
.B(n_1270),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1852),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1853),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_1718),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1872),
.B(n_1001),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1735),
.Y(n_2123)
);

BUFx6f_ASAP7_75t_L g2124 ( 
.A(n_1733),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1739),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1927),
.B(n_1270),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_1919),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1730),
.B(n_1152),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1855),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1862),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1866),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1877),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1858),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_1770),
.B(n_1069),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1867),
.B(n_1070),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1752),
.B(n_1003),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1790),
.B(n_1005),
.Y(n_2137)
);

CKINVDCx8_ASAP7_75t_R g2138 ( 
.A(n_1831),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1858),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_1736),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1879),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1858),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1733),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1892),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1880),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1882),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1886),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1891),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1766),
.B(n_1854),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_1904),
.B(n_1863),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1845),
.B(n_1889),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1937),
.B(n_1381),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1892),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1892),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1819),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1896),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_1767),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1764),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_1843),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1893),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1893),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1897),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1909),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1893),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1777),
.B(n_1152),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1910),
.B(n_1007),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1911),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_1875),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1918),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1918),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1918),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1843),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1913),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1934),
.B(n_1012),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1915),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_1844),
.Y(n_2176)
);

XNOR2x2_ASAP7_75t_L g2177 ( 
.A(n_1884),
.B(n_975),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1922),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1924),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1925),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1936),
.A2(n_1074),
.B(n_1071),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1839),
.B(n_1158),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1726),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_1726),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1850),
.B(n_1158),
.Y(n_2185)
);

BUFx2_ASAP7_75t_L g2186 ( 
.A(n_1901),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1933),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1933),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1727),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1727),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1747),
.B(n_1015),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1932),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1932),
.Y(n_2193)
);

INVxp67_ASAP7_75t_L g2194 ( 
.A(n_1747),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1846),
.B(n_1016),
.Y(n_2195)
);

BUFx4f_ASAP7_75t_L g2196 ( 
.A(n_1846),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1864),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1864),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1873),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1873),
.Y(n_2200)
);

INVx6_ASAP7_75t_L g2201 ( 
.A(n_1902),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1902),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1903),
.B(n_1017),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1903),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1842),
.Y(n_2205)
);

AND2x6_ASAP7_75t_L g2206 ( 
.A(n_1824),
.B(n_1076),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_1768),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1842),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1812),
.Y(n_2209)
);

OA21x2_ASAP7_75t_L g2210 ( 
.A1(n_1758),
.A2(n_1086),
.B(n_1079),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1812),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1812),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1812),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1812),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_1731),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_1824),
.A2(n_1019),
.B1(n_1021),
.B2(n_1018),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1768),
.B(n_1182),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1796),
.B(n_1024),
.Y(n_2218)
);

CKINVDCx20_ASAP7_75t_R g2219 ( 
.A(n_1757),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1812),
.Y(n_2220)
);

NAND2xp33_ASAP7_75t_SL g2221 ( 
.A(n_1716),
.B(n_1026),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1782),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1812),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1812),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1796),
.B(n_1030),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1768),
.B(n_1182),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1842),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1812),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1842),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1796),
.B(n_1032),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1782),
.B(n_1381),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_SL g2232 ( 
.A1(n_1783),
.A2(n_1230),
.B1(n_1241),
.B2(n_1227),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1812),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1812),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1796),
.B(n_1035),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1812),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1824),
.B(n_1097),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1737),
.A2(n_1037),
.B1(n_1038),
.B2(n_1036),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1842),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1812),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1812),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1955),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1956),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1947),
.Y(n_2244)
);

INVx4_ASAP7_75t_L g2245 ( 
.A(n_1954),
.Y(n_2245)
);

INVx4_ASAP7_75t_L g2246 ( 
.A(n_1954),
.Y(n_2246)
);

AND2x6_ASAP7_75t_L g2247 ( 
.A(n_2098),
.B(n_1102),
.Y(n_2247)
);

NAND2x1p5_ASAP7_75t_L g2248 ( 
.A(n_2014),
.B(n_976),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_1991),
.B(n_1246),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_SL g2250 ( 
.A1(n_1938),
.A2(n_975),
.B(n_1103),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2029),
.A2(n_1570),
.B1(n_1276),
.B2(n_1300),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2106),
.B(n_1039),
.Y(n_2252)
);

NAND2xp33_ASAP7_75t_L g2253 ( 
.A(n_2241),
.B(n_1041),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2107),
.B(n_1043),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_2085),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1939),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2205),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_L g2258 ( 
.A1(n_2140),
.A2(n_1450),
.B1(n_1108),
.B2(n_1109),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2045),
.B(n_1044),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2109),
.B(n_1046),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_2030),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2208),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2030),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2207),
.B(n_1253),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2115),
.B(n_1058),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2014),
.B(n_1320),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2043),
.B(n_1321),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2051),
.B(n_1333),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2227),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2054),
.B(n_1433),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2229),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2239),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2047),
.B(n_1460),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2049),
.B(n_1472),
.Y(n_2274)
);

INVx2_ASAP7_75t_SL g2275 ( 
.A(n_2085),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2127),
.B(n_996),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2056),
.B(n_1483),
.Y(n_2277)
);

INVx4_ASAP7_75t_L g2278 ( 
.A(n_2052),
.Y(n_2278)
);

NAND2xp33_ASAP7_75t_L g2279 ( 
.A(n_2241),
.B(n_1060),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2021),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2181),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2052),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2149),
.B(n_1491),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1945),
.B(n_1063),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_2083),
.B(n_1496),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2059),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2059),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2215),
.B(n_1066),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2117),
.B(n_1067),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_2087),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1958),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2033),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_2040),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2125),
.B(n_1068),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1988),
.B(n_1072),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2157),
.B(n_2087),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_2065),
.Y(n_2297)
);

AND2x2_ASAP7_75t_SL g2298 ( 
.A(n_2040),
.B(n_1106),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2140),
.A2(n_1111),
.B1(n_1113),
.B2(n_1110),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2206),
.A2(n_1129),
.B1(n_1131),
.B2(n_1121),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2042),
.B(n_1083),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2081),
.Y(n_2302)
);

INVx4_ASAP7_75t_L g2303 ( 
.A(n_2065),
.Y(n_2303)
);

BUFx3_ASAP7_75t_L g2304 ( 
.A(n_2168),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2032),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_2042),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_2002),
.B(n_1078),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2019),
.B(n_1081),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1976),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2219),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2018),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2020),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_2080),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2025),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2019),
.B(n_1140),
.Y(n_2315)
);

BUFx8_ASAP7_75t_SL g2316 ( 
.A(n_2031),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1949),
.Y(n_2317)
);

INVx4_ASAP7_75t_L g2318 ( 
.A(n_2080),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1950),
.Y(n_2319)
);

INVxp67_ASAP7_75t_SL g2320 ( 
.A(n_1996),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2026),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2072),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2028),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2071),
.B(n_1173),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2036),
.B(n_1082),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2082),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2222),
.Y(n_2327)
);

INVx3_ASAP7_75t_L g2328 ( 
.A(n_2090),
.Y(n_2328)
);

AND2x6_ASAP7_75t_L g2329 ( 
.A(n_2124),
.B(n_1132),
.Y(n_2329)
);

OAI21xp33_ASAP7_75t_SL g2330 ( 
.A1(n_1940),
.A2(n_1138),
.B(n_1133),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2034),
.B(n_1379),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2086),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2206),
.A2(n_1146),
.B1(n_1154),
.B2(n_1142),
.Y(n_2333)
);

INVx1_ASAP7_75t_SL g2334 ( 
.A(n_2023),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_1972),
.Y(n_2335)
);

INVx2_ASAP7_75t_SL g2336 ( 
.A(n_2172),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1962),
.B(n_1085),
.Y(n_2337)
);

INVx4_ASAP7_75t_L g2338 ( 
.A(n_2090),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1964),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2022),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1996),
.B(n_1087),
.Y(n_2341)
);

CKINVDCx20_ASAP7_75t_R g2342 ( 
.A(n_2066),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2217),
.B(n_1090),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2226),
.B(n_1092),
.Y(n_2344)
);

AOI22xp33_ASAP7_75t_SL g2345 ( 
.A1(n_2104),
.A2(n_2206),
.B1(n_2232),
.B2(n_1963),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2037),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2046),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1968),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2007),
.B(n_1094),
.Y(n_2349)
);

AND2x6_ASAP7_75t_L g2350 ( 
.A(n_2124),
.B(n_1157),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2143),
.B(n_1095),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2104),
.A2(n_1167),
.B1(n_1168),
.B2(n_1162),
.Y(n_2352)
);

INVx6_ASAP7_75t_L g2353 ( 
.A(n_2009),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2165),
.B(n_1096),
.Y(n_2354)
);

BUFx2_ASAP7_75t_L g2355 ( 
.A(n_2104),
.Y(n_2355)
);

INVxp67_ASAP7_75t_L g2356 ( 
.A(n_2155),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1970),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1971),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1977),
.Y(n_2359)
);

INVx5_ASAP7_75t_L g2360 ( 
.A(n_2009),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2143),
.B(n_1099),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1981),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1944),
.B(n_1101),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2069),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2153),
.B(n_1105),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1982),
.Y(n_2366)
);

XOR2xp5_ASAP7_75t_L g2367 ( 
.A(n_2078),
.B(n_1112),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2153),
.B(n_2161),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2159),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1983),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1984),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1986),
.Y(n_2372)
);

BUFx8_ASAP7_75t_SL g2373 ( 
.A(n_2186),
.Y(n_2373)
);

INVx5_ASAP7_75t_L g2374 ( 
.A(n_1957),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2044),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2111),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2092),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_2110),
.Y(n_2378)
);

AND2x6_ASAP7_75t_L g2379 ( 
.A(n_2161),
.B(n_1170),
.Y(n_2379)
);

OR2x2_ASAP7_75t_L g2380 ( 
.A(n_2094),
.B(n_1197),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2116),
.Y(n_2381)
);

NAND2xp33_ASAP7_75t_L g2382 ( 
.A(n_1967),
.B(n_1114),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1993),
.Y(n_2383)
);

AND3x2_ASAP7_75t_L g2384 ( 
.A(n_2186),
.B(n_1178),
.C(n_1176),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1994),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_1944),
.A2(n_2237),
.B1(n_2150),
.B2(n_2134),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2169),
.B(n_1116),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2121),
.B(n_2058),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2119),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2122),
.B(n_1122),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2120),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2110),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_2114),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1997),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2101),
.B(n_1242),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2138),
.Y(n_2396)
);

BUFx10_ASAP7_75t_L g2397 ( 
.A(n_1995),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2024),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2135),
.B(n_1123),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2129),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2237),
.B(n_1379),
.Y(n_2401)
);

AND2x2_ASAP7_75t_SL g2402 ( 
.A(n_2185),
.B(n_2128),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2027),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2135),
.B(n_1125),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2053),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2055),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2057),
.Y(n_2407)
);

INVxp67_ASAP7_75t_SL g2408 ( 
.A(n_1967),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2134),
.B(n_1446),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2136),
.B(n_1128),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2196),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2063),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_2112),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2130),
.Y(n_2414)
);

INVx5_ASAP7_75t_L g2415 ( 
.A(n_2113),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2064),
.Y(n_2416)
);

INVx4_ASAP7_75t_SL g2417 ( 
.A(n_2169),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2068),
.A2(n_1181),
.B1(n_1183),
.B2(n_1179),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2084),
.B(n_1130),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2070),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2131),
.Y(n_2421)
);

INVx4_ASAP7_75t_SL g2422 ( 
.A(n_2050),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2003),
.B(n_1136),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2216),
.B(n_1446),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2132),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2073),
.B(n_1137),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2158),
.B(n_1139),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2075),
.B(n_1543),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_1959),
.Y(n_2429)
);

BUFx10_ASAP7_75t_L g2430 ( 
.A(n_1969),
.Y(n_2430)
);

OR2x6_ASAP7_75t_L g2431 ( 
.A(n_2176),
.B(n_1187),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2076),
.B(n_1141),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_1998),
.B(n_1143),
.Y(n_2433)
);

BUFx4f_ASAP7_75t_L g2434 ( 
.A(n_2091),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2077),
.Y(n_2435)
);

AND2x6_ASAP7_75t_L g2436 ( 
.A(n_2133),
.B(n_1190),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_1942),
.B(n_1148),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_1990),
.B(n_1992),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2182),
.B(n_1149),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_2102),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2015),
.B(n_2095),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2048),
.A2(n_1201),
.B1(n_1203),
.B2(n_1191),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_1960),
.Y(n_2443)
);

CKINVDCx20_ASAP7_75t_R g2444 ( 
.A(n_2006),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2141),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1975),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2238),
.B(n_1543),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2096),
.B(n_1150),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_1961),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2061),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_2102),
.Y(n_2451)
);

INVx4_ASAP7_75t_L g2452 ( 
.A(n_2103),
.Y(n_2452)
);

BUFx2_ASAP7_75t_L g2453 ( 
.A(n_2221),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2035),
.B(n_1151),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2088),
.B(n_1153),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2062),
.Y(n_2456)
);

OR2x6_ASAP7_75t_L g2457 ( 
.A(n_2152),
.B(n_1209),
.Y(n_2457)
);

NOR3xp33_ASAP7_75t_L g2458 ( 
.A(n_2074),
.B(n_1577),
.C(n_1558),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2218),
.Y(n_2459)
);

CKINVDCx20_ASAP7_75t_R g2460 ( 
.A(n_2225),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2230),
.B(n_1159),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2173),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2177),
.Y(n_2463)
);

AND2x6_ASAP7_75t_L g2464 ( 
.A(n_2139),
.B(n_1212),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2039),
.B(n_1160),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2175),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2235),
.B(n_2137),
.Y(n_2467)
);

BUFx3_ASAP7_75t_L g2468 ( 
.A(n_1952),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2041),
.B(n_1161),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2178),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2108),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2118),
.B(n_2126),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2151),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2079),
.B(n_1163),
.Y(n_2474)
);

AND2x6_ASAP7_75t_L g2475 ( 
.A(n_2142),
.B(n_1215),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2103),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2180),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2166),
.B(n_1164),
.Y(n_2478)
);

BUFx2_ASAP7_75t_L g2479 ( 
.A(n_2174),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_1966),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2093),
.B(n_1169),
.Y(n_2481)
);

AOI22xp33_ASAP7_75t_L g2482 ( 
.A1(n_2097),
.A2(n_2099),
.B1(n_2211),
.B2(n_2209),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2145),
.Y(n_2483)
);

INVx3_ASAP7_75t_L g2484 ( 
.A(n_1973),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2146),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2147),
.B(n_1244),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2000),
.B(n_1171),
.Y(n_2487)
);

INVx1_ASAP7_75t_SL g2488 ( 
.A(n_2191),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_1978),
.Y(n_2489)
);

AND3x2_ASAP7_75t_L g2490 ( 
.A(n_2212),
.B(n_1224),
.C(n_1217),
.Y(n_2490)
);

INVxp33_ASAP7_75t_L g2491 ( 
.A(n_2195),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2123),
.B(n_1172),
.Y(n_2492)
);

AOI22xp33_ASAP7_75t_L g2493 ( 
.A1(n_2213),
.A2(n_1237),
.B1(n_1249),
.B2(n_1232),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2148),
.B(n_2156),
.Y(n_2494)
);

INVx5_ASAP7_75t_L g2495 ( 
.A(n_2123),
.Y(n_2495)
);

AND2x6_ASAP7_75t_L g2496 ( 
.A(n_2144),
.B(n_2154),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2162),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2214),
.B(n_1174),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2004),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_1974),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2005),
.Y(n_2501)
);

BUFx6f_ASAP7_75t_L g2502 ( 
.A(n_2184),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2163),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2038),
.B(n_1177),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2167),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2010),
.Y(n_2506)
);

OR2x2_ASAP7_75t_L g2507 ( 
.A(n_2203),
.B(n_1322),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2179),
.B(n_1180),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_1941),
.Y(n_2509)
);

INVxp67_ASAP7_75t_L g2510 ( 
.A(n_1974),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_1943),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2220),
.B(n_1184),
.Y(n_2512)
);

BUFx3_ASAP7_75t_L g2513 ( 
.A(n_2001),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1999),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_1948),
.Y(n_2515)
);

NAND2xp33_ASAP7_75t_L g2516 ( 
.A(n_2223),
.B(n_1186),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_1951),
.Y(n_2517)
);

BUFx10_ASAP7_75t_L g2518 ( 
.A(n_2160),
.Y(n_2518)
);

INVx4_ASAP7_75t_L g2519 ( 
.A(n_2184),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_L g2520 ( 
.A1(n_2224),
.A2(n_1252),
.B1(n_1257),
.B2(n_1250),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2228),
.B(n_1188),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_1953),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2210),
.B(n_1331),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2100),
.B(n_1189),
.Y(n_2524)
);

BUFx10_ASAP7_75t_L g2525 ( 
.A(n_2164),
.Y(n_2525)
);

INVx3_ASAP7_75t_L g2526 ( 
.A(n_1980),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2233),
.B(n_1193),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2234),
.B(n_1194),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1965),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2210),
.B(n_1467),
.Y(n_2530)
);

AOI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2240),
.A2(n_2236),
.B1(n_2170),
.B2(n_2171),
.Y(n_2531)
);

INVx1_ASAP7_75t_SL g2532 ( 
.A(n_2011),
.Y(n_2532)
);

INVx8_ASAP7_75t_L g2533 ( 
.A(n_2231),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_1946),
.Y(n_2534)
);

INVx6_ASAP7_75t_L g2535 ( 
.A(n_2201),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2105),
.B(n_1195),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_1985),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2012),
.B(n_1199),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_L g2539 ( 
.A(n_2201),
.Y(n_2539)
);

AOI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_1987),
.A2(n_1205),
.B1(n_1210),
.B2(n_1202),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_1989),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2008),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2013),
.B(n_1468),
.Y(n_2543)
);

INVx6_ASAP7_75t_L g2544 ( 
.A(n_2194),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2016),
.B(n_1500),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2017),
.Y(n_2546)
);

AND3x2_ASAP7_75t_L g2547 ( 
.A(n_2060),
.B(n_1261),
.C(n_1259),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_1979),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2067),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2089),
.Y(n_2550)
);

INVxp67_ASAP7_75t_SL g2551 ( 
.A(n_2183),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2189),
.B(n_1214),
.Y(n_2552)
);

INVx5_ASAP7_75t_L g2553 ( 
.A(n_2187),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2197),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2198),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_2188),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2199),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_SL g2558 ( 
.A(n_2200),
.B(n_1216),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2204),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2190),
.B(n_1218),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2202),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2192),
.B(n_1219),
.Y(n_2562)
);

INVx3_ASAP7_75t_L g2563 ( 
.A(n_2193),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1955),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_1991),
.B(n_1220),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_1991),
.B(n_1221),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_1991),
.B(n_1222),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_1955),
.Y(n_2568)
);

OR2x6_ASAP7_75t_L g2569 ( 
.A(n_2031),
.B(n_1263),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_1939),
.Y(n_2570)
);

XNOR2xp5_ASAP7_75t_L g2571 ( 
.A(n_2023),
.B(n_1),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_1991),
.B(n_1223),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_1991),
.B(n_1225),
.Y(n_2573)
);

BUFx10_ASAP7_75t_L g2574 ( 
.A(n_2090),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2029),
.B(n_1226),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_1954),
.Y(n_2576)
);

OR2x6_ASAP7_75t_L g2577 ( 
.A(n_2031),
.B(n_1267),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2029),
.B(n_1231),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_1939),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2127),
.B(n_1233),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1955),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2127),
.B(n_1234),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1955),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_1955),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1955),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2029),
.B(n_1236),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2014),
.B(n_1268),
.Y(n_2587)
);

INVx5_ASAP7_75t_L g2588 ( 
.A(n_2031),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2085),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_1991),
.B(n_1245),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2014),
.B(n_1269),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_1954),
.Y(n_2592)
);

OR2x6_ASAP7_75t_L g2593 ( 
.A(n_2031),
.B(n_1271),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2029),
.A2(n_1277),
.B1(n_1278),
.B2(n_1274),
.Y(n_2594)
);

BUFx4f_ASAP7_75t_L g2595 ( 
.A(n_2031),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1955),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_1955),
.Y(n_2597)
);

NOR2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2031),
.B(n_1574),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2047),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2127),
.B(n_1247),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2029),
.B(n_1251),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_1939),
.Y(n_2602)
);

INVx4_ASAP7_75t_L g2603 ( 
.A(n_1954),
.Y(n_2603)
);

AND3x1_ASAP7_75t_L g2604 ( 
.A(n_2185),
.B(n_1280),
.C(n_1279),
.Y(n_2604)
);

NAND2xp33_ASAP7_75t_L g2605 ( 
.A(n_2241),
.B(n_1254),
.Y(n_2605)
);

INVx3_ASAP7_75t_L g2606 ( 
.A(n_1954),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2029),
.B(n_1255),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_1939),
.Y(n_2608)
);

OAI22xp33_ASAP7_75t_SL g2609 ( 
.A1(n_2140),
.A2(n_1258),
.B1(n_1262),
.B2(n_1256),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_1939),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_1939),
.Y(n_2611)
);

BUFx6f_ASAP7_75t_L g2612 ( 
.A(n_1954),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_1955),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1955),
.Y(n_2614)
);

INVxp33_ASAP7_75t_L g2615 ( 
.A(n_2047),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_1939),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2029),
.A2(n_1289),
.B1(n_1292),
.B2(n_1284),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_1954),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_1939),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2029),
.B(n_1264),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_1991),
.B(n_1265),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_1955),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2283),
.B(n_1273),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2247),
.B(n_1275),
.Y(n_2624)
);

INVx1_ASAP7_75t_SL g2625 ( 
.A(n_2599),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2277),
.B(n_1281),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2386),
.A2(n_1283),
.B1(n_1286),
.B2(n_1282),
.Y(n_2627)
);

INVxp67_ASAP7_75t_L g2628 ( 
.A(n_2431),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2247),
.B(n_1288),
.Y(n_2629)
);

NOR2xp33_ASAP7_75t_L g2630 ( 
.A(n_2267),
.B(n_1291),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2274),
.B(n_2285),
.Y(n_2631)
);

OR2x6_ASAP7_75t_L g2632 ( 
.A(n_2353),
.B(n_1301),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2347),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2250),
.A2(n_2441),
.B(n_2330),
.C(n_2450),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2242),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2247),
.B(n_1293),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2243),
.B(n_1294),
.Y(n_2637)
);

OR2x2_ASAP7_75t_L g2638 ( 
.A(n_2251),
.B(n_1295),
.Y(n_2638)
);

OR2x2_ASAP7_75t_L g2639 ( 
.A(n_2364),
.B(n_2334),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2292),
.B(n_1297),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2298),
.A2(n_1303),
.B1(n_1304),
.B2(n_1302),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2369),
.B(n_1554),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2564),
.B(n_2568),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2306),
.B(n_2356),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2309),
.Y(n_2645)
);

OAI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2431),
.A2(n_1306),
.B1(n_1309),
.B2(n_1305),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2581),
.B(n_1310),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_2293),
.B(n_1311),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2615),
.A2(n_1314),
.B1(n_1316),
.B2(n_1312),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2249),
.B(n_1323),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2346),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2332),
.A2(n_1327),
.B1(n_1336),
.B2(n_1325),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2375),
.Y(n_2653)
);

OAI221xp5_ASAP7_75t_L g2654 ( 
.A1(n_2299),
.A2(n_2258),
.B1(n_2345),
.B2(n_2352),
.C(n_2617),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2583),
.B(n_2584),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2585),
.B(n_2596),
.Y(n_2656)
);

OR2x6_ASAP7_75t_L g2657 ( 
.A(n_2353),
.B(n_1317),
.Y(n_2657)
);

AO221x1_ASAP7_75t_L g2658 ( 
.A1(n_2355),
.A2(n_1444),
.B1(n_1525),
.B2(n_1421),
.C(n_1381),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2597),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2613),
.B(n_1337),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2502),
.B(n_2263),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2614),
.B(n_2622),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2302),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2305),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2405),
.B(n_2406),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2273),
.B(n_1338),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2407),
.B(n_1341),
.Y(n_2667)
);

INVx2_ASAP7_75t_SL g2668 ( 
.A(n_2574),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2264),
.B(n_1343),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2412),
.B(n_1347),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2463),
.A2(n_1350),
.B1(n_1352),
.B2(n_1349),
.Y(n_2671)
);

AO221x1_ASAP7_75t_L g2672 ( 
.A1(n_2453),
.A2(n_1444),
.B1(n_1525),
.B2(n_1421),
.C(n_1381),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2416),
.B(n_1353),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2244),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2502),
.B(n_1571),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2420),
.B(n_1354),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2423),
.A2(n_1358),
.B1(n_1360),
.B2(n_1356),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2311),
.Y(n_2678)
);

AOI221xp5_ASAP7_75t_L g2679 ( 
.A1(n_2594),
.A2(n_1332),
.B1(n_1339),
.B2(n_1330),
.C(n_1319),
.Y(n_2679)
);

INVx2_ASAP7_75t_SL g2680 ( 
.A(n_2588),
.Y(n_2680)
);

BUFx3_ASAP7_75t_L g2681 ( 
.A(n_2588),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2435),
.B(n_2312),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2268),
.B(n_1362),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2314),
.B(n_1364),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2270),
.B(n_1365),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2424),
.A2(n_1368),
.B1(n_1369),
.B2(n_1366),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2509),
.A2(n_1373),
.B1(n_1375),
.B2(n_1371),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2321),
.B(n_1376),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2323),
.Y(n_2689)
);

NAND2xp33_ASAP7_75t_L g2690 ( 
.A(n_2440),
.B(n_1580),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2263),
.B(n_2286),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2339),
.B(n_1377),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_R g2693 ( 
.A(n_2340),
.B(n_1378),
.Y(n_2693)
);

A2O1A1Ixp33_ASAP7_75t_L g2694 ( 
.A1(n_2456),
.A2(n_1344),
.B(n_1359),
.C(n_1340),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2252),
.B(n_1380),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2566),
.B(n_2567),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2322),
.Y(n_2697)
);

INVx4_ASAP7_75t_L g2698 ( 
.A(n_2286),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2326),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2254),
.B(n_1382),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2313),
.B(n_1556),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2348),
.Y(n_2702)
);

A2O1A1Ixp33_ASAP7_75t_L g2703 ( 
.A1(n_2446),
.A2(n_1363),
.B(n_1384),
.C(n_1361),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2511),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2534),
.Y(n_2705)
);

NOR2xp67_ASAP7_75t_SL g2706 ( 
.A(n_2360),
.B(n_1566),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2313),
.B(n_1383),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2280),
.Y(n_2708)
);

INVx2_ASAP7_75t_SL g2709 ( 
.A(n_2595),
.Y(n_2709)
);

AO22x2_ASAP7_75t_L g2710 ( 
.A1(n_2367),
.A2(n_1387),
.B1(n_1388),
.B2(n_1385),
.Y(n_2710)
);

AO22x2_ASAP7_75t_L g2711 ( 
.A1(n_2510),
.A2(n_1395),
.B1(n_1398),
.B2(n_1390),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2259),
.B(n_1386),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2467),
.B(n_1391),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2460),
.A2(n_1393),
.B1(n_1394),
.B2(n_1392),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2260),
.B(n_1396),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2281),
.Y(n_2716)
);

AOI22xp33_ASAP7_75t_L g2717 ( 
.A1(n_2409),
.A2(n_2428),
.B1(n_2402),
.B2(n_2307),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2357),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2358),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2388),
.B(n_1397),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2359),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2362),
.Y(n_2722)
);

AOI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2300),
.A2(n_1400),
.B1(n_1401),
.B2(n_1399),
.Y(n_2723)
);

INVxp67_ASAP7_75t_L g2724 ( 
.A(n_2276),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2256),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2366),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2612),
.Y(n_2727)
);

NAND3xp33_ASAP7_75t_L g2728 ( 
.A(n_2433),
.B(n_1444),
.C(n_1421),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2459),
.B(n_2578),
.Y(n_2729)
);

BUFx8_ASAP7_75t_L g2730 ( 
.A(n_2335),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2262),
.Y(n_2731)
);

OAI221xp5_ASAP7_75t_L g2732 ( 
.A1(n_2333),
.A2(n_1405),
.B1(n_1411),
.B2(n_1407),
.C(n_1403),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2370),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_2301),
.B(n_1415),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2272),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2601),
.B(n_2607),
.Y(n_2736)
);

NOR2xp67_ASAP7_75t_L g2737 ( 
.A(n_2495),
.B(n_1),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_SL g2738 ( 
.A(n_2558),
.B(n_1560),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2620),
.B(n_1418),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2371),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2600),
.B(n_1419),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2570),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2372),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2331),
.B(n_1420),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2493),
.B(n_1426),
.Y(n_2745)
);

AOI22xp33_ASAP7_75t_L g2746 ( 
.A1(n_2401),
.A2(n_1432),
.B1(n_1437),
.B2(n_1429),
.Y(n_2746)
);

INVx2_ASAP7_75t_SL g2747 ( 
.A(n_2360),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2520),
.B(n_1438),
.Y(n_2748)
);

NOR3xp33_ASAP7_75t_L g2749 ( 
.A(n_2609),
.B(n_1563),
.C(n_1561),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2579),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2304),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2572),
.B(n_2621),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2383),
.B(n_1442),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2385),
.B(n_1445),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2248),
.B(n_1447),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2602),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2399),
.A2(n_1451),
.B1(n_1452),
.B2(n_1449),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2394),
.B(n_1455),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2600),
.B(n_2580),
.Y(n_2759)
);

INVxp67_ASAP7_75t_L g2760 ( 
.A(n_2380),
.Y(n_2760)
);

AND3x1_ASAP7_75t_L g2761 ( 
.A(n_2396),
.B(n_1412),
.C(n_1404),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2486),
.B(n_2488),
.Y(n_2762)
);

OR2x6_ASAP7_75t_L g2763 ( 
.A(n_2338),
.B(n_1416),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2337),
.B(n_1456),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2404),
.A2(n_1462),
.B1(n_1463),
.B2(n_1457),
.Y(n_2765)
);

O2A1O1Ixp5_ASAP7_75t_L g2766 ( 
.A1(n_2341),
.A2(n_1425),
.B(n_1427),
.C(n_1417),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2479),
.B(n_1465),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2612),
.B(n_1575),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2434),
.B(n_1578),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2447),
.A2(n_1470),
.B1(n_1474),
.B2(n_1469),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2390),
.B(n_1475),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2342),
.Y(n_2772)
);

OAI21xp33_ASAP7_75t_L g2773 ( 
.A1(n_2325),
.A2(n_1481),
.B(n_1476),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2462),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2265),
.B(n_1482),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2378),
.B(n_1544),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2608),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2587),
.A2(n_1485),
.B1(n_1488),
.B2(n_1484),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2466),
.Y(n_2779)
);

INVxp67_ASAP7_75t_L g2780 ( 
.A(n_2395),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2470),
.Y(n_2781)
);

BUFx2_ASAP7_75t_L g2782 ( 
.A(n_2266),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2477),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2398),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2392),
.B(n_1489),
.Y(n_2785)
);

INVxp67_ASAP7_75t_L g2786 ( 
.A(n_2582),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2289),
.B(n_1494),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2294),
.B(n_1498),
.Y(n_2788)
);

NAND3xp33_ASAP7_75t_L g2789 ( 
.A(n_2410),
.B(n_1444),
.C(n_1421),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2403),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2257),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2269),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2440),
.Y(n_2793)
);

NOR3xp33_ASAP7_75t_L g2794 ( 
.A(n_2349),
.B(n_1435),
.C(n_1434),
.Y(n_2794)
);

INVxp67_ASAP7_75t_SL g2795 ( 
.A(n_2522),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2271),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2295),
.B(n_2426),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2565),
.B(n_1503),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2324),
.B(n_1535),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2432),
.B(n_1507),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2473),
.B(n_1508),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2610),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2255),
.B(n_1539),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2393),
.B(n_1509),
.Y(n_2804)
);

INVxp67_ASAP7_75t_SL g2805 ( 
.A(n_2522),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2438),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2354),
.B(n_1510),
.Y(n_2807)
);

NOR3xp33_ASAP7_75t_L g2808 ( 
.A(n_2343),
.B(n_2344),
.C(n_2419),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2573),
.B(n_2590),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2611),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2275),
.B(n_1546),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2491),
.B(n_1515),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2616),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2619),
.Y(n_2814)
);

INVx8_ASAP7_75t_L g2815 ( 
.A(n_2569),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2461),
.B(n_1516),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2483),
.Y(n_2817)
);

OAI21xp33_ASAP7_75t_L g2818 ( 
.A1(n_2448),
.A2(n_1518),
.B(n_1517),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2363),
.B(n_1521),
.Y(n_2819)
);

NOR2xp67_ASAP7_75t_L g2820 ( 
.A(n_2495),
.B(n_1),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2439),
.B(n_1522),
.Y(n_2821)
);

OAI221xp5_ASAP7_75t_L g2822 ( 
.A1(n_2442),
.A2(n_2507),
.B1(n_2455),
.B2(n_2458),
.C(n_2575),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2290),
.Y(n_2823)
);

BUFx3_ASAP7_75t_L g2824 ( 
.A(n_2316),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2589),
.B(n_1526),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2376),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2418),
.B(n_1528),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2485),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2505),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2478),
.B(n_1529),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2381),
.Y(n_2831)
);

OR2x6_ASAP7_75t_L g2832 ( 
.A(n_2569),
.B(n_2577),
.Y(n_2832)
);

INVx2_ASAP7_75t_SL g2833 ( 
.A(n_2374),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2389),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2586),
.B(n_2543),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2444),
.B(n_2430),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2391),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2374),
.B(n_1531),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2400),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2414),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2315),
.B(n_1537),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2604),
.A2(n_1550),
.B1(n_1572),
.B2(n_1547),
.Y(n_2842)
);

NAND2xp33_ASAP7_75t_L g2843 ( 
.A(n_2329),
.B(n_1525),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2421),
.Y(n_2844)
);

OR2x6_ASAP7_75t_L g2845 ( 
.A(n_2577),
.B(n_1436),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2425),
.Y(n_2846)
);

HB1xp67_ASAP7_75t_L g2847 ( 
.A(n_2593),
.Y(n_2847)
);

NAND2xp33_ASAP7_75t_L g2848 ( 
.A(n_2329),
.B(n_1525),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2545),
.B(n_1542),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2445),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2310),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2591),
.B(n_1545),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2443),
.B(n_1551),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2540),
.B(n_1439),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2397),
.B(n_1565),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2497),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2449),
.B(n_1440),
.Y(n_2857)
);

BUFx5_ASAP7_75t_L g2858 ( 
.A(n_2496),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2427),
.B(n_1487),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2413),
.B(n_1490),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2527),
.B(n_1492),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2503),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2494),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_SL g2864 ( 
.A(n_2336),
.B(n_1443),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2413),
.B(n_1497),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2592),
.B(n_1499),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2528),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2481),
.B(n_1501),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2524),
.B(n_1505),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2415),
.B(n_2296),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2415),
.B(n_1512),
.Y(n_2871)
);

INVx1_ASAP7_75t_SL g2872 ( 
.A(n_2544),
.Y(n_2872)
);

INVx2_ASAP7_75t_SL g2873 ( 
.A(n_2328),
.Y(n_2873)
);

INVx2_ASAP7_75t_SL g2874 ( 
.A(n_2544),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2523),
.B(n_1458),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2474),
.B(n_2472),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2519),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2469),
.B(n_1527),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2508),
.Y(n_2879)
);

A2O1A1Ixp33_ASAP7_75t_L g2880 ( 
.A1(n_2514),
.A2(n_1461),
.B(n_1464),
.C(n_1459),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2487),
.B(n_2504),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2454),
.B(n_1557),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2465),
.B(n_1471),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2530),
.B(n_1473),
.Y(n_2884)
);

NOR2xp67_ASAP7_75t_L g2885 ( 
.A(n_2451),
.B(n_2),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2437),
.B(n_1477),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2490),
.B(n_1493),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2317),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2452),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2377),
.B(n_2471),
.Y(n_2890)
);

HB1xp67_ASAP7_75t_L g2891 ( 
.A(n_2593),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2560),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2278),
.B(n_1524),
.Y(n_2893)
);

INVxp67_ASAP7_75t_L g2894 ( 
.A(n_2571),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2516),
.B(n_1530),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2457),
.B(n_2498),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2319),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2562),
.Y(n_2898)
);

NAND3xp33_ASAP7_75t_L g2899 ( 
.A(n_2382),
.B(n_2279),
.C(n_2253),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2554),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2457),
.B(n_1533),
.Y(n_2901)
);

INVxp67_ASAP7_75t_SL g2902 ( 
.A(n_2500),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2303),
.B(n_2318),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2329),
.A2(n_1536),
.B1(n_4),
.B2(n_2),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2512),
.B(n_2),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2521),
.B(n_3),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2559),
.Y(n_2907)
);

INVx1_ASAP7_75t_SL g2908 ( 
.A(n_2350),
.Y(n_2908)
);

NOR3xp33_ASAP7_75t_L g2909 ( 
.A(n_2308),
.B(n_6),
.C(n_5),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2536),
.B(n_3),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2422),
.B(n_3),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2245),
.B(n_7),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_SL g2913 ( 
.A(n_2291),
.B(n_5),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2246),
.B(n_7),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2538),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2547),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2529),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2576),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2603),
.B(n_7),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2546),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2429),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2284),
.B(n_5),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2539),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2422),
.B(n_8),
.Y(n_2924)
);

AND2x4_ASAP7_75t_L g2925 ( 
.A(n_2417),
.B(n_8),
.Y(n_2925)
);

INVxp67_ASAP7_75t_L g2926 ( 
.A(n_2350),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2436),
.B(n_9),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2552),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_SL g2929 ( 
.A(n_2417),
.B(n_10),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2539),
.B(n_2261),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2288),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_L g2932 ( 
.A(n_2541),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2436),
.B(n_9),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2327),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2436),
.B(n_9),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2555),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2282),
.B(n_10),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2541),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2287),
.B(n_10),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2464),
.B(n_11),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2549),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2464),
.B(n_11),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2550),
.Y(n_2943)
);

NAND3xp33_ASAP7_75t_L g2944 ( 
.A(n_2605),
.B(n_12),
.C(n_13),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2464),
.B(n_12),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2297),
.B(n_12),
.Y(n_2946)
);

NAND2xp33_ASAP7_75t_L g2947 ( 
.A(n_2350),
.B(n_14),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2606),
.B(n_13),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2561),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2411),
.B(n_15),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2475),
.B(n_14),
.Y(n_2951)
);

INVxp67_ASAP7_75t_L g2952 ( 
.A(n_2379),
.Y(n_2952)
);

INVxp67_ASAP7_75t_L g2953 ( 
.A(n_2379),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2618),
.B(n_16),
.Y(n_2954)
);

BUFx8_ASAP7_75t_L g2955 ( 
.A(n_2379),
.Y(n_2955)
);

BUFx6f_ASAP7_75t_L g2956 ( 
.A(n_2476),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2475),
.B(n_15),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2475),
.B(n_15),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2482),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2532),
.B(n_17),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2518),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2513),
.B(n_19),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_SL g2963 ( 
.A(n_2468),
.B(n_20),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2556),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2351),
.B(n_18),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2533),
.A2(n_2361),
.B1(n_2387),
.B2(n_2365),
.Y(n_2966)
);

INVxp67_ASAP7_75t_L g2967 ( 
.A(n_2480),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2506),
.B(n_18),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2551),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2484),
.B(n_20),
.Y(n_2970)
);

NAND3xp33_ASAP7_75t_L g2971 ( 
.A(n_2531),
.B(n_21),
.C(n_22),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2525),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2548),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2489),
.B(n_22),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2499),
.B(n_23),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2501),
.B(n_23),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2533),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2492),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2598),
.B(n_23),
.Y(n_2979)
);

AND2x6_ASAP7_75t_SL g2980 ( 
.A(n_2373),
.B(n_24),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2384),
.B(n_24),
.Y(n_2981)
);

BUFx5_ASAP7_75t_L g2982 ( 
.A(n_2496),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2496),
.B(n_25),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2535),
.B(n_25),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2535),
.Y(n_2985)
);

NAND2xp33_ASAP7_75t_L g2986 ( 
.A(n_2556),
.B(n_2368),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2553),
.B(n_2557),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2515),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2553),
.B(n_25),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2517),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2526),
.B(n_26),
.Y(n_2991)
);

OR2x6_ASAP7_75t_L g2992 ( 
.A(n_2537),
.B(n_26),
.Y(n_2992)
);

NAND2x1p5_ASAP7_75t_L g2993 ( 
.A(n_2542),
.B(n_2563),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2320),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2408),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2247),
.B(n_26),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2247),
.B(n_27),
.Y(n_2997)
);

INVx2_ASAP7_75t_SL g2998 ( 
.A(n_2574),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2283),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2369),
.B(n_28),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2347),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2369),
.B(n_29),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2309),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2309),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2309),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2347),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2247),
.B(n_27),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_SL g3008 ( 
.A(n_2369),
.B(n_31),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2316),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2347),
.Y(n_3010)
);

BUFx6f_ASAP7_75t_L g3011 ( 
.A(n_2502),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2369),
.B(n_31),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2283),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2247),
.B(n_32),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2247),
.B(n_33),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2309),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2247),
.B(n_33),
.Y(n_3017)
);

INVxp67_ASAP7_75t_L g3018 ( 
.A(n_2599),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2283),
.B(n_33),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_SL g3020 ( 
.A(n_2369),
.B(n_35),
.Y(n_3020)
);

O2A1O1Ixp33_ASAP7_75t_L g3021 ( 
.A1(n_2250),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2309),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2369),
.B(n_35),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2283),
.B(n_34),
.Y(n_3024)
);

CKINVDCx20_ASAP7_75t_R g3025 ( 
.A(n_2316),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2347),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_L g3027 ( 
.A(n_2283),
.B(n_36),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2283),
.B(n_36),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2247),
.B(n_37),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2247),
.B(n_37),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2247),
.B(n_37),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2347),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2247),
.B(n_38),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2347),
.Y(n_3034)
);

HB1xp67_ASAP7_75t_L g3035 ( 
.A(n_2599),
.Y(n_3035)
);

INVx2_ASAP7_75t_SL g3036 ( 
.A(n_2574),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2283),
.B(n_38),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2347),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2588),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2309),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2283),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_3041)
);

BUFx6f_ASAP7_75t_SL g3042 ( 
.A(n_2335),
.Y(n_3042)
);

NOR2xp67_ASAP7_75t_L g3043 ( 
.A(n_2495),
.B(n_40),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2247),
.B(n_40),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2283),
.B(n_41),
.Y(n_3045)
);

OAI221xp5_ASAP7_75t_L g3046 ( 
.A1(n_2283),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2247),
.B(n_41),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2247),
.B(n_42),
.Y(n_3048)
);

OAI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2251),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2283),
.B(n_43),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2369),
.B(n_45),
.Y(n_3051)
);

INVxp67_ASAP7_75t_SL g3052 ( 
.A(n_2251),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2283),
.B(n_44),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2347),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2347),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2283),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2309),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2247),
.B(n_46),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2247),
.B(n_47),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2247),
.B(n_47),
.Y(n_3060)
);

NOR3xp33_ASAP7_75t_L g3061 ( 
.A(n_2283),
.B(n_50),
.C(n_49),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_2251),
.B(n_48),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2369),
.B(n_50),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2369),
.B(n_50),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2347),
.Y(n_3065)
);

NAND2xp33_ASAP7_75t_SL g3066 ( 
.A(n_2444),
.B(n_49),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2502),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2283),
.B(n_49),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2347),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2247),
.B(n_51),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2309),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2247),
.B(n_51),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2369),
.B(n_52),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2369),
.B(n_52),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2347),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2247),
.B(n_51),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2347),
.Y(n_3077)
);

INVx3_ASAP7_75t_L g3078 ( 
.A(n_2502),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2347),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_2574),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2347),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2247),
.B(n_52),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_2369),
.B(n_54),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2309),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2369),
.B(n_54),
.Y(n_3085)
);

NAND2xp33_ASAP7_75t_L g3086 ( 
.A(n_2502),
.B(n_55),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_2574),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2283),
.B(n_53),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2298),
.B(n_53),
.Y(n_3089)
);

NOR2xp33_ASAP7_75t_L g3090 ( 
.A(n_2283),
.B(n_53),
.Y(n_3090)
);

NOR2xp67_ASAP7_75t_SL g3091 ( 
.A(n_2588),
.B(n_55),
.Y(n_3091)
);

INVx4_ASAP7_75t_L g3092 ( 
.A(n_2588),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2283),
.B(n_55),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2247),
.B(n_56),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2347),
.Y(n_3095)
);

INVxp67_ASAP7_75t_L g3096 ( 
.A(n_2599),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2502),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2247),
.B(n_56),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2283),
.B(n_56),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2309),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2309),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2247),
.B(n_57),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2298),
.B(n_58),
.Y(n_3103)
);

NAND2xp33_ASAP7_75t_L g3104 ( 
.A(n_2502),
.B(n_59),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_SL g3105 ( 
.A(n_2595),
.B(n_58),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_SL g3106 ( 
.A(n_2335),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2309),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2347),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2347),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2574),
.Y(n_3110)
);

OR2x6_ASAP7_75t_L g3111 ( 
.A(n_2353),
.B(n_59),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2283),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2247),
.B(n_60),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2347),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_L g3115 ( 
.A1(n_2283),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2247),
.B(n_61),
.Y(n_3116)
);

AND2x6_ASAP7_75t_SL g3117 ( 
.A(n_2569),
.B(n_62),
.Y(n_3117)
);

AOI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2283),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2369),
.B(n_64),
.Y(n_3119)
);

CKINVDCx5p33_ASAP7_75t_R g3120 ( 
.A(n_2316),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2422),
.B(n_63),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_SL g3122 ( 
.A1(n_2345),
.A2(n_66),
.B1(n_67),
.B2(n_65),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2347),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2283),
.B(n_63),
.Y(n_3124)
);

NOR2xp33_ASAP7_75t_L g3125 ( 
.A(n_2283),
.B(n_65),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2298),
.B(n_67),
.Y(n_3126)
);

AOI22xp33_ASAP7_75t_L g3127 ( 
.A1(n_2283),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2347),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2347),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2247),
.B(n_68),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2247),
.B(n_68),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2247),
.B(n_69),
.Y(n_3132)
);

OR2x2_ASAP7_75t_L g3133 ( 
.A(n_2251),
.B(n_69),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2247),
.B(n_70),
.Y(n_3134)
);

A2O1A1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2250),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_2298),
.B(n_70),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2247),
.B(n_71),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2347),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_2251),
.B(n_71),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2283),
.B(n_72),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2247),
.B(n_73),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2283),
.B(n_73),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2247),
.B(n_73),
.Y(n_3143)
);

BUFx3_ASAP7_75t_L g3144 ( 
.A(n_2588),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2283),
.B(n_74),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2247),
.B(n_74),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2369),
.B(n_75),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2369),
.B(n_75),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2283),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2369),
.B(n_77),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2347),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2347),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2369),
.B(n_77),
.Y(n_3153)
);

NOR2x1p5_ASAP7_75t_L g3154 ( 
.A(n_2335),
.B(n_76),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2369),
.B(n_79),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2247),
.B(n_76),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_2283),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2247),
.B(n_80),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2309),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2309),
.Y(n_3160)
);

AO22x2_ASAP7_75t_L g3161 ( 
.A1(n_2251),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2247),
.B(n_82),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2369),
.B(n_83),
.Y(n_3163)
);

AOI22xp5_ASAP7_75t_L g3164 ( 
.A1(n_2283),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2369),
.B(n_85),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2309),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2247),
.B(n_84),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2309),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2283),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_2369),
.B(n_87),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2369),
.B(n_87),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2347),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2309),
.Y(n_3173)
);

INVxp67_ASAP7_75t_L g3174 ( 
.A(n_2599),
.Y(n_3174)
);

INVx2_ASAP7_75t_SL g3175 ( 
.A(n_2574),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2347),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2309),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2309),
.Y(n_3178)
);

CKINVDCx5p33_ASAP7_75t_R g3179 ( 
.A(n_2316),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2283),
.B(n_86),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2247),
.B(n_87),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2247),
.B(n_88),
.Y(n_3182)
);

NOR2xp67_ASAP7_75t_L g3183 ( 
.A(n_2495),
.B(n_88),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2309),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2247),
.B(n_89),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2247),
.B(n_89),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2309),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2347),
.Y(n_3188)
);

AOI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2283),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3189)
);

NOR3xp33_ASAP7_75t_L g3190 ( 
.A(n_2283),
.B(n_92),
.C(n_91),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_SL g3191 ( 
.A(n_2369),
.B(n_91),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2347),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2283),
.B(n_90),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2309),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2369),
.B(n_94),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2283),
.A2(n_96),
.B1(n_93),
.B2(n_95),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2247),
.B(n_93),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_2298),
.B(n_93),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_SL g3199 ( 
.A(n_2595),
.B(n_96),
.Y(n_3199)
);

INVxp67_ASAP7_75t_L g3200 ( 
.A(n_2599),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2247),
.B(n_96),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2247),
.B(n_97),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2347),
.Y(n_3203)
);

BUFx3_ASAP7_75t_L g3204 ( 
.A(n_2588),
.Y(n_3204)
);

AOI22xp33_ASAP7_75t_L g3205 ( 
.A1(n_2283),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2347),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2347),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2369),
.B(n_100),
.Y(n_3208)
);

NOR2x1p5_ASAP7_75t_L g3209 ( 
.A(n_2335),
.B(n_99),
.Y(n_3209)
);

INVxp67_ASAP7_75t_SL g3210 ( 
.A(n_2251),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2247),
.B(n_99),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_2283),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2247),
.B(n_101),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_2369),
.B(n_102),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_2247),
.B(n_101),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2247),
.B(n_102),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2347),
.Y(n_3217)
);

NAND2xp33_ASAP7_75t_L g3218 ( 
.A(n_2502),
.B(n_104),
.Y(n_3218)
);

INVx2_ASAP7_75t_SL g3219 ( 
.A(n_2574),
.Y(n_3219)
);

NAND2x1_ASAP7_75t_L g3220 ( 
.A(n_2502),
.B(n_103),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_2422),
.B(n_103),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2247),
.B(n_104),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2247),
.B(n_104),
.Y(n_3223)
);

NAND3xp33_ASAP7_75t_L g3224 ( 
.A(n_2433),
.B(n_105),
.C(n_106),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2309),
.Y(n_3225)
);

OR2x2_ASAP7_75t_L g3226 ( 
.A(n_2251),
.B(n_105),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2247),
.B(n_105),
.Y(n_3227)
);

NOR2xp67_ASAP7_75t_L g3228 ( 
.A(n_2495),
.B(n_106),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2309),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2247),
.B(n_107),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2369),
.B(n_108),
.Y(n_3231)
);

NAND3xp33_ASAP7_75t_L g3232 ( 
.A(n_2433),
.B(n_107),
.C(n_109),
.Y(n_3232)
);

INVxp67_ASAP7_75t_L g3233 ( 
.A(n_2599),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_L g3234 ( 
.A(n_2283),
.B(n_107),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2386),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2247),
.B(n_109),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2309),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2309),
.Y(n_3238)
);

INVx4_ASAP7_75t_L g3239 ( 
.A(n_2588),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2309),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2247),
.B(n_110),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2369),
.B(n_111),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2247),
.B(n_110),
.Y(n_3243)
);

INVx8_ASAP7_75t_L g3244 ( 
.A(n_2588),
.Y(n_3244)
);

NAND2xp33_ASAP7_75t_L g3245 ( 
.A(n_2502),
.B(n_112),
.Y(n_3245)
);

BUFx5_ASAP7_75t_L g3246 ( 
.A(n_2496),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2283),
.B(n_111),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2347),
.Y(n_3248)
);

INVx2_ASAP7_75t_SL g3249 ( 
.A(n_2574),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2369),
.B(n_113),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_SL g3251 ( 
.A(n_2369),
.B(n_113),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_2316),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_2283),
.B(n_112),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2347),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2283),
.B(n_112),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2247),
.B(n_113),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2247),
.B(n_114),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2247),
.B(n_114),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2247),
.B(n_114),
.Y(n_3259)
);

NOR3xp33_ASAP7_75t_L g3260 ( 
.A(n_2283),
.B(n_117),
.C(n_116),
.Y(n_3260)
);

AOI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_2283),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2247),
.B(n_115),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2309),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2347),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2806),
.B(n_116),
.Y(n_3265)
);

AND2x6_ASAP7_75t_SL g3266 ( 
.A(n_2832),
.B(n_117),
.Y(n_3266)
);

OR2x6_ASAP7_75t_L g3267 ( 
.A(n_3244),
.B(n_118),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2762),
.B(n_2696),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_3244),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2752),
.B(n_118),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2633),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2659),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2674),
.Y(n_3273)
);

NOR2x2_ASAP7_75t_L g3274 ( 
.A(n_2832),
.B(n_120),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2645),
.Y(n_3275)
);

NAND2x1p5_ASAP7_75t_L g3276 ( 
.A(n_3092),
.B(n_119),
.Y(n_3276)
);

AND2x4_ASAP7_75t_L g3277 ( 
.A(n_2867),
.B(n_120),
.Y(n_3277)
);

HB1xp67_ASAP7_75t_L g3278 ( 
.A(n_2625),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2759),
.B(n_120),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3052),
.B(n_121),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3210),
.B(n_121),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_2832),
.Y(n_3282)
);

INVx4_ASAP7_75t_L g3283 ( 
.A(n_3244),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_3035),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3001),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_2631),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_3286)
);

HB1xp67_ASAP7_75t_L g3287 ( 
.A(n_3018),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2736),
.B(n_122),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2634),
.A2(n_122),
.B(n_123),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_2879),
.B(n_123),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3006),
.B(n_3010),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_3011),
.Y(n_3292)
);

NOR2xp67_ASAP7_75t_L g3293 ( 
.A(n_3092),
.B(n_3239),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3089),
.B(n_3103),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_2646),
.B(n_144),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_2730),
.Y(n_3296)
);

INVx6_ASAP7_75t_L g3297 ( 
.A(n_2730),
.Y(n_3297)
);

OR2x2_ASAP7_75t_L g3298 ( 
.A(n_2760),
.B(n_124),
.Y(n_3298)
);

CKINVDCx5p33_ASAP7_75t_R g3299 ( 
.A(n_3025),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_3011),
.Y(n_3300)
);

HB1xp67_ASAP7_75t_L g3301 ( 
.A(n_3096),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2651),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_3011),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2653),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3026),
.Y(n_3305)
);

BUFx4f_ASAP7_75t_L g3306 ( 
.A(n_2815),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_2915),
.B(n_124),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2704),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3032),
.B(n_3034),
.Y(n_3309)
);

NAND3xp33_ASAP7_75t_L g3310 ( 
.A(n_3061),
.B(n_3260),
.C(n_3190),
.Y(n_3310)
);

BUFx8_ASAP7_75t_L g3311 ( 
.A(n_3042),
.Y(n_3311)
);

BUFx3_ASAP7_75t_L g3312 ( 
.A(n_2681),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3038),
.B(n_124),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_2628),
.B(n_125),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3054),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3055),
.B(n_3065),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2705),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3069),
.B(n_125),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3067),
.B(n_144),
.Y(n_3319)
);

BUFx2_ASAP7_75t_L g3320 ( 
.A(n_2845),
.Y(n_3320)
);

AND2x4_ASAP7_75t_L g3321 ( 
.A(n_2698),
.B(n_126),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3075),
.B(n_127),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3077),
.Y(n_3323)
);

HB1xp67_ASAP7_75t_L g3324 ( 
.A(n_3174),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3079),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3081),
.B(n_127),
.Y(n_3326)
);

OR2x2_ASAP7_75t_L g3327 ( 
.A(n_2780),
.B(n_128),
.Y(n_3327)
);

HB1xp67_ASAP7_75t_L g3328 ( 
.A(n_3200),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_2654),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3095),
.B(n_128),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3126),
.B(n_129),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3108),
.B(n_130),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_3067),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3109),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3114),
.B(n_131),
.Y(n_3335)
);

BUFx3_ASAP7_75t_L g3336 ( 
.A(n_3039),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3003),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_2724),
.B(n_131),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_2782),
.B(n_132),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_SL g3340 ( 
.A1(n_2815),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3136),
.B(n_134),
.Y(n_3341)
);

AND2x4_ASAP7_75t_L g3342 ( 
.A(n_2698),
.B(n_134),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_2727),
.B(n_135),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2786),
.B(n_135),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3004),
.Y(n_3345)
);

A2O1A1Ixp33_ASAP7_75t_L g3346 ( 
.A1(n_3021),
.A2(n_138),
.B(n_135),
.C(n_137),
.Y(n_3346)
);

BUFx6f_ASAP7_75t_L g3347 ( 
.A(n_3067),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_2992),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3123),
.B(n_137),
.Y(n_3349)
);

BUFx3_ASAP7_75t_L g3350 ( 
.A(n_3144),
.Y(n_3350)
);

NOR2x2_ASAP7_75t_L g3351 ( 
.A(n_2845),
.B(n_140),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3128),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3129),
.B(n_139),
.Y(n_3353)
);

BUFx6f_ASAP7_75t_L g3354 ( 
.A(n_3097),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3005),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3138),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3151),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3152),
.B(n_3172),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3016),
.Y(n_3359)
);

OAI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_2845),
.A2(n_3111),
.B1(n_2992),
.B2(n_2913),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3176),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3188),
.Y(n_3362)
);

CKINVDCx8_ASAP7_75t_R g3363 ( 
.A(n_2815),
.Y(n_3363)
);

INVxp67_ASAP7_75t_L g3364 ( 
.A(n_2639),
.Y(n_3364)
);

INVx5_ASAP7_75t_L g3365 ( 
.A(n_3239),
.Y(n_3365)
);

BUFx6f_ASAP7_75t_L g3366 ( 
.A(n_3097),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_2992),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_3367)
);

OAI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2797),
.A2(n_2881),
.B(n_2766),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3192),
.Y(n_3369)
);

AOI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_2809),
.A2(n_3019),
.B1(n_3027),
.B2(n_3024),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3028),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_2632),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3097),
.B(n_146),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_2727),
.B(n_141),
.Y(n_3374)
);

BUFx2_ASAP7_75t_L g3375 ( 
.A(n_2632),
.Y(n_3375)
);

XNOR2xp5_ASAP7_75t_L g3376 ( 
.A(n_3154),
.B(n_147),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_2822),
.B(n_147),
.Y(n_3377)
);

AND2x4_ASAP7_75t_L g3378 ( 
.A(n_2892),
.B(n_148),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3203),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3206),
.B(n_3207),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3217),
.B(n_148),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_2894),
.B(n_149),
.Y(n_3382)
);

NOR2x1p5_ASAP7_75t_L g3383 ( 
.A(n_2824),
.B(n_3009),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3248),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_2623),
.B(n_149),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3254),
.B(n_150),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3264),
.Y(n_3387)
);

NAND2x1p5_ASAP7_75t_L g3388 ( 
.A(n_3204),
.B(n_150),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2635),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2729),
.B(n_151),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3037),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_3391)
);

AND2x6_ASAP7_75t_SL g3392 ( 
.A(n_3111),
.B(n_152),
.Y(n_3392)
);

AO21x1_ASAP7_75t_L g3393 ( 
.A1(n_2947),
.A2(n_153),
.B(n_154),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_2716),
.A2(n_156),
.B(n_157),
.Y(n_3394)
);

OR2x2_ASAP7_75t_L g3395 ( 
.A(n_2638),
.B(n_158),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_2842),
.B(n_161),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3022),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2663),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2664),
.B(n_161),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2678),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3040),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_2772),
.B(n_164),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2689),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3045),
.A2(n_3053),
.B1(n_3068),
.B2(n_3050),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_2932),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_2680),
.Y(n_3406)
);

NAND3xp33_ASAP7_75t_L g3407 ( 
.A(n_3088),
.B(n_164),
.C(n_165),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_2842),
.B(n_2847),
.Y(n_3408)
);

INVxp67_ASAP7_75t_SL g3409 ( 
.A(n_2902),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_2891),
.B(n_3233),
.Y(n_3410)
);

AND2x4_ASAP7_75t_L g3411 ( 
.A(n_2898),
.B(n_165),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2702),
.Y(n_3412)
);

BUFx6f_ASAP7_75t_L g3413 ( 
.A(n_2932),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2643),
.B(n_166),
.Y(n_3414)
);

NAND2xp33_ASAP7_75t_L g3415 ( 
.A(n_2858),
.B(n_953),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2718),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_2863),
.B(n_166),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3057),
.Y(n_3418)
);

AOI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_2741),
.A2(n_3090),
.B1(n_3099),
.B2(n_3093),
.Y(n_3419)
);

INVx4_ASAP7_75t_L g3420 ( 
.A(n_3042),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2719),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3124),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3422)
);

NOR2xp33_ASAP7_75t_R g3423 ( 
.A(n_3120),
.B(n_954),
.Y(n_3423)
);

HB1xp67_ASAP7_75t_L g3424 ( 
.A(n_3111),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3071),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2655),
.B(n_167),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_2904),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2721),
.Y(n_3428)
);

AO21x1_ASAP7_75t_L g3429 ( 
.A1(n_2843),
.A2(n_170),
.B(n_171),
.Y(n_3429)
);

CKINVDCx5p33_ASAP7_75t_R g3430 ( 
.A(n_3179),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_2714),
.B(n_172),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3084),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2722),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_2656),
.B(n_172),
.Y(n_3434)
);

HB1xp67_ASAP7_75t_L g3435 ( 
.A(n_2632),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_3125),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_2734),
.B(n_173),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_2657),
.Y(n_3438)
);

BUFx2_ASAP7_75t_L g3439 ( 
.A(n_2657),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2726),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2733),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_2662),
.B(n_174),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2740),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2743),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_3252),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_2657),
.B(n_175),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2665),
.B(n_176),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_SL g3448 ( 
.A1(n_2710),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3448)
);

OAI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3105),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_3449)
);

BUFx2_ASAP7_75t_L g3450 ( 
.A(n_2763),
.Y(n_3450)
);

NOR3xp33_ASAP7_75t_L g3451 ( 
.A(n_3046),
.B(n_3122),
.C(n_3140),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2774),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_3142),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3453)
);

NAND2x1p5_ASAP7_75t_L g3454 ( 
.A(n_2709),
.B(n_180),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_2955),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_L g3456 ( 
.A1(n_3145),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2779),
.Y(n_3457)
);

OAI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_2904),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2682),
.B(n_184),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3100),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_2781),
.B(n_185),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_2763),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2783),
.B(n_187),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3101),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_SL g3465 ( 
.A(n_2851),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3107),
.Y(n_3466)
);

NAND3xp33_ASAP7_75t_SL g3467 ( 
.A(n_3199),
.B(n_187),
.C(n_188),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3180),
.B(n_188),
.Y(n_3468)
);

HB1xp67_ASAP7_75t_L g3469 ( 
.A(n_2763),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3193),
.B(n_189),
.Y(n_3470)
);

BUFx2_ASAP7_75t_L g3471 ( 
.A(n_2955),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_R g3472 ( 
.A(n_3106),
.B(n_961),
.Y(n_3472)
);

HB1xp67_ASAP7_75t_L g3473 ( 
.A(n_2872),
.Y(n_3473)
);

BUFx6f_ASAP7_75t_L g3474 ( 
.A(n_2932),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_2784),
.Y(n_3475)
);

OR2x2_ASAP7_75t_L g3476 ( 
.A(n_2713),
.B(n_190),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3159),
.Y(n_3477)
);

OAI22xp5_ASAP7_75t_SL g3478 ( 
.A1(n_2761),
.A2(n_199),
.B1(n_207),
.B2(n_191),
.Y(n_3478)
);

NAND2x1p5_ASAP7_75t_L g3479 ( 
.A(n_2668),
.B(n_191),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3234),
.B(n_192),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3247),
.B(n_192),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_2790),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_2626),
.B(n_193),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_2908),
.B(n_193),
.Y(n_3484)
);

INVxp67_ASAP7_75t_L g3485 ( 
.A(n_2755),
.Y(n_3485)
);

AO22x1_ASAP7_75t_L g3486 ( 
.A1(n_3121),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3253),
.B(n_3255),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_3066),
.B(n_194),
.Y(n_3488)
);

OR2x6_ASAP7_75t_L g3489 ( 
.A(n_3209),
.B(n_196),
.Y(n_3489)
);

HB1xp67_ASAP7_75t_L g3490 ( 
.A(n_2751),
.Y(n_3490)
);

NOR2xp33_ASAP7_75t_L g3491 ( 
.A(n_2630),
.B(n_197),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_2749),
.A2(n_200),
.B1(n_197),
.B2(n_198),
.Y(n_3492)
);

CKINVDCx5p33_ASAP7_75t_R g3493 ( 
.A(n_3106),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_2817),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3160),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_2833),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3166),
.Y(n_3497)
);

AOI221xp5_ASAP7_75t_SL g3498 ( 
.A1(n_3135),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_3498)
);

AND2x2_ASAP7_75t_SL g3499 ( 
.A(n_2848),
.B(n_201),
.Y(n_3499)
);

INVx1_ASAP7_75t_SL g3500 ( 
.A(n_2693),
.Y(n_3500)
);

CKINVDCx20_ASAP7_75t_R g3501 ( 
.A(n_2998),
.Y(n_3501)
);

HB1xp67_ASAP7_75t_L g3502 ( 
.A(n_2874),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3168),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_2828),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3198),
.B(n_203),
.Y(n_3505)
);

BUFx12f_ASAP7_75t_L g3506 ( 
.A(n_3117),
.Y(n_3506)
);

BUFx3_ASAP7_75t_L g3507 ( 
.A(n_3036),
.Y(n_3507)
);

NOR3xp33_ASAP7_75t_L g3508 ( 
.A(n_2808),
.B(n_204),
.C(n_205),
.Y(n_3508)
);

BUFx2_ASAP7_75t_L g3509 ( 
.A(n_3080),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_3121),
.B(n_204),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_2717),
.B(n_205),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_SL g3512 ( 
.A(n_3221),
.B(n_206),
.Y(n_3512)
);

OR2x2_ASAP7_75t_SL g3513 ( 
.A(n_3062),
.B(n_961),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3173),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2829),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_2791),
.Y(n_3516)
);

INVx5_ASAP7_75t_L g3517 ( 
.A(n_2938),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_2710),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_2792),
.Y(n_3519)
);

AOI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_2888),
.A2(n_209),
.B(n_210),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_2799),
.B(n_211),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2703),
.B(n_211),
.Y(n_3522)
);

NAND3xp33_ASAP7_75t_SL g3523 ( 
.A(n_2999),
.B(n_212),
.C(n_213),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_2859),
.B(n_2694),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2880),
.B(n_213),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2796),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3177),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_2900),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2794),
.B(n_214),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3178),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3184),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_2907),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2697),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3187),
.Y(n_3534)
);

CKINVDCx20_ASAP7_75t_R g3535 ( 
.A(n_3087),
.Y(n_3535)
);

INVx1_ASAP7_75t_SL g3536 ( 
.A(n_2644),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2699),
.Y(n_3537)
);

INVx3_ASAP7_75t_L g3538 ( 
.A(n_2956),
.Y(n_3538)
);

INVx2_ASAP7_75t_SL g3539 ( 
.A(n_2956),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3194),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_2810),
.Y(n_3541)
);

AOI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_2669),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_2896),
.B(n_215),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3221),
.B(n_216),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_2666),
.B(n_217),
.Y(n_3545)
);

INVx3_ASAP7_75t_L g3546 ( 
.A(n_2956),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_2814),
.Y(n_3547)
);

INVx5_ASAP7_75t_L g3548 ( 
.A(n_2938),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_2849),
.B(n_2835),
.Y(n_3549)
);

AND2x4_ASAP7_75t_L g3550 ( 
.A(n_2977),
.B(n_217),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_2834),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_2876),
.B(n_218),
.Y(n_3552)
);

INVx3_ASAP7_75t_L g3553 ( 
.A(n_3110),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2861),
.B(n_219),
.Y(n_3554)
);

OAI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_2711),
.A2(n_223),
.B1(n_219),
.B2(n_222),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_2931),
.B(n_223),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_2938),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_2869),
.B(n_224),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_2878),
.B(n_224),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_2999),
.B(n_225),
.Y(n_3560)
);

OAI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_2711),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3561)
);

BUFx3_ASAP7_75t_L g3562 ( 
.A(n_3175),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2837),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2650),
.B(n_226),
.Y(n_3564)
);

NOR2x1p5_ASAP7_75t_L g3565 ( 
.A(n_3133),
.B(n_228),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3225),
.Y(n_3566)
);

NOR3xp33_ASAP7_75t_SL g3567 ( 
.A(n_2836),
.B(n_228),
.C(n_229),
.Y(n_3567)
);

AND2x6_ASAP7_75t_SL g3568 ( 
.A(n_2979),
.B(n_229),
.Y(n_3568)
);

INVx5_ASAP7_75t_L g3569 ( 
.A(n_2964),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3219),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3139),
.B(n_231),
.Y(n_3571)
);

INVx4_ASAP7_75t_L g3572 ( 
.A(n_2923),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3013),
.B(n_233),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_SL g3574 ( 
.A(n_2925),
.B(n_2737),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3013),
.B(n_233),
.Y(n_3575)
);

HB1xp67_ASAP7_75t_L g3576 ( 
.A(n_3249),
.Y(n_3576)
);

INVx2_ASAP7_75t_SL g3577 ( 
.A(n_2918),
.Y(n_3577)
);

CKINVDCx5p33_ASAP7_75t_R g3578 ( 
.A(n_2980),
.Y(n_3578)
);

AND2x4_ASAP7_75t_L g3579 ( 
.A(n_3078),
.B(n_234),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_2909),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3078),
.B(n_237),
.Y(n_3581)
);

NOR3xp33_ASAP7_75t_SL g3582 ( 
.A(n_3049),
.B(n_238),
.C(n_239),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_2683),
.A2(n_2685),
.B1(n_2807),
.B2(n_2641),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_2798),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_3584)
);

OR2x6_ASAP7_75t_L g3585 ( 
.A(n_2925),
.B(n_240),
.Y(n_3585)
);

INVx3_ASAP7_75t_L g3586 ( 
.A(n_2923),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3118),
.B(n_242),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3226),
.B(n_243),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_2648),
.B(n_243),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3118),
.B(n_244),
.Y(n_3590)
);

OAI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2875),
.A2(n_245),
.B(n_246),
.Y(n_3591)
);

BUFx6f_ASAP7_75t_L g3592 ( 
.A(n_2964),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_2839),
.Y(n_3593)
);

INVx2_ASAP7_75t_SL g3594 ( 
.A(n_2923),
.Y(n_3594)
);

INVx2_ASAP7_75t_SL g3595 ( 
.A(n_2747),
.Y(n_3595)
);

INVx3_ASAP7_75t_L g3596 ( 
.A(n_2877),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_2737),
.B(n_247),
.Y(n_3597)
);

O2A1O1Ixp5_ASAP7_75t_L g3598 ( 
.A1(n_2884),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_2840),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2844),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2846),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_2820),
.B(n_248),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3189),
.B(n_249),
.Y(n_3603)
);

CKINVDCx5p33_ASAP7_75t_R g3604 ( 
.A(n_2981),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_2850),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3189),
.B(n_250),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_2868),
.B(n_250),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_2679),
.B(n_251),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_2856),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3229),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2723),
.B(n_252),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3237),
.Y(n_3612)
);

AOI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_2812),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_2885),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3161),
.Y(n_3615)
);

OR2x2_ASAP7_75t_L g3616 ( 
.A(n_2767),
.B(n_255),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3161),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3238),
.Y(n_3618)
);

BUFx2_ASAP7_75t_L g3619 ( 
.A(n_2967),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_2723),
.B(n_256),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_2820),
.B(n_257),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_2725),
.Y(n_3622)
);

BUFx3_ASAP7_75t_L g3623 ( 
.A(n_2877),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3041),
.B(n_257),
.Y(n_3624)
);

BUFx6f_ASAP7_75t_L g3625 ( 
.A(n_2964),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3043),
.B(n_258),
.Y(n_3626)
);

BUFx10_ASAP7_75t_L g3627 ( 
.A(n_2870),
.Y(n_3627)
);

AOI22xp33_ASAP7_75t_L g3628 ( 
.A1(n_2922),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_2901),
.B(n_259),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_2889),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2731),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_2735),
.Y(n_3632)
);

OAI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3164),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3169),
.B(n_262),
.Y(n_3634)
);

OAI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3224),
.A2(n_263),
.B(n_264),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3196),
.B(n_263),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_SL g3637 ( 
.A1(n_2996),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3043),
.B(n_266),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_2742),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_2854),
.B(n_268),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_2750),
.Y(n_3641)
);

INVx5_ASAP7_75t_L g3642 ( 
.A(n_2793),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3056),
.B(n_268),
.Y(n_3643)
);

NOR2xp67_ASAP7_75t_L g3644 ( 
.A(n_2961),
.B(n_269),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_R g3645 ( 
.A(n_2690),
.B(n_954),
.Y(n_3645)
);

BUFx6f_ASAP7_75t_L g3646 ( 
.A(n_2793),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3112),
.B(n_269),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2756),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_2777),
.Y(n_3649)
);

HB1xp67_ASAP7_75t_L g3650 ( 
.A(n_2885),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3240),
.Y(n_3651)
);

AOI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_2897),
.A2(n_270),
.B(n_271),
.Y(n_3652)
);

AND2x2_ASAP7_75t_SL g3653 ( 
.A(n_3086),
.B(n_270),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3183),
.B(n_272),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_2852),
.B(n_273),
.Y(n_3655)
);

INVx3_ASAP7_75t_L g3656 ( 
.A(n_2889),
.Y(n_3656)
);

BUFx2_ASAP7_75t_L g3657 ( 
.A(n_2823),
.Y(n_3657)
);

INVx1_ASAP7_75t_SL g3658 ( 
.A(n_2825),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3115),
.B(n_273),
.Y(n_3659)
);

INVx4_ASAP7_75t_L g3660 ( 
.A(n_2993),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3127),
.B(n_274),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3183),
.B(n_276),
.Y(n_3662)
);

AOI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_2841),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3663)
);

INVx6_ASAP7_75t_L g3664 ( 
.A(n_2984),
.Y(n_3664)
);

INVx2_ASAP7_75t_SL g3665 ( 
.A(n_2873),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3149),
.B(n_279),
.Y(n_3666)
);

OR2x2_ASAP7_75t_L g3667 ( 
.A(n_2627),
.B(n_280),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3157),
.B(n_280),
.Y(n_3668)
);

AOI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_2855),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3205),
.B(n_281),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3212),
.B(n_3261),
.Y(n_3671)
);

NOR2xp33_ASAP7_75t_L g3672 ( 
.A(n_2642),
.B(n_282),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_2745),
.B(n_283),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_2785),
.B(n_284),
.Y(n_3674)
);

INVx1_ASAP7_75t_SL g3675 ( 
.A(n_2989),
.Y(n_3675)
);

OAI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3232),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3263),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_2708),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_2802),
.Y(n_3679)
);

AND2x4_ASAP7_75t_L g3680 ( 
.A(n_2978),
.B(n_2928),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_2972),
.B(n_285),
.Y(n_3681)
);

AND2x4_ASAP7_75t_L g3682 ( 
.A(n_2990),
.B(n_2988),
.Y(n_3682)
);

AOI22xp5_ASAP7_75t_L g3683 ( 
.A1(n_2686),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_2866),
.B(n_288),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3228),
.B(n_290),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_2813),
.Y(n_3686)
);

INVx2_ASAP7_75t_SL g3687 ( 
.A(n_2903),
.Y(n_3687)
);

CKINVDCx16_ASAP7_75t_R g3688 ( 
.A(n_2652),
.Y(n_3688)
);

INVx4_ASAP7_75t_L g3689 ( 
.A(n_2826),
.Y(n_3689)
);

NOR3xp33_ASAP7_75t_L g3690 ( 
.A(n_3000),
.B(n_291),
.C(n_292),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_2853),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_2831),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2748),
.B(n_292),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_2857),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_2969),
.Y(n_3695)
);

BUFx6f_ASAP7_75t_L g3696 ( 
.A(n_3220),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_SL g3697 ( 
.A(n_3228),
.B(n_293),
.Y(n_3697)
);

AOI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_2986),
.A2(n_293),
.B(n_294),
.Y(n_3698)
);

NOR3xp33_ASAP7_75t_SL g3699 ( 
.A(n_2887),
.B(n_294),
.C(n_296),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_2862),
.Y(n_3700)
);

INVx2_ASAP7_75t_SL g3701 ( 
.A(n_2890),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_2882),
.B(n_296),
.Y(n_3702)
);

BUFx4f_ASAP7_75t_L g3703 ( 
.A(n_2916),
.Y(n_3703)
);

CKINVDCx5p33_ASAP7_75t_R g3704 ( 
.A(n_2985),
.Y(n_3704)
);

BUFx3_ASAP7_75t_L g3705 ( 
.A(n_2934),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_2883),
.B(n_297),
.Y(n_3706)
);

NAND3xp33_ASAP7_75t_SL g3707 ( 
.A(n_2677),
.B(n_297),
.C(n_299),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_2949),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_2886),
.B(n_300),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_2624),
.B(n_302),
.Y(n_3710)
);

AND2x4_ASAP7_75t_L g3711 ( 
.A(n_2921),
.B(n_302),
.Y(n_3711)
);

CKINVDCx20_ASAP7_75t_R g3712 ( 
.A(n_2738),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2692),
.B(n_303),
.Y(n_3713)
);

OR2x6_ASAP7_75t_L g3714 ( 
.A(n_2926),
.B(n_303),
.Y(n_3714)
);

AO21x1_ASAP7_75t_L g3715 ( 
.A1(n_2959),
.A2(n_304),
.B(n_305),
.Y(n_3715)
);

CKINVDCx6p67_ASAP7_75t_R g3716 ( 
.A(n_2838),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3262),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_2695),
.B(n_304),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_2700),
.B(n_306),
.Y(n_3719)
);

BUFx12f_ASAP7_75t_SL g3720 ( 
.A(n_2706),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_2960),
.Y(n_3721)
);

HB1xp67_ASAP7_75t_L g3722 ( 
.A(n_2997),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_2917),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_2936),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_2970),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_R g3726 ( 
.A(n_3104),
.B(n_956),
.Y(n_3726)
);

AND2x4_ASAP7_75t_L g3727 ( 
.A(n_2691),
.B(n_306),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_2712),
.B(n_307),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_2974),
.Y(n_3729)
);

CKINVDCx16_ASAP7_75t_R g3730 ( 
.A(n_3235),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3002),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_2827),
.B(n_309),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_SL g3733 ( 
.A(n_2629),
.B(n_310),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_2636),
.B(n_311),
.Y(n_3734)
);

AOI22xp5_ASAP7_75t_L g3735 ( 
.A1(n_3008),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3735)
);

NOR2x1p5_ASAP7_75t_L g3736 ( 
.A(n_3007),
.B(n_312),
.Y(n_3736)
);

BUFx3_ASAP7_75t_L g3737 ( 
.A(n_2968),
.Y(n_3737)
);

BUFx12f_ASAP7_75t_L g3738 ( 
.A(n_3091),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_2975),
.Y(n_3739)
);

INVx2_ASAP7_75t_SL g3740 ( 
.A(n_2987),
.Y(n_3740)
);

A2O1A1Ixp33_ASAP7_75t_L g3741 ( 
.A1(n_2971),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_2976),
.Y(n_3742)
);

INVxp67_ASAP7_75t_L g3743 ( 
.A(n_3014),
.Y(n_3743)
);

BUFx4f_ASAP7_75t_L g3744 ( 
.A(n_2973),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_2715),
.B(n_316),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_2739),
.B(n_316),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_2770),
.B(n_317),
.Y(n_3747)
);

NAND2xp33_ASAP7_75t_SL g3748 ( 
.A(n_3015),
.B(n_318),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_2920),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_2941),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_2943),
.Y(n_3751)
);

NOR2x2_ASAP7_75t_L g3752 ( 
.A(n_2778),
.B(n_320),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_2773),
.B(n_320),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_2994),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_2775),
.B(n_321),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_2787),
.B(n_322),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_2995),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_2910),
.Y(n_3758)
);

OAI22x1_ASAP7_75t_L g3759 ( 
.A1(n_2929),
.A2(n_326),
.B1(n_327),
.B2(n_324),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_2905),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_2788),
.B(n_323),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_2728),
.A2(n_324),
.B(n_327),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_R g3763 ( 
.A(n_3218),
.B(n_963),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_2819),
.B(n_328),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_2637),
.B(n_329),
.Y(n_3765)
);

OR2x4_ASAP7_75t_L g3766 ( 
.A(n_2965),
.B(n_329),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_2640),
.B(n_330),
.Y(n_3767)
);

NAND2xp33_ASAP7_75t_L g3768 ( 
.A(n_2858),
.B(n_331),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_SL g3769 ( 
.A(n_2952),
.B(n_332),
.Y(n_3769)
);

AND2x6_ASAP7_75t_SL g3770 ( 
.A(n_2860),
.B(n_333),
.Y(n_3770)
);

BUFx4f_ASAP7_75t_L g3771 ( 
.A(n_2769),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_2906),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_2789),
.A2(n_333),
.B(n_334),
.Y(n_3773)
);

INVxp67_ASAP7_75t_L g3774 ( 
.A(n_3017),
.Y(n_3774)
);

AND2x4_ASAP7_75t_L g3775 ( 
.A(n_2661),
.B(n_334),
.Y(n_3775)
);

OAI22xp5_ASAP7_75t_SL g3776 ( 
.A1(n_3029),
.A2(n_344),
.B1(n_353),
.B2(n_335),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_2991),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_2672),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_2744),
.B(n_2816),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_2937),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_2953),
.B(n_2858),
.Y(n_3781)
);

BUFx2_ASAP7_75t_L g3782 ( 
.A(n_3030),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_2658),
.Y(n_3783)
);

NAND2x2_ASAP7_75t_L g3784 ( 
.A(n_2911),
.B(n_335),
.Y(n_3784)
);

AOI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_3012),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_2939),
.Y(n_3786)
);

AOI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3020),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.Y(n_3787)
);

BUFx4f_ASAP7_75t_L g3788 ( 
.A(n_2966),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3023),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_3789)
);

BUFx3_ASAP7_75t_L g3790 ( 
.A(n_2924),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_2983),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3031),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_SL g3793 ( 
.A(n_2858),
.B(n_341),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_2647),
.B(n_343),
.Y(n_3794)
);

HB1xp67_ASAP7_75t_L g3795 ( 
.A(n_3033),
.Y(n_3795)
);

INVx3_ASAP7_75t_L g3796 ( 
.A(n_2858),
.Y(n_3796)
);

OR2x2_ASAP7_75t_L g3797 ( 
.A(n_2801),
.B(n_344),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_SL g3798 ( 
.A(n_2982),
.B(n_345),
.Y(n_3798)
);

AND3x1_ASAP7_75t_L g3799 ( 
.A(n_2821),
.B(n_345),
.C(n_347),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_2660),
.B(n_348),
.Y(n_3800)
);

INVx5_ASAP7_75t_L g3801 ( 
.A(n_3245),
.Y(n_3801)
);

INVxp67_ASAP7_75t_SL g3802 ( 
.A(n_3044),
.Y(n_3802)
);

AOI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3051),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3803)
);

OR2x6_ASAP7_75t_L g3804 ( 
.A(n_2963),
.B(n_350),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_2667),
.B(n_351),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_2946),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_L g3807 ( 
.A1(n_3063),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_3807)
);

INVx2_ASAP7_75t_SL g3808 ( 
.A(n_2675),
.Y(n_3808)
);

OR2x6_ASAP7_75t_L g3809 ( 
.A(n_3047),
.B(n_352),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_2948),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3048),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_2670),
.B(n_2673),
.Y(n_3812)
);

NOR2x1_ASAP7_75t_L g3813 ( 
.A(n_2944),
.B(n_354),
.Y(n_3813)
);

INVx4_ASAP7_75t_L g3814 ( 
.A(n_2982),
.Y(n_3814)
);

OR2x2_ASAP7_75t_L g3815 ( 
.A(n_2687),
.B(n_355),
.Y(n_3815)
);

BUFx3_ASAP7_75t_L g3816 ( 
.A(n_3058),
.Y(n_3816)
);

NAND3xp33_ASAP7_75t_SL g3817 ( 
.A(n_3059),
.B(n_355),
.C(n_356),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3060),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3064),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2676),
.B(n_359),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3070),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_3821)
);

OR2x4_ASAP7_75t_L g3822 ( 
.A(n_2865),
.B(n_362),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3268),
.B(n_3073),
.Y(n_3823)
);

BUFx3_ASAP7_75t_L g3824 ( 
.A(n_3283),
.Y(n_3824)
);

CKINVDCx12_ASAP7_75t_R g3825 ( 
.A(n_3267),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3294),
.B(n_2649),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3272),
.Y(n_3827)
);

BUFx2_ASAP7_75t_L g3828 ( 
.A(n_3744),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3271),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_3297),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3278),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3285),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3305),
.Y(n_3833)
);

NAND2x1p5_ASAP7_75t_L g3834 ( 
.A(n_3306),
.B(n_3365),
.Y(n_3834)
);

AND2x4_ASAP7_75t_SL g3835 ( 
.A(n_3267),
.B(n_2746),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3549),
.B(n_3074),
.Y(n_3836)
);

INVx2_ASAP7_75t_SL g3837 ( 
.A(n_3297),
.Y(n_3837)
);

BUFx2_ASAP7_75t_L g3838 ( 
.A(n_3365),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3779),
.B(n_3083),
.Y(n_3839)
);

BUFx8_ASAP7_75t_L g3840 ( 
.A(n_3465),
.Y(n_3840)
);

BUFx8_ASAP7_75t_L g3841 ( 
.A(n_3471),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3365),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3364),
.B(n_3085),
.Y(n_3843)
);

CKINVDCx5p33_ASAP7_75t_R g3844 ( 
.A(n_3296),
.Y(n_3844)
);

OAI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3310),
.A2(n_3242),
.B(n_3231),
.Y(n_3845)
);

AND2x4_ASAP7_75t_L g3846 ( 
.A(n_3293),
.B(n_2893),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3360),
.B(n_3072),
.Y(n_3847)
);

BUFx3_ASAP7_75t_L g3848 ( 
.A(n_3311),
.Y(n_3848)
);

BUFx6f_ASAP7_75t_L g3849 ( 
.A(n_3292),
.Y(n_3849)
);

BUFx6f_ASAP7_75t_L g3850 ( 
.A(n_3292),
.Y(n_3850)
);

HB1xp67_ASAP7_75t_L g3851 ( 
.A(n_3284),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3315),
.Y(n_3852)
);

BUFx3_ASAP7_75t_L g3853 ( 
.A(n_3311),
.Y(n_3853)
);

O2A1O1Ixp33_ASAP7_75t_L g3854 ( 
.A1(n_3487),
.A2(n_3251),
.B(n_3250),
.C(n_3147),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3323),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3331),
.B(n_3119),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_R g3857 ( 
.A(n_3363),
.B(n_3076),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3451),
.A2(n_3148),
.B1(n_3153),
.B2(n_3150),
.Y(n_3858)
);

INVx3_ASAP7_75t_L g3859 ( 
.A(n_3269),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3370),
.B(n_3155),
.Y(n_3860)
);

BUFx6f_ASAP7_75t_L g3861 ( 
.A(n_3292),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3691),
.B(n_3694),
.Y(n_3862)
);

AND2x4_ASAP7_75t_L g3863 ( 
.A(n_3501),
.B(n_2701),
.Y(n_3863)
);

HB1xp67_ASAP7_75t_L g3864 ( 
.A(n_3435),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3299),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3325),
.Y(n_3866)
);

NOR2xp33_ASAP7_75t_L g3867 ( 
.A(n_3688),
.B(n_2732),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3334),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3352),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3658),
.B(n_3163),
.Y(n_3870)
);

BUFx6f_ASAP7_75t_L g3871 ( 
.A(n_3300),
.Y(n_3871)
);

CKINVDCx6p67_ASAP7_75t_R g3872 ( 
.A(n_3489),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3356),
.Y(n_3873)
);

OR2x2_ASAP7_75t_L g3874 ( 
.A(n_3395),
.B(n_3215),
.Y(n_3874)
);

HB1xp67_ASAP7_75t_L g3875 ( 
.A(n_3462),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3273),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3357),
.B(n_3165),
.Y(n_3877)
);

OAI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3499),
.A2(n_3094),
.B1(n_3098),
.B2(n_3082),
.Y(n_3878)
);

CKINVDCx5p33_ASAP7_75t_R g3879 ( 
.A(n_3430),
.Y(n_3879)
);

CKINVDCx5p33_ASAP7_75t_R g3880 ( 
.A(n_3445),
.Y(n_3880)
);

BUFx12f_ASAP7_75t_L g3881 ( 
.A(n_3493),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3653),
.B(n_3102),
.Y(n_3882)
);

INVx4_ASAP7_75t_L g3883 ( 
.A(n_3312),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3415),
.A2(n_2805),
.B(n_2795),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3361),
.B(n_3170),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3528),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3801),
.B(n_3113),
.Y(n_3887)
);

OR2x6_ASAP7_75t_L g3888 ( 
.A(n_3489),
.B(n_3116),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_SL g3889 ( 
.A(n_3801),
.B(n_3130),
.Y(n_3889)
);

AND3x1_ASAP7_75t_SL g3890 ( 
.A(n_3383),
.B(n_362),
.C(n_363),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3362),
.Y(n_3891)
);

BUFx3_ASAP7_75t_L g3892 ( 
.A(n_3535),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3369),
.B(n_3379),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3384),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3341),
.B(n_3171),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_3801),
.B(n_3131),
.Y(n_3896)
);

BUFx6f_ASAP7_75t_L g3897 ( 
.A(n_3300),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3532),
.Y(n_3898)
);

CKINVDCx5p33_ASAP7_75t_R g3899 ( 
.A(n_3506),
.Y(n_3899)
);

INVx4_ASAP7_75t_L g3900 ( 
.A(n_3336),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3469),
.Y(n_3901)
);

NOR2xp67_ASAP7_75t_L g3902 ( 
.A(n_3282),
.B(n_3132),
.Y(n_3902)
);

HB1xp67_ASAP7_75t_L g3903 ( 
.A(n_3287),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3387),
.B(n_3191),
.Y(n_3904)
);

BUFx3_ASAP7_75t_L g3905 ( 
.A(n_3350),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3533),
.Y(n_3906)
);

AOI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3730),
.A2(n_3195),
.B1(n_3214),
.B2(n_3208),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_3301),
.Y(n_3908)
);

OR2x6_ASAP7_75t_L g3909 ( 
.A(n_3585),
.B(n_3134),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3505),
.B(n_3137),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3507),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3277),
.B(n_3141),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3389),
.B(n_3398),
.Y(n_3913)
);

OR2x6_ASAP7_75t_L g3914 ( 
.A(n_3585),
.B(n_3143),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3562),
.Y(n_3915)
);

BUFx6f_ASAP7_75t_L g3916 ( 
.A(n_3300),
.Y(n_3916)
);

INVx1_ASAP7_75t_SL g3917 ( 
.A(n_3509),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3537),
.Y(n_3918)
);

BUFx6f_ASAP7_75t_L g3919 ( 
.A(n_3303),
.Y(n_3919)
);

INVx3_ASAP7_75t_L g3920 ( 
.A(n_3660),
.Y(n_3920)
);

BUFx6f_ASAP7_75t_L g3921 ( 
.A(n_3303),
.Y(n_3921)
);

AOI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3565),
.A2(n_3146),
.B1(n_3158),
.B2(n_3156),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3400),
.B(n_2684),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3726),
.B(n_3162),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3377),
.A2(n_3181),
.B(n_3182),
.C(n_3167),
.Y(n_3925)
);

HB1xp67_ASAP7_75t_L g3926 ( 
.A(n_3324),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3403),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3541),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3412),
.Y(n_3929)
);

INVxp67_ASAP7_75t_L g3930 ( 
.A(n_3328),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3416),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3763),
.B(n_3185),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3421),
.Y(n_3933)
);

INVx3_ASAP7_75t_L g3934 ( 
.A(n_3406),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_R g3935 ( 
.A(n_3720),
.B(n_3186),
.Y(n_3935)
);

INVx3_ASAP7_75t_L g3936 ( 
.A(n_3623),
.Y(n_3936)
);

A2O1A1Ixp33_ASAP7_75t_L g3937 ( 
.A1(n_3419),
.A2(n_3201),
.B(n_3202),
.C(n_3197),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3547),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3378),
.B(n_3211),
.Y(n_3939)
);

OR2x6_ASAP7_75t_L g3940 ( 
.A(n_3738),
.B(n_3213),
.Y(n_3940)
);

CKINVDCx5p33_ASAP7_75t_R g3941 ( 
.A(n_3578),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_3303),
.Y(n_3942)
);

OAI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_3404),
.A2(n_3222),
.B1(n_3223),
.B2(n_3216),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3428),
.Y(n_3944)
);

HB1xp67_ASAP7_75t_L g3945 ( 
.A(n_3450),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3433),
.B(n_2688),
.Y(n_3946)
);

OAI22xp5_ASAP7_75t_SL g3947 ( 
.A1(n_3376),
.A2(n_3230),
.B1(n_3236),
.B2(n_3227),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3788),
.A2(n_3241),
.B1(n_3256),
.B2(n_3243),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3440),
.B(n_2895),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3378),
.B(n_3257),
.Y(n_3950)
);

INVx4_ASAP7_75t_L g3951 ( 
.A(n_3392),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3333),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3441),
.B(n_3258),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3372),
.Y(n_3954)
);

NOR2xp33_ASAP7_75t_L g3955 ( 
.A(n_3485),
.B(n_3320),
.Y(n_3955)
);

OR2x6_ASAP7_75t_L g3956 ( 
.A(n_3455),
.B(n_3259),
.Y(n_3956)
);

INVx1_ASAP7_75t_SL g3957 ( 
.A(n_3619),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3443),
.B(n_2753),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3551),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3444),
.B(n_2754),
.Y(n_3960)
);

BUFx3_ASAP7_75t_L g3961 ( 
.A(n_3577),
.Y(n_3961)
);

BUFx6f_ASAP7_75t_L g3962 ( 
.A(n_3333),
.Y(n_3962)
);

A2O1A1Ixp33_ASAP7_75t_L g3963 ( 
.A1(n_3385),
.A2(n_2927),
.B(n_2935),
.C(n_2933),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3452),
.B(n_2758),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3457),
.Y(n_3965)
);

BUFx6f_ASAP7_75t_L g3966 ( 
.A(n_3333),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3563),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3695),
.B(n_2871),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3291),
.B(n_2671),
.Y(n_3969)
);

INVx3_ASAP7_75t_L g3970 ( 
.A(n_3689),
.Y(n_3970)
);

AOI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3583),
.A2(n_2962),
.B1(n_2912),
.B2(n_2919),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3475),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3593),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3309),
.B(n_2720),
.Y(n_3974)
);

HB1xp67_ASAP7_75t_L g3975 ( 
.A(n_3375),
.Y(n_3975)
);

NOR3xp33_ASAP7_75t_L g3976 ( 
.A(n_3467),
.B(n_2914),
.C(n_2950),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3438),
.Y(n_3977)
);

INVx3_ASAP7_75t_L g3978 ( 
.A(n_3703),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3316),
.B(n_3358),
.Y(n_3979)
);

INVx2_ASAP7_75t_SL g3980 ( 
.A(n_3539),
.Y(n_3980)
);

OAI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3513),
.A2(n_2940),
.B1(n_2945),
.B2(n_2942),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3439),
.B(n_2776),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3380),
.B(n_2818),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_R g3984 ( 
.A(n_3500),
.B(n_2951),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3482),
.B(n_2757),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3347),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3494),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3504),
.Y(n_3988)
);

NAND2x1p5_ASAP7_75t_L g3989 ( 
.A(n_3420),
.B(n_2707),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3408),
.B(n_2864),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3515),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3516),
.B(n_2765),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3411),
.B(n_2982),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3519),
.B(n_2764),
.Y(n_3994)
);

HB1xp67_ASAP7_75t_L g3995 ( 
.A(n_3657),
.Y(n_3995)
);

NOR2xp33_ASAP7_75t_L g3996 ( 
.A(n_3664),
.B(n_2803),
.Y(n_3996)
);

CKINVDCx8_ASAP7_75t_R g3997 ( 
.A(n_3266),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3526),
.B(n_2800),
.Y(n_3998)
);

OR2x2_ASAP7_75t_L g3999 ( 
.A(n_3277),
.B(n_2957),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3599),
.Y(n_4000)
);

HB1xp67_ASAP7_75t_L g4001 ( 
.A(n_3409),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3600),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3601),
.Y(n_4003)
);

BUFx8_ASAP7_75t_L g4004 ( 
.A(n_3402),
.Y(n_4004)
);

INVx3_ASAP7_75t_L g4005 ( 
.A(n_3716),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3605),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3288),
.B(n_2830),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3664),
.B(n_2811),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3609),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3723),
.Y(n_4010)
);

AOI22xp33_ASAP7_75t_L g4011 ( 
.A1(n_3615),
.A2(n_3617),
.B1(n_3508),
.B2(n_3483),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3812),
.B(n_2954),
.Y(n_4012)
);

BUFx2_ASAP7_75t_L g4013 ( 
.A(n_3538),
.Y(n_4013)
);

BUFx6f_ASAP7_75t_L g4014 ( 
.A(n_3347),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3275),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3724),
.Y(n_4016)
);

AND2x4_ASAP7_75t_L g4017 ( 
.A(n_3570),
.B(n_2768),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3511),
.B(n_2771),
.Y(n_4018)
);

BUFx4f_ASAP7_75t_L g4019 ( 
.A(n_3388),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3302),
.Y(n_4020)
);

OR2x6_ASAP7_75t_L g4021 ( 
.A(n_3276),
.B(n_2958),
.Y(n_4021)
);

BUFx4f_ASAP7_75t_L g4022 ( 
.A(n_3479),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3304),
.Y(n_4023)
);

AOI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3431),
.A2(n_2804),
.B1(n_2899),
.B2(n_2930),
.Y(n_4024)
);

BUFx6f_ASAP7_75t_L g4025 ( 
.A(n_3347),
.Y(n_4025)
);

INVx4_ASAP7_75t_L g4026 ( 
.A(n_3546),
.Y(n_4026)
);

BUFx3_ASAP7_75t_L g4027 ( 
.A(n_3553),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3524),
.B(n_2982),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_SL g4029 ( 
.A(n_3411),
.B(n_2982),
.Y(n_4029)
);

NOR2xp67_ASAP7_75t_L g4030 ( 
.A(n_3496),
.B(n_363),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3279),
.B(n_3246),
.Y(n_4031)
);

INVx3_ASAP7_75t_L g4032 ( 
.A(n_3771),
.Y(n_4032)
);

AOI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3307),
.A2(n_3246),
.B1(n_366),
.B2(n_364),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_L g4034 ( 
.A1(n_3491),
.A2(n_3246),
.B1(n_367),
.B2(n_365),
.Y(n_4034)
);

INVx3_ASAP7_75t_L g4035 ( 
.A(n_3596),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3622),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3777),
.B(n_3246),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3608),
.B(n_3246),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3631),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_SL g4040 ( 
.A(n_3417),
.B(n_366),
.Y(n_4040)
);

BUFx2_ASAP7_75t_L g4041 ( 
.A(n_3572),
.Y(n_4041)
);

BUFx3_ASAP7_75t_L g4042 ( 
.A(n_3576),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3632),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3307),
.B(n_368),
.Y(n_4044)
);

BUFx6f_ASAP7_75t_L g4045 ( 
.A(n_3354),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3308),
.Y(n_4046)
);

BUFx6f_ASAP7_75t_L g4047 ( 
.A(n_3354),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3290),
.B(n_368),
.Y(n_4048)
);

INVx3_ASAP7_75t_L g4049 ( 
.A(n_3656),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3675),
.B(n_369),
.Y(n_4050)
);

BUFx6f_ASAP7_75t_L g4051 ( 
.A(n_3354),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3639),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3760),
.B(n_369),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3758),
.B(n_3571),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3588),
.B(n_370),
.Y(n_4055)
);

HB1xp67_ASAP7_75t_L g4056 ( 
.A(n_3290),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3368),
.B(n_370),
.Y(n_4057)
);

OR2x2_ASAP7_75t_L g4058 ( 
.A(n_3446),
.B(n_371),
.Y(n_4058)
);

CKINVDCx5p33_ASAP7_75t_R g4059 ( 
.A(n_3423),
.Y(n_4059)
);

INVx3_ASAP7_75t_L g4060 ( 
.A(n_3321),
.Y(n_4060)
);

INVx2_ASAP7_75t_SL g4061 ( 
.A(n_3321),
.Y(n_4061)
);

BUFx3_ASAP7_75t_L g4062 ( 
.A(n_3704),
.Y(n_4062)
);

NOR2xp33_ASAP7_75t_L g4063 ( 
.A(n_3604),
.B(n_371),
.Y(n_4063)
);

INVx3_ASAP7_75t_L g4064 ( 
.A(n_3342),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3317),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3337),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3732),
.B(n_3344),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3641),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3490),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3366),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3780),
.B(n_372),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3648),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3649),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3679),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3786),
.B(n_3806),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3810),
.B(n_372),
.Y(n_4076)
);

BUFx6f_ASAP7_75t_L g4077 ( 
.A(n_3366),
.Y(n_4077)
);

AOI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_3564),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_4078)
);

INVx3_ASAP7_75t_L g4079 ( 
.A(n_3342),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3345),
.Y(n_4080)
);

OR2x4_ASAP7_75t_L g4081 ( 
.A(n_3382),
.B(n_374),
.Y(n_4081)
);

AND2x6_ASAP7_75t_SL g4082 ( 
.A(n_3714),
.B(n_958),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3686),
.Y(n_4083)
);

BUFx6f_ASAP7_75t_L g4084 ( 
.A(n_3366),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3721),
.B(n_376),
.Y(n_4085)
);

CKINVDCx5p33_ASAP7_75t_R g4086 ( 
.A(n_3472),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3737),
.B(n_377),
.Y(n_4087)
);

A2O1A1Ixp33_ASAP7_75t_L g4088 ( 
.A1(n_3768),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3684),
.B(n_379),
.Y(n_4089)
);

NAND2x1p5_ASAP7_75t_L g4090 ( 
.A(n_3517),
.B(n_380),
.Y(n_4090)
);

INVx3_ASAP7_75t_L g4091 ( 
.A(n_3343),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3265),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3270),
.B(n_381),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3280),
.B(n_381),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3355),
.Y(n_4095)
);

BUFx3_ASAP7_75t_L g4096 ( 
.A(n_3595),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3281),
.B(n_382),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3772),
.B(n_3747),
.Y(n_4098)
);

OR2x6_ASAP7_75t_L g4099 ( 
.A(n_3714),
.B(n_382),
.Y(n_4099)
);

AOI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_3417),
.A2(n_386),
.B1(n_383),
.B2(n_385),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3725),
.B(n_383),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3729),
.B(n_387),
.Y(n_4102)
);

BUFx2_ASAP7_75t_L g4103 ( 
.A(n_3424),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3359),
.Y(n_4104)
);

AND2x4_ASAP7_75t_L g4105 ( 
.A(n_3550),
.B(n_387),
.Y(n_4105)
);

NAND3xp33_ASAP7_75t_SL g4106 ( 
.A(n_3645),
.B(n_388),
.C(n_389),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3397),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3401),
.Y(n_4108)
);

NOR2xp33_ASAP7_75t_L g4109 ( 
.A(n_3766),
.B(n_388),
.Y(n_4109)
);

O2A1O1Ixp33_ASAP7_75t_L g4110 ( 
.A1(n_3529),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_4110)
);

INVx2_ASAP7_75t_SL g4111 ( 
.A(n_3343),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3739),
.B(n_390),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_3655),
.B(n_393),
.Y(n_4113)
);

AO22x1_ASAP7_75t_L g4114 ( 
.A1(n_3550),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_4114)
);

AND2x4_ASAP7_75t_L g4115 ( 
.A(n_3630),
.B(n_395),
.Y(n_4115)
);

OR2x6_ASAP7_75t_L g4116 ( 
.A(n_3454),
.B(n_3809),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3313),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_3298),
.B(n_397),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_3743),
.B(n_397),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3418),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3523),
.A2(n_3295),
.B1(n_3690),
.B2(n_3396),
.Y(n_4121)
);

INVx2_ASAP7_75t_SL g4122 ( 
.A(n_3374),
.Y(n_4122)
);

AND2x6_ASAP7_75t_SL g4123 ( 
.A(n_3681),
.B(n_966),
.Y(n_4123)
);

OAI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3329),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4124)
);

AO22x1_ASAP7_75t_L g4125 ( 
.A1(n_3681),
.A2(n_402),
.B1(n_398),
.B2(n_401),
.Y(n_4125)
);

NOR2x1p5_ASAP7_75t_SL g4126 ( 
.A(n_3783),
.B(n_401),
.Y(n_4126)
);

AOI22xp5_ASAP7_75t_SL g4127 ( 
.A1(n_3274),
.A2(n_3351),
.B1(n_3752),
.B2(n_3486),
.Y(n_4127)
);

AND2x4_ASAP7_75t_L g4128 ( 
.A(n_3712),
.B(n_402),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3318),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3289),
.A2(n_3671),
.B(n_3598),
.Y(n_4130)
);

INVxp67_ASAP7_75t_L g4131 ( 
.A(n_3327),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3322),
.Y(n_4132)
);

OR2x6_ASAP7_75t_L g4133 ( 
.A(n_3809),
.B(n_403),
.Y(n_4133)
);

OR2x2_ASAP7_75t_L g4134 ( 
.A(n_3338),
.B(n_403),
.Y(n_4134)
);

INVx3_ASAP7_75t_L g4135 ( 
.A(n_3374),
.Y(n_4135)
);

INVx3_ASAP7_75t_L g4136 ( 
.A(n_3705),
.Y(n_4136)
);

AOI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_3543),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3425),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3742),
.B(n_404),
.Y(n_4139)
);

INVx5_ASAP7_75t_L g4140 ( 
.A(n_3405),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_3545),
.B(n_3674),
.Y(n_4141)
);

OAI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_3346),
.A2(n_406),
.B(n_407),
.Y(n_4142)
);

INVx3_ASAP7_75t_L g4143 ( 
.A(n_3579),
.Y(n_4143)
);

INVx1_ASAP7_75t_SL g4144 ( 
.A(n_3473),
.Y(n_4144)
);

BUFx6f_ASAP7_75t_L g4145 ( 
.A(n_3517),
.Y(n_4145)
);

AND2x4_ASAP7_75t_L g4146 ( 
.A(n_3736),
.B(n_407),
.Y(n_4146)
);

INVx1_ASAP7_75t_SL g4147 ( 
.A(n_3627),
.Y(n_4147)
);

INVx1_ASAP7_75t_SL g4148 ( 
.A(n_3502),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_3432),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3460),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3464),
.Y(n_4151)
);

AND2x6_ASAP7_75t_L g4152 ( 
.A(n_3727),
.B(n_408),
.Y(n_4152)
);

INVx2_ASAP7_75t_SL g4153 ( 
.A(n_3579),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_3748),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_4154)
);

AND2x4_ASAP7_75t_L g4155 ( 
.A(n_3711),
.B(n_409),
.Y(n_4155)
);

OR2x2_ASAP7_75t_SL g4156 ( 
.A(n_3667),
.B(n_3817),
.Y(n_4156)
);

OAI21x1_ASAP7_75t_L g4157 ( 
.A1(n_3796),
.A2(n_3778),
.B(n_3781),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3326),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3466),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_3568),
.Y(n_4160)
);

INVxp67_ASAP7_75t_L g4161 ( 
.A(n_3339),
.Y(n_4161)
);

INVx4_ASAP7_75t_L g4162 ( 
.A(n_3517),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3717),
.B(n_3722),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3795),
.B(n_410),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3330),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3782),
.B(n_411),
.Y(n_4166)
);

INVx1_ASAP7_75t_SL g4167 ( 
.A(n_3410),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3332),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3335),
.Y(n_4169)
);

AND2x4_ASAP7_75t_L g4170 ( 
.A(n_3711),
.B(n_414),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3774),
.B(n_414),
.Y(n_4171)
);

HB1xp67_ASAP7_75t_L g4172 ( 
.A(n_3708),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3349),
.Y(n_4173)
);

INVx4_ASAP7_75t_L g4174 ( 
.A(n_3548),
.Y(n_4174)
);

HB1xp67_ASAP7_75t_L g4175 ( 
.A(n_3754),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3353),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3477),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_3804),
.B(n_415),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3558),
.B(n_3390),
.Y(n_4179)
);

BUFx3_ASAP7_75t_L g4180 ( 
.A(n_3665),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3495),
.Y(n_4181)
);

BUFx2_ASAP7_75t_L g4182 ( 
.A(n_3548),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3554),
.B(n_416),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3559),
.B(n_417),
.Y(n_4184)
);

INVx4_ASAP7_75t_L g4185 ( 
.A(n_3548),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_L g4186 ( 
.A(n_3822),
.B(n_417),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_3497),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_L g4188 ( 
.A(n_3536),
.B(n_418),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3503),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3514),
.Y(n_4190)
);

AND2x4_ASAP7_75t_L g4191 ( 
.A(n_3804),
.B(n_419),
.Y(n_4191)
);

AND3x1_ASAP7_75t_SL g4192 ( 
.A(n_3770),
.B(n_420),
.C(n_421),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_3790),
.B(n_420),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3527),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3530),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3531),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3534),
.Y(n_4197)
);

INVx3_ASAP7_75t_L g4198 ( 
.A(n_3581),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_3707),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_4199)
);

INVx2_ASAP7_75t_SL g4200 ( 
.A(n_3581),
.Y(n_4200)
);

BUFx2_ASAP7_75t_L g4201 ( 
.A(n_3569),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_3629),
.B(n_423),
.Y(n_4202)
);

BUFx12f_ASAP7_75t_L g4203 ( 
.A(n_3701),
.Y(n_4203)
);

OAI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_3448),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_4204)
);

AND2x4_ASAP7_75t_L g4205 ( 
.A(n_3816),
.B(n_426),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_3540),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3566),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_3699),
.B(n_428),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3610),
.Y(n_4209)
);

HB1xp67_ASAP7_75t_L g4210 ( 
.A(n_3757),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_3808),
.B(n_428),
.Y(n_4211)
);

BUFx6f_ASAP7_75t_L g4212 ( 
.A(n_3569),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3607),
.B(n_429),
.Y(n_4213)
);

OR2x4_ASAP7_75t_L g4214 ( 
.A(n_3314),
.B(n_429),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3612),
.Y(n_4215)
);

INVx4_ASAP7_75t_L g4216 ( 
.A(n_3569),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3476),
.B(n_430),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3618),
.Y(n_4218)
);

BUFx12f_ASAP7_75t_L g4219 ( 
.A(n_3680),
.Y(n_4219)
);

INVx2_ASAP7_75t_SL g4220 ( 
.A(n_3642),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3651),
.Y(n_4221)
);

HB1xp67_ASAP7_75t_L g4222 ( 
.A(n_3677),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_3678),
.Y(n_4223)
);

AO221x1_ASAP7_75t_L g4224 ( 
.A1(n_3449),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.C(n_434),
.Y(n_4224)
);

AO32x2_ASAP7_75t_L g4225 ( 
.A1(n_3981),
.A2(n_3555),
.A3(n_3561),
.B1(n_3776),
.B2(n_3478),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4141),
.B(n_3556),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_L g4227 ( 
.A1(n_4157),
.A2(n_3813),
.B(n_3574),
.Y(n_4227)
);

AOI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_3947),
.A2(n_3799),
.B1(n_3348),
.B2(n_3367),
.Y(n_4228)
);

OAI21x1_ASAP7_75t_L g4229 ( 
.A1(n_3887),
.A2(n_3798),
.B(n_3793),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_3979),
.B(n_3556),
.Y(n_4230)
);

BUFx12f_ASAP7_75t_L g4231 ( 
.A(n_3840),
.Y(n_4231)
);

NOR2x1_ASAP7_75t_SL g4232 ( 
.A(n_4116),
.B(n_3510),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3829),
.Y(n_4233)
);

AO21x1_ASAP7_75t_L g4234 ( 
.A1(n_3878),
.A2(n_3775),
.B(n_3727),
.Y(n_4234)
);

AO21x2_ASAP7_75t_L g4235 ( 
.A1(n_4057),
.A2(n_3635),
.B(n_3393),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3862),
.B(n_3802),
.Y(n_4236)
);

HB1xp67_ASAP7_75t_L g4237 ( 
.A(n_4001),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_3993),
.A2(n_3650),
.B(n_3614),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3827),
.Y(n_4239)
);

AO31x2_ASAP7_75t_L g4240 ( 
.A1(n_4028),
.A2(n_3429),
.A3(n_3715),
.B(n_3741),
.Y(n_4240)
);

INVx4_ASAP7_75t_L g4241 ( 
.A(n_3824),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4075),
.B(n_3792),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4054),
.B(n_3811),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_3876),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3832),
.B(n_3818),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_3925),
.A2(n_3937),
.B(n_3963),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_SL g4247 ( 
.A1(n_4099),
.A2(n_3458),
.B(n_3427),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_4029),
.A2(n_3602),
.B(n_3597),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_3826),
.B(n_3680),
.Y(n_4249)
);

BUFx12f_ASAP7_75t_L g4250 ( 
.A(n_3865),
.Y(n_4250)
);

INVx3_ASAP7_75t_L g4251 ( 
.A(n_3834),
.Y(n_4251)
);

NAND2x1_ASAP7_75t_L g4252 ( 
.A(n_4152),
.B(n_3775),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_3833),
.B(n_3560),
.Y(n_4253)
);

CKINVDCx8_ASAP7_75t_R g4254 ( 
.A(n_4082),
.Y(n_4254)
);

AOI211x1_ASAP7_75t_L g4255 ( 
.A1(n_4125),
.A2(n_3512),
.B(n_3544),
.C(n_3488),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3852),
.B(n_3573),
.Y(n_4256)
);

AO21x2_ASAP7_75t_L g4257 ( 
.A1(n_3847),
.A2(n_3626),
.B(n_3621),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_4015),
.Y(n_4258)
);

OAI21x1_ASAP7_75t_L g4259 ( 
.A1(n_3889),
.A2(n_3896),
.B(n_3884),
.Y(n_4259)
);

OAI22x1_ASAP7_75t_L g4260 ( 
.A1(n_3951),
.A2(n_3663),
.B1(n_3286),
.B2(n_3669),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_SL g4261 ( 
.A(n_4127),
.B(n_3567),
.Y(n_4261)
);

OAI21x1_ASAP7_75t_L g4262 ( 
.A1(n_4130),
.A2(n_3791),
.B(n_3773),
.Y(n_4262)
);

NAND2x1p5_ASAP7_75t_L g4263 ( 
.A(n_3848),
.B(n_3642),
.Y(n_4263)
);

OAI21x1_ASAP7_75t_L g4264 ( 
.A1(n_4037),
.A2(n_3762),
.B(n_3698),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_3939),
.A2(n_3654),
.B(n_3638),
.Y(n_4265)
);

AOI21xp33_ASAP7_75t_L g4266 ( 
.A1(n_3854),
.A2(n_3470),
.B(n_3468),
.Y(n_4266)
);

AOI21xp33_ASAP7_75t_L g4267 ( 
.A1(n_3943),
.A2(n_3481),
.B(n_3480),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_3950),
.A2(n_3685),
.B(n_3662),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3855),
.B(n_3575),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3866),
.B(n_3587),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4038),
.A2(n_3697),
.B(n_3413),
.Y(n_4271)
);

OAI21x1_ASAP7_75t_L g4272 ( 
.A1(n_4031),
.A2(n_3520),
.B(n_3394),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3868),
.Y(n_4273)
);

OAI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_4088),
.A2(n_3407),
.B(n_3582),
.Y(n_4274)
);

INVx2_ASAP7_75t_SL g4275 ( 
.A(n_3841),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4048),
.B(n_3518),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4113),
.B(n_3692),
.Y(n_4277)
);

NAND3xp33_ASAP7_75t_SL g4278 ( 
.A(n_3997),
.B(n_3340),
.C(n_3613),
.Y(n_4278)
);

BUFx2_ASAP7_75t_L g4279 ( 
.A(n_3838),
.Y(n_4279)
);

INVx3_ASAP7_75t_L g4280 ( 
.A(n_3883),
.Y(n_4280)
);

OAI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_3845),
.A2(n_3498),
.B(n_3676),
.Y(n_4281)
);

OAI21x1_ASAP7_75t_L g4282 ( 
.A1(n_3906),
.A2(n_3652),
.B(n_3373),
.Y(n_4282)
);

OAI21x1_ASAP7_75t_L g4283 ( 
.A1(n_3918),
.A2(n_3319),
.B(n_3586),
.Y(n_4283)
);

OAI22xp5_ASAP7_75t_L g4284 ( 
.A1(n_4133),
.A2(n_3784),
.B1(n_3590),
.B2(n_3606),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4020),
.Y(n_4285)
);

OAI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4142),
.A2(n_3821),
.B(n_3753),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3869),
.B(n_3603),
.Y(n_4287)
);

AND2x4_ASAP7_75t_L g4288 ( 
.A(n_4116),
.B(n_3594),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3873),
.B(n_3751),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_SL g4290 ( 
.A(n_4022),
.B(n_3644),
.Y(n_4290)
);

OAI21x1_ASAP7_75t_L g4291 ( 
.A1(n_3928),
.A2(n_3749),
.B(n_3700),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_3891),
.Y(n_4292)
);

INVx6_ASAP7_75t_L g4293 ( 
.A(n_3900),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_3894),
.B(n_3381),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3927),
.Y(n_4295)
);

OAI21x1_ASAP7_75t_L g4296 ( 
.A1(n_3938),
.A2(n_3750),
.B(n_3399),
.Y(n_4296)
);

NOR4xp25_ASAP7_75t_L g4297 ( 
.A(n_4109),
.B(n_3633),
.C(n_3706),
.D(n_3702),
.Y(n_4297)
);

OAI21x1_ASAP7_75t_L g4298 ( 
.A1(n_3959),
.A2(n_3461),
.B(n_3386),
.Y(n_4298)
);

OAI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_4199),
.A2(n_3591),
.B(n_3683),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4175),
.A2(n_3413),
.B(n_3405),
.Y(n_4300)
);

OAI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_3858),
.A2(n_3634),
.B(n_3624),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4210),
.A2(n_3413),
.B(n_3405),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3929),
.B(n_3463),
.Y(n_4303)
);

OAI22xp5_ASAP7_75t_L g4304 ( 
.A1(n_4133),
.A2(n_3542),
.B1(n_3422),
.B2(n_3580),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_4179),
.A2(n_3557),
.B(n_3474),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_SL g4306 ( 
.A(n_3935),
.B(n_3637),
.C(n_3371),
.Y(n_4306)
);

NAND2x1_ASAP7_75t_L g4307 ( 
.A(n_4152),
.B(n_3814),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_3931),
.B(n_3414),
.Y(n_4308)
);

OAI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4121),
.A2(n_3636),
.B(n_3735),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_3882),
.A2(n_3557),
.B(n_3474),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_SL g4311 ( 
.A(n_4019),
.B(n_3474),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_L g4312 ( 
.A1(n_4222),
.A2(n_3592),
.B(n_3557),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3933),
.Y(n_4313)
);

OAI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_3971),
.A2(n_3787),
.B(n_3785),
.Y(n_4314)
);

INVx2_ASAP7_75t_SL g4315 ( 
.A(n_3853),
.Y(n_4315)
);

AOI21x1_ASAP7_75t_L g4316 ( 
.A1(n_3842),
.A2(n_3484),
.B(n_3759),
.Y(n_4316)
);

AO31x2_ASAP7_75t_L g4317 ( 
.A1(n_3968),
.A2(n_3525),
.A3(n_3522),
.B(n_3426),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3944),
.B(n_3434),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_SL g4319 ( 
.A(n_3970),
.B(n_3592),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_3965),
.B(n_3442),
.Y(n_4320)
);

OAI21x1_ASAP7_75t_L g4321 ( 
.A1(n_3967),
.A2(n_4003),
.B(n_3973),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_3924),
.A2(n_3625),
.B(n_3592),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3972),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_3844),
.Y(n_4324)
);

INVx3_ASAP7_75t_SL g4325 ( 
.A(n_3872),
.Y(n_4325)
);

OAI21x1_ASAP7_75t_L g4326 ( 
.A1(n_4006),
.A2(n_3459),
.B(n_3447),
.Y(n_4326)
);

OAI21x1_ASAP7_75t_SL g4327 ( 
.A1(n_4033),
.A2(n_3620),
.B(n_3611),
.Y(n_4327)
);

INVx4_ASAP7_75t_L g4328 ( 
.A(n_3920),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_3932),
.A2(n_3625),
.B(n_3718),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4023),
.Y(n_4330)
);

BUFx2_ASAP7_75t_L g4331 ( 
.A(n_4069),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3987),
.B(n_3552),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_3899),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_3988),
.B(n_3682),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_3991),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4046),
.Y(n_4336)
);

BUFx2_ASAP7_75t_L g4337 ( 
.A(n_4042),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_3851),
.B(n_3815),
.Y(n_4338)
);

OAI21x1_ASAP7_75t_L g4339 ( 
.A1(n_3886),
.A2(n_3733),
.B(n_3710),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4010),
.B(n_4000),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4065),
.Y(n_4341)
);

INVx4_ASAP7_75t_L g4342 ( 
.A(n_3905),
.Y(n_4342)
);

OAI21x1_ASAP7_75t_L g4343 ( 
.A1(n_3898),
.A2(n_3734),
.B(n_3769),
.Y(n_4343)
);

OAI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4011),
.A2(n_3819),
.B(n_3789),
.Y(n_4344)
);

OAI21xp5_ASAP7_75t_L g4345 ( 
.A1(n_3976),
.A2(n_3709),
.B(n_3719),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4089),
.B(n_3682),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4002),
.B(n_3616),
.Y(n_4347)
);

OAI21x1_ASAP7_75t_L g4348 ( 
.A1(n_4009),
.A2(n_3647),
.B(n_3643),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4092),
.B(n_3437),
.Y(n_4349)
);

AND2x4_ASAP7_75t_L g4350 ( 
.A(n_4062),
.B(n_3642),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_3910),
.B(n_3740),
.Y(n_4351)
);

BUFx8_ASAP7_75t_SL g4352 ( 
.A(n_3879),
.Y(n_4352)
);

INVx3_ASAP7_75t_L g4353 ( 
.A(n_3961),
.Y(n_4353)
);

AOI211x1_ASAP7_75t_L g4354 ( 
.A1(n_4114),
.A2(n_4208),
.B(n_4106),
.C(n_4040),
.Y(n_4354)
);

OAI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4110),
.A2(n_3745),
.B(n_3728),
.Y(n_4355)
);

OAI21x1_ASAP7_75t_SL g4356 ( 
.A1(n_4061),
.A2(n_3584),
.B(n_3436),
.Y(n_4356)
);

OAI21x1_ASAP7_75t_L g4357 ( 
.A1(n_4016),
.A2(n_4039),
.B(n_4036),
.Y(n_4357)
);

AOI22xp5_ASAP7_75t_L g4358 ( 
.A1(n_3867),
.A2(n_3521),
.B1(n_3672),
.B2(n_3589),
.Y(n_4358)
);

OAI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4099),
.A2(n_3453),
.B1(n_3456),
.B2(n_3391),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3893),
.Y(n_4360)
);

INVx3_ASAP7_75t_L g4361 ( 
.A(n_4219),
.Y(n_4361)
);

AOI31xp67_ASAP7_75t_L g4362 ( 
.A1(n_4024),
.A2(n_3659),
.A3(n_3666),
.B(n_3661),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4117),
.B(n_3797),
.Y(n_4363)
);

OAI21x1_ASAP7_75t_L g4364 ( 
.A1(n_4043),
.A2(n_3670),
.B(n_3668),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4129),
.B(n_4132),
.Y(n_4365)
);

INVxp67_ASAP7_75t_L g4366 ( 
.A(n_3995),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4158),
.B(n_3492),
.Y(n_4367)
);

INVx1_ASAP7_75t_SL g4368 ( 
.A(n_3828),
.Y(n_4368)
);

INVx5_ASAP7_75t_L g4369 ( 
.A(n_4145),
.Y(n_4369)
);

INVxp67_ASAP7_75t_L g4370 ( 
.A(n_3903),
.Y(n_4370)
);

CKINVDCx20_ASAP7_75t_R g4371 ( 
.A(n_3892),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_3913),
.Y(n_4372)
);

OAI21x1_ASAP7_75t_L g4373 ( 
.A1(n_4052),
.A2(n_3765),
.B(n_3713),
.Y(n_4373)
);

INVx1_ASAP7_75t_SL g4374 ( 
.A(n_3911),
.Y(n_4374)
);

INVxp67_ASAP7_75t_SL g4375 ( 
.A(n_4056),
.Y(n_4375)
);

OAI21x1_ASAP7_75t_SL g4376 ( 
.A1(n_4111),
.A2(n_3628),
.B(n_3731),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4044),
.B(n_431),
.Y(n_4377)
);

OAI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_3860),
.A2(n_3755),
.B(n_3746),
.Y(n_4378)
);

OAI21x1_ASAP7_75t_L g4379 ( 
.A1(n_4068),
.A2(n_3794),
.B(n_3767),
.Y(n_4379)
);

OAI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_4018),
.A2(n_4124),
.B(n_4007),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4165),
.B(n_3640),
.Y(n_4381)
);

AOI21x1_ASAP7_75t_L g4382 ( 
.A1(n_4182),
.A2(n_3761),
.B(n_3756),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_4168),
.B(n_4169),
.Y(n_4383)
);

OAI21xp5_ASAP7_75t_L g4384 ( 
.A1(n_3907),
.A2(n_3764),
.B(n_3800),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4173),
.B(n_3673),
.Y(n_4385)
);

A2O1A1Ixp33_ASAP7_75t_L g4386 ( 
.A1(n_4030),
.A2(n_3807),
.B(n_3803),
.C(n_3805),
.Y(n_4386)
);

OAI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_4204),
.A2(n_3820),
.B(n_3693),
.Y(n_4387)
);

AO31x2_ASAP7_75t_L g4388 ( 
.A1(n_4098),
.A2(n_3625),
.A3(n_3696),
.B(n_3646),
.Y(n_4388)
);

OAI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_3839),
.A2(n_3687),
.B(n_3696),
.Y(n_4389)
);

O2A1O1Ixp5_ASAP7_75t_SL g4390 ( 
.A1(n_3908),
.A2(n_3696),
.B(n_435),
.C(n_432),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4176),
.B(n_3646),
.Y(n_4391)
);

OAI21x1_ASAP7_75t_L g4392 ( 
.A1(n_4072),
.A2(n_444),
.B(n_433),
.Y(n_4392)
);

NOR4xp25_ASAP7_75t_L g4393 ( 
.A(n_3930),
.B(n_438),
.C(n_436),
.D(n_437),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4073),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_4074),
.B(n_436),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4083),
.B(n_437),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4066),
.Y(n_4397)
);

AOI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_4153),
.A2(n_4200),
.B(n_4198),
.Y(n_4398)
);

AO31x2_ASAP7_75t_L g4399 ( 
.A1(n_4080),
.A2(n_440),
.A3(n_438),
.B(n_439),
.Y(n_4399)
);

AND2x4_ASAP7_75t_L g4400 ( 
.A(n_4136),
.B(n_4041),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_4143),
.A2(n_4104),
.B(n_4095),
.Y(n_4401)
);

O2A1O1Ixp5_ASAP7_75t_L g4402 ( 
.A1(n_4162),
.A2(n_4185),
.B(n_4216),
.C(n_4174),
.Y(n_4402)
);

BUFx2_ASAP7_75t_L g4403 ( 
.A(n_4201),
.Y(n_4403)
);

OAI21x1_ASAP7_75t_L g4404 ( 
.A1(n_4107),
.A2(n_450),
.B(n_440),
.Y(n_4404)
);

OAI21x1_ASAP7_75t_L g4405 ( 
.A1(n_4108),
.A2(n_452),
.B(n_442),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4131),
.B(n_443),
.Y(n_4406)
);

OAI21x1_ASAP7_75t_L g4407 ( 
.A1(n_4120),
.A2(n_453),
.B(n_443),
.Y(n_4407)
);

BUFx12f_ASAP7_75t_L g4408 ( 
.A(n_3880),
.Y(n_4408)
);

NAND2xp33_ASAP7_75t_SL g4409 ( 
.A(n_3984),
.B(n_444),
.Y(n_4409)
);

O2A1O1Ixp5_ASAP7_75t_SL g4410 ( 
.A1(n_3926),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_4410)
);

AND2x2_ASAP7_75t_SL g4411 ( 
.A(n_4178),
.B(n_962),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_3874),
.B(n_4177),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4181),
.B(n_445),
.Y(n_4413)
);

INVxp67_ASAP7_75t_L g4414 ( 
.A(n_3957),
.Y(n_4414)
);

HB1xp67_ASAP7_75t_L g4415 ( 
.A(n_3831),
.Y(n_4415)
);

AND2x4_ASAP7_75t_L g4416 ( 
.A(n_4096),
.B(n_446),
.Y(n_4416)
);

BUFx2_ASAP7_75t_L g4417 ( 
.A(n_4145),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4189),
.Y(n_4418)
);

AOI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_4138),
.A2(n_449),
.B(n_451),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4190),
.Y(n_4420)
);

OAI21xp5_ASAP7_75t_L g4421 ( 
.A1(n_3990),
.A2(n_451),
.B(n_452),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4197),
.B(n_4207),
.Y(n_4422)
);

NOR2xp33_ASAP7_75t_L g4423 ( 
.A(n_4081),
.B(n_945),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_L g4424 ( 
.A1(n_4149),
.A2(n_462),
.B(n_454),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4105),
.B(n_454),
.Y(n_4425)
);

OAI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4034),
.A2(n_455),
.B(n_456),
.Y(n_4426)
);

BUFx2_ASAP7_75t_L g4427 ( 
.A(n_4212),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4150),
.A2(n_456),
.B(n_457),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4209),
.B(n_457),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4151),
.A2(n_4187),
.B(n_4159),
.Y(n_4430)
);

INVx8_ASAP7_75t_L g4431 ( 
.A(n_4123),
.Y(n_4431)
);

AOI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_4194),
.A2(n_4196),
.B(n_4195),
.Y(n_4432)
);

OA21x2_ASAP7_75t_L g4433 ( 
.A1(n_3948),
.A2(n_458),
.B(n_459),
.Y(n_4433)
);

INVx3_ASAP7_75t_L g4434 ( 
.A(n_4212),
.Y(n_4434)
);

OAI21x1_ASAP7_75t_L g4435 ( 
.A1(n_4206),
.A2(n_468),
.B(n_459),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4215),
.B(n_460),
.Y(n_4436)
);

AOI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_4221),
.A2(n_460),
.B(n_461),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4218),
.B(n_463),
.Y(n_4438)
);

CKINVDCx5p33_ASAP7_75t_R g4439 ( 
.A(n_3881),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4223),
.Y(n_4440)
);

OAI21x1_ASAP7_75t_SL g4441 ( 
.A1(n_4122),
.A2(n_463),
.B(n_464),
.Y(n_4441)
);

OAI21x1_ASAP7_75t_L g4442 ( 
.A1(n_4060),
.A2(n_473),
.B(n_465),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3912),
.B(n_466),
.Y(n_4443)
);

OAI21x1_ASAP7_75t_L g4444 ( 
.A1(n_4064),
.A2(n_476),
.B(n_467),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_SL g4445 ( 
.A(n_4140),
.B(n_468),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4163),
.B(n_469),
.Y(n_4446)
);

AO32x2_ASAP7_75t_L g4447 ( 
.A1(n_3915),
.A2(n_471),
.A3(n_469),
.B1(n_470),
.B2(n_472),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4079),
.A2(n_484),
.B(n_470),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_3856),
.B(n_474),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_3849),
.Y(n_4450)
);

HB1xp67_ASAP7_75t_L g4451 ( 
.A(n_4172),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_3922),
.B(n_474),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_3941),
.Y(n_4453)
);

OAI21x1_ASAP7_75t_L g4454 ( 
.A1(n_4091),
.A2(n_486),
.B(n_475),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4144),
.B(n_475),
.Y(n_4455)
);

OA22x2_ASAP7_75t_L g4456 ( 
.A1(n_3888),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_4456)
);

OAI21x1_ASAP7_75t_L g4457 ( 
.A1(n_4135),
.A2(n_487),
.B(n_478),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3895),
.B(n_479),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4148),
.B(n_480),
.Y(n_4459)
);

OAI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_4154),
.A2(n_481),
.B(n_483),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_3953),
.B(n_3949),
.Y(n_4461)
);

A2O1A1Ixp33_ASAP7_75t_L g4462 ( 
.A1(n_4191),
.A2(n_484),
.B(n_481),
.C(n_483),
.Y(n_4462)
);

AND2x2_ASAP7_75t_SL g4463 ( 
.A(n_4155),
.B(n_967),
.Y(n_4463)
);

BUFx3_ASAP7_75t_L g4464 ( 
.A(n_3830),
.Y(n_4464)
);

NOR2xp67_ASAP7_75t_L g4465 ( 
.A(n_4005),
.B(n_485),
.Y(n_4465)
);

OR2x6_ASAP7_75t_L g4466 ( 
.A(n_4021),
.B(n_485),
.Y(n_4466)
);

OA22x2_ASAP7_75t_L g4467 ( 
.A1(n_3888),
.A2(n_488),
.B1(n_486),
.B2(n_487),
.Y(n_4467)
);

OAI21x1_ASAP7_75t_SL g4468 ( 
.A1(n_4100),
.A2(n_489),
.B(n_490),
.Y(n_4468)
);

OAI21x1_ASAP7_75t_L g4469 ( 
.A1(n_4090),
.A2(n_501),
.B(n_489),
.Y(n_4469)
);

INVxp67_ASAP7_75t_SL g4470 ( 
.A(n_3875),
.Y(n_4470)
);

NAND2x1p5_ASAP7_75t_L g4471 ( 
.A(n_3934),
.B(n_491),
.Y(n_4471)
);

OAI21x1_ASAP7_75t_L g4472 ( 
.A1(n_3999),
.A2(n_502),
.B(n_491),
.Y(n_4472)
);

OAI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_4202),
.A2(n_495),
.B(n_496),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_3923),
.B(n_497),
.Y(n_4474)
);

AOI21xp5_ASAP7_75t_L g4475 ( 
.A1(n_3909),
.A2(n_497),
.B(n_498),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4103),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_3946),
.B(n_3958),
.Y(n_4477)
);

OAI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_4161),
.A2(n_4119),
.B(n_4012),
.Y(n_4478)
);

BUFx2_ASAP7_75t_SL g4479 ( 
.A(n_3837),
.Y(n_4479)
);

OAI21x1_ASAP7_75t_L g4480 ( 
.A1(n_4053),
.A2(n_506),
.B(n_498),
.Y(n_4480)
);

OAI21x1_ASAP7_75t_L g4481 ( 
.A1(n_3877),
.A2(n_507),
.B(n_499),
.Y(n_4481)
);

AO31x2_ASAP7_75t_L g4482 ( 
.A1(n_4094),
.A2(n_501),
.A3(n_499),
.B(n_500),
.Y(n_4482)
);

NAND2x1p5_ASAP7_75t_L g4483 ( 
.A(n_3978),
.B(n_500),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_SL g4484 ( 
.A(n_4140),
.B(n_502),
.Y(n_4484)
);

AO31x2_ASAP7_75t_L g4485 ( 
.A1(n_4097),
.A2(n_4184),
.A3(n_4213),
.B(n_4183),
.Y(n_4485)
);

NOR2x1_ASAP7_75t_SL g4486 ( 
.A(n_4021),
.B(n_3956),
.Y(n_4486)
);

OAI21x1_ASAP7_75t_L g4487 ( 
.A1(n_3885),
.A2(n_511),
.B(n_503),
.Y(n_4487)
);

OAI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_4137),
.A2(n_503),
.B(n_504),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_SL g4489 ( 
.A(n_3902),
.B(n_504),
.Y(n_4489)
);

AND2x4_ASAP7_75t_L g4490 ( 
.A(n_3936),
.B(n_505),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_3835),
.B(n_4214),
.Y(n_4491)
);

AOI221xp5_ASAP7_75t_SL g4492 ( 
.A1(n_4186),
.A2(n_953),
.B1(n_944),
.B2(n_508),
.C(n_506),
.Y(n_4492)
);

O2A1O1Ixp5_ASAP7_75t_L g4493 ( 
.A1(n_4026),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_4493)
);

OAI21x1_ASAP7_75t_L g4494 ( 
.A1(n_3904),
.A2(n_4085),
.B(n_4101),
.Y(n_4494)
);

BUFx6f_ASAP7_75t_L g4495 ( 
.A(n_4180),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_3864),
.Y(n_4496)
);

AOI21xp33_ASAP7_75t_L g4497 ( 
.A1(n_3909),
.A2(n_509),
.B(n_510),
.Y(n_4497)
);

NOR2x1_ASAP7_75t_SL g4498 ( 
.A(n_3956),
.B(n_3914),
.Y(n_4498)
);

OAI21xp33_ASAP7_75t_L g4499 ( 
.A1(n_4126),
.A2(n_510),
.B(n_511),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_3960),
.B(n_512),
.Y(n_4500)
);

AO31x2_ASAP7_75t_L g4501 ( 
.A1(n_4013),
.A2(n_516),
.A3(n_513),
.B(n_514),
.Y(n_4501)
);

AO21x1_ASAP7_75t_L g4502 ( 
.A1(n_4146),
.A2(n_4170),
.B(n_4193),
.Y(n_4502)
);

NOR2xp33_ASAP7_75t_L g4503 ( 
.A(n_4032),
.B(n_959),
.Y(n_4503)
);

INVxp67_ASAP7_75t_L g4504 ( 
.A(n_3955),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_4160),
.B(n_4147),
.Y(n_4505)
);

OAI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_3836),
.A2(n_517),
.B(n_518),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_3964),
.B(n_518),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4164),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4067),
.B(n_519),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_3849),
.Y(n_4510)
);

OAI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_4078),
.A2(n_520),
.B(n_521),
.Y(n_4511)
);

AOI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_3914),
.A2(n_522),
.B(n_523),
.Y(n_4512)
);

OA21x2_ASAP7_75t_L g4513 ( 
.A1(n_4224),
.A2(n_523),
.B(n_524),
.Y(n_4513)
);

INVx4_ASAP7_75t_L g4514 ( 
.A(n_4027),
.Y(n_4514)
);

INVx1_ASAP7_75t_SL g4515 ( 
.A(n_3917),
.Y(n_4515)
);

AOI221xp5_ASAP7_75t_L g4516 ( 
.A1(n_4297),
.A2(n_4087),
.B1(n_4055),
.B2(n_4211),
.C(n_4217),
.Y(n_4516)
);

INVx1_ASAP7_75t_SL g4517 ( 
.A(n_4293),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_4360),
.B(n_4372),
.Y(n_4518)
);

BUFx3_ASAP7_75t_L g4519 ( 
.A(n_4293),
.Y(n_4519)
);

BUFx12f_ASAP7_75t_L g4520 ( 
.A(n_4231),
.Y(n_4520)
);

OAI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4463),
.A2(n_4156),
.B1(n_4167),
.B2(n_4205),
.Y(n_4521)
);

NAND3xp33_ASAP7_75t_L g4522 ( 
.A(n_4261),
.B(n_4188),
.C(n_4004),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4239),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4237),
.B(n_3901),
.Y(n_4524)
);

BUFx2_ASAP7_75t_L g4525 ( 
.A(n_4279),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4249),
.B(n_3945),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4233),
.Y(n_4527)
);

INVx5_ASAP7_75t_L g4528 ( 
.A(n_4241),
.Y(n_4528)
);

INVx3_ASAP7_75t_L g4529 ( 
.A(n_4328),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4412),
.B(n_3954),
.Y(n_4530)
);

AND2x4_ASAP7_75t_L g4531 ( 
.A(n_4486),
.B(n_3977),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_4244),
.Y(n_4532)
);

AOI22xp33_ASAP7_75t_L g4533 ( 
.A1(n_4306),
.A2(n_4152),
.B1(n_4128),
.B2(n_3975),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_4352),
.Y(n_4534)
);

BUFx2_ASAP7_75t_L g4535 ( 
.A(n_4403),
.Y(n_4535)
);

BUFx3_ASAP7_75t_L g4536 ( 
.A(n_4280),
.Y(n_4536)
);

AOI21x1_ASAP7_75t_L g4537 ( 
.A1(n_4382),
.A2(n_3940),
.B(n_4115),
.Y(n_4537)
);

HB1xp67_ASAP7_75t_L g4538 ( 
.A(n_4451),
.Y(n_4538)
);

CKINVDCx20_ASAP7_75t_R g4539 ( 
.A(n_4371),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_4252),
.A2(n_4220),
.B(n_3983),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4461),
.B(n_4058),
.Y(n_4541)
);

BUFx2_ASAP7_75t_L g4542 ( 
.A(n_4331),
.Y(n_4542)
);

NOR2xp67_ASAP7_75t_L g4543 ( 
.A(n_4342),
.B(n_4086),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4418),
.B(n_4118),
.Y(n_4544)
);

INVxp67_ASAP7_75t_SL g4545 ( 
.A(n_4415),
.Y(n_4545)
);

INVx4_ASAP7_75t_SL g4546 ( 
.A(n_4325),
.Y(n_4546)
);

OAI22xp5_ASAP7_75t_L g4547 ( 
.A1(n_4228),
.A2(n_4059),
.B1(n_3940),
.B2(n_4166),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4351),
.B(n_3980),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4420),
.B(n_4394),
.Y(n_4549)
);

AOI21xp5_ASAP7_75t_L g4550 ( 
.A1(n_4307),
.A2(n_3861),
.B(n_3850),
.Y(n_4550)
);

OAI22xp5_ASAP7_75t_SL g4551 ( 
.A1(n_4254),
.A2(n_3825),
.B1(n_4063),
.B2(n_4203),
.Y(n_4551)
);

AOI22xp33_ASAP7_75t_L g4552 ( 
.A1(n_4234),
.A2(n_3969),
.B1(n_3982),
.B2(n_3823),
.Y(n_4552)
);

AND2x4_ASAP7_75t_L g4553 ( 
.A(n_4498),
.B(n_3846),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4226),
.B(n_4035),
.Y(n_4554)
);

BUFx6f_ASAP7_75t_L g4555 ( 
.A(n_4495),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4258),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_L g4557 ( 
.A(n_4374),
.B(n_3863),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4285),
.Y(n_4558)
);

AOI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_4278),
.A2(n_4192),
.B1(n_3890),
.B2(n_3974),
.Y(n_4559)
);

INVx2_ASAP7_75t_SL g4560 ( 
.A(n_4495),
.Y(n_4560)
);

BUFx3_ASAP7_75t_L g4561 ( 
.A(n_4464),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_4333),
.Y(n_4562)
);

BUFx2_ASAP7_75t_L g4563 ( 
.A(n_4337),
.Y(n_4563)
);

AND2x4_ASAP7_75t_L g4564 ( 
.A(n_4400),
.B(n_4049),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4273),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4330),
.Y(n_4566)
);

INVx5_ASAP7_75t_L g4567 ( 
.A(n_4466),
.Y(n_4567)
);

HB1xp67_ASAP7_75t_L g4568 ( 
.A(n_4370),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4292),
.B(n_4134),
.Y(n_4569)
);

AND2x4_ASAP7_75t_L g4570 ( 
.A(n_4417),
.B(n_3850),
.Y(n_4570)
);

BUFx3_ASAP7_75t_L g4571 ( 
.A(n_4514),
.Y(n_4571)
);

OR2x2_ASAP7_75t_L g4572 ( 
.A(n_4470),
.B(n_4050),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4295),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4336),
.Y(n_4574)
);

INVx3_ASAP7_75t_L g4575 ( 
.A(n_4251),
.Y(n_4575)
);

BUFx6f_ASAP7_75t_L g4576 ( 
.A(n_4369),
.Y(n_4576)
);

AND2x4_ASAP7_75t_L g4577 ( 
.A(n_4427),
.B(n_3861),
.Y(n_4577)
);

BUFx3_ASAP7_75t_L g4578 ( 
.A(n_4275),
.Y(n_4578)
);

OR2x6_ASAP7_75t_L g4579 ( 
.A(n_4466),
.B(n_3989),
.Y(n_4579)
);

AOI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4246),
.A2(n_3897),
.B(n_3871),
.Y(n_4580)
);

BUFx6f_ASAP7_75t_L g4581 ( 
.A(n_4369),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4313),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4323),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4335),
.Y(n_4584)
);

NOR2xp33_ASAP7_75t_L g4585 ( 
.A(n_4431),
.B(n_3859),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_SL g4586 ( 
.A(n_4502),
.B(n_3857),
.Y(n_4586)
);

AOI21x1_ASAP7_75t_L g4587 ( 
.A1(n_4316),
.A2(n_3870),
.B(n_4171),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4319),
.A2(n_3897),
.B(n_3871),
.Y(n_4588)
);

BUFx2_ASAP7_75t_L g4589 ( 
.A(n_4369),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4496),
.B(n_4071),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4477),
.B(n_3994),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4366),
.B(n_4076),
.Y(n_4592)
);

A2O1A1Ixp33_ASAP7_75t_L g4593 ( 
.A1(n_4409),
.A2(n_3996),
.B(n_4008),
.C(n_4017),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4341),
.Y(n_4594)
);

BUFx3_ASAP7_75t_L g4595 ( 
.A(n_4353),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4340),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4515),
.B(n_3916),
.Y(n_4597)
);

AOI21xp5_ASAP7_75t_SL g4598 ( 
.A1(n_4232),
.A2(n_3919),
.B(n_3916),
.Y(n_4598)
);

NAND3xp33_ASAP7_75t_L g4599 ( 
.A(n_4354),
.B(n_4093),
.C(n_4102),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4357),
.Y(n_4600)
);

NOR2xp33_ASAP7_75t_L g4601 ( 
.A(n_4431),
.B(n_3843),
.Y(n_4601)
);

INVx1_ASAP7_75t_SL g4602 ( 
.A(n_4479),
.Y(n_4602)
);

OAI21x1_ASAP7_75t_L g4603 ( 
.A1(n_4227),
.A2(n_4259),
.B(n_4262),
.Y(n_4603)
);

BUFx12f_ASAP7_75t_L g4604 ( 
.A(n_4324),
.Y(n_4604)
);

BUFx3_ASAP7_75t_L g4605 ( 
.A(n_4315),
.Y(n_4605)
);

BUFx4_ASAP7_75t_SL g4606 ( 
.A(n_4439),
.Y(n_4606)
);

OAI31xp33_ASAP7_75t_L g4607 ( 
.A1(n_4284),
.A2(n_3998),
.A3(n_3992),
.B(n_3985),
.Y(n_4607)
);

BUFx3_ASAP7_75t_L g4608 ( 
.A(n_4361),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4365),
.B(n_4112),
.Y(n_4609)
);

A2O1A1Ixp33_ASAP7_75t_L g4610 ( 
.A1(n_4411),
.A2(n_4139),
.B(n_3921),
.C(n_3942),
.Y(n_4610)
);

AOI21xp5_ASAP7_75t_L g4611 ( 
.A1(n_4300),
.A2(n_3921),
.B(n_3919),
.Y(n_4611)
);

OAI22xp5_ASAP7_75t_L g4612 ( 
.A1(n_4247),
.A2(n_3952),
.B1(n_3962),
.B2(n_3942),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4346),
.B(n_3952),
.Y(n_4613)
);

AND2x4_ASAP7_75t_L g4614 ( 
.A(n_4350),
.B(n_3962),
.Y(n_4614)
);

BUFx6f_ASAP7_75t_L g4615 ( 
.A(n_4288),
.Y(n_4615)
);

AOI22xp33_ASAP7_75t_SL g4616 ( 
.A1(n_4456),
.A2(n_3986),
.B1(n_4014),
.B2(n_3966),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4321),
.Y(n_4617)
);

BUFx4_ASAP7_75t_SL g4618 ( 
.A(n_4453),
.Y(n_4618)
);

AND2x4_ASAP7_75t_L g4619 ( 
.A(n_4414),
.B(n_3966),
.Y(n_4619)
);

AOI22xp33_ASAP7_75t_L g4620 ( 
.A1(n_4304),
.A2(n_4359),
.B1(n_4260),
.B2(n_4467),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4397),
.Y(n_4621)
);

INVx3_ASAP7_75t_L g4622 ( 
.A(n_4263),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4277),
.B(n_3986),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4383),
.B(n_4014),
.Y(n_4624)
);

OAI21x1_ASAP7_75t_L g4625 ( 
.A1(n_4272),
.A2(n_4283),
.B(n_4229),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_4408),
.Y(n_4626)
);

NAND2xp33_ASAP7_75t_L g4627 ( 
.A(n_4471),
.B(n_4025),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_L g4628 ( 
.A(n_4440),
.B(n_4025),
.Y(n_4628)
);

BUFx3_ASAP7_75t_L g4629 ( 
.A(n_4250),
.Y(n_4629)
);

OR2x2_ASAP7_75t_L g4630 ( 
.A(n_4476),
.B(n_4045),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4449),
.B(n_4045),
.Y(n_4631)
);

AND2x4_ASAP7_75t_L g4632 ( 
.A(n_4434),
.B(n_4047),
.Y(n_4632)
);

AO32x1_ASAP7_75t_L g4633 ( 
.A1(n_4508),
.A2(n_4070),
.A3(n_4077),
.B1(n_4051),
.B2(n_4047),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_L g4634 ( 
.A(n_4491),
.B(n_524),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4338),
.B(n_4051),
.Y(n_4635)
);

HB1xp67_ASAP7_75t_L g4636 ( 
.A(n_4375),
.Y(n_4636)
);

BUFx3_ASAP7_75t_L g4637 ( 
.A(n_4368),
.Y(n_4637)
);

AOI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_4302),
.A2(n_4077),
.B(n_4070),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4312),
.A2(n_4084),
.B(n_525),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4422),
.Y(n_4640)
);

INVx3_ASAP7_75t_L g4641 ( 
.A(n_4490),
.Y(n_4641)
);

HB1xp67_ASAP7_75t_L g4642 ( 
.A(n_4388),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4504),
.B(n_4084),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4291),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4243),
.B(n_525),
.Y(n_4645)
);

OAI22xp5_ASAP7_75t_L g4646 ( 
.A1(n_4255),
.A2(n_528),
.B1(n_526),
.B2(n_527),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4334),
.B(n_949),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4289),
.Y(n_4648)
);

AND2x4_ASAP7_75t_L g4649 ( 
.A(n_4450),
.B(n_528),
.Y(n_4649)
);

OR2x6_ASAP7_75t_L g4650 ( 
.A(n_4483),
.B(n_4465),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4245),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4388),
.Y(n_4652)
);

BUFx2_ASAP7_75t_L g4653 ( 
.A(n_4510),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4236),
.B(n_529),
.Y(n_4654)
);

BUFx2_ASAP7_75t_L g4655 ( 
.A(n_4389),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4276),
.B(n_952),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4242),
.Y(n_4657)
);

BUFx6f_ASAP7_75t_L g4658 ( 
.A(n_4311),
.Y(n_4658)
);

INVx5_ASAP7_75t_L g4659 ( 
.A(n_4416),
.Y(n_4659)
);

OAI22xp5_ASAP7_75t_L g4660 ( 
.A1(n_4462),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4395),
.Y(n_4661)
);

AND2x4_ASAP7_75t_L g4662 ( 
.A(n_4398),
.B(n_531),
.Y(n_4662)
);

INVx3_ASAP7_75t_L g4663 ( 
.A(n_4377),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4478),
.B(n_959),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4396),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4253),
.Y(n_4666)
);

OAI22xp33_ASAP7_75t_SL g4667 ( 
.A1(n_4489),
.A2(n_536),
.B1(n_533),
.B2(n_535),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4256),
.Y(n_4668)
);

NOR2xp33_ASAP7_75t_SL g4669 ( 
.A(n_4505),
.B(n_533),
.Y(n_4669)
);

AND2x4_ASAP7_75t_L g4670 ( 
.A(n_4391),
.B(n_535),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4230),
.B(n_967),
.Y(n_4671)
);

OR2x6_ASAP7_75t_L g4672 ( 
.A(n_4290),
.B(n_4469),
.Y(n_4672)
);

BUFx6f_ASAP7_75t_L g4673 ( 
.A(n_4443),
.Y(n_4673)
);

AOI22xp33_ASAP7_75t_L g4674 ( 
.A1(n_4309),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4425),
.B(n_941),
.Y(n_4675)
);

BUFx2_ASAP7_75t_L g4676 ( 
.A(n_4347),
.Y(n_4676)
);

AND2x4_ASAP7_75t_L g4677 ( 
.A(n_4401),
.B(n_538),
.Y(n_4677)
);

A2O1A1Ixp33_ASAP7_75t_L g4678 ( 
.A1(n_4473),
.A2(n_944),
.B(n_945),
.C(n_943),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4421),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4423),
.B(n_947),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4322),
.A2(n_539),
.B(n_542),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4269),
.Y(n_4682)
);

BUFx2_ASAP7_75t_L g4683 ( 
.A(n_4447),
.Y(n_4683)
);

CKINVDCx5p33_ASAP7_75t_R g4684 ( 
.A(n_4503),
.Y(n_4684)
);

INVx3_ASAP7_75t_SL g4685 ( 
.A(n_4445),
.Y(n_4685)
);

OAI22xp5_ASAP7_75t_L g4686 ( 
.A1(n_4506),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_4686)
);

OAI21x1_ASAP7_75t_L g4687 ( 
.A1(n_4238),
.A2(n_543),
.B(n_544),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4296),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4270),
.B(n_545),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4287),
.Y(n_4690)
);

NAND2x1p5_ASAP7_75t_L g4691 ( 
.A(n_4484),
.B(n_547),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4430),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4310),
.A2(n_547),
.B(n_548),
.Y(n_4693)
);

INVx3_ASAP7_75t_L g4694 ( 
.A(n_4442),
.Y(n_4694)
);

NOR2xp33_ASAP7_75t_L g4695 ( 
.A(n_4458),
.B(n_548),
.Y(n_4695)
);

OAI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4493),
.A2(n_549),
.B(n_550),
.Y(n_4696)
);

NAND2x1p5_ASAP7_75t_L g4697 ( 
.A(n_4444),
.B(n_549),
.Y(n_4697)
);

O2A1O1Ixp33_ASAP7_75t_L g4698 ( 
.A1(n_4345),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4363),
.B(n_4385),
.Y(n_4699)
);

INVx5_ASAP7_75t_L g4700 ( 
.A(n_4402),
.Y(n_4700)
);

OR2x6_ASAP7_75t_L g4701 ( 
.A(n_4441),
.B(n_553),
.Y(n_4701)
);

AOI21xp5_ASAP7_75t_L g4702 ( 
.A1(n_4305),
.A2(n_554),
.B(n_555),
.Y(n_4702)
);

INVx2_ASAP7_75t_SL g4703 ( 
.A(n_4459),
.Y(n_4703)
);

INVx2_ASAP7_75t_L g4704 ( 
.A(n_4294),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4349),
.B(n_554),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4286),
.A2(n_555),
.B(n_556),
.Y(n_4706)
);

NAND3xp33_ASAP7_75t_L g4707 ( 
.A(n_4492),
.B(n_556),
.C(n_557),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4303),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4432),
.Y(n_4709)
);

A2O1A1Ixp33_ASAP7_75t_L g4710 ( 
.A1(n_4610),
.A2(n_4512),
.B(n_4475),
.C(n_4497),
.Y(n_4710)
);

AOI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4586),
.A2(n_4499),
.B(n_4268),
.Y(n_4711)
);

AND2x4_ASAP7_75t_L g4712 ( 
.A(n_4542),
.B(n_4329),
.Y(n_4712)
);

OAI22xp5_ASAP7_75t_L g4713 ( 
.A1(n_4620),
.A2(n_4358),
.B1(n_4511),
.B2(n_4488),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4523),
.Y(n_4714)
);

A2O1A1Ixp33_ASAP7_75t_L g4715 ( 
.A1(n_4607),
.A2(n_4274),
.B(n_4426),
.C(n_4380),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4526),
.B(n_4455),
.Y(n_4716)
);

A2O1A1Ixp33_ASAP7_75t_L g4717 ( 
.A1(n_4521),
.A2(n_4460),
.B(n_4344),
.C(n_4265),
.Y(n_4717)
);

OA21x2_ASAP7_75t_L g4718 ( 
.A1(n_4603),
.A2(n_4326),
.B(n_4373),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4532),
.Y(n_4719)
);

NAND2x1p5_ASAP7_75t_L g4720 ( 
.A(n_4528),
.B(n_4448),
.Y(n_4720)
);

AOI21xp5_ASAP7_75t_L g4721 ( 
.A1(n_4633),
.A2(n_4281),
.B(n_4271),
.Y(n_4721)
);

AOI21xp5_ASAP7_75t_SL g4722 ( 
.A1(n_4612),
.A2(n_4513),
.B(n_4433),
.Y(n_4722)
);

A2O1A1Ixp33_ASAP7_75t_L g4723 ( 
.A1(n_4669),
.A2(n_4472),
.B(n_4454),
.C(n_4457),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_L g4724 ( 
.A(n_4666),
.B(n_4308),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4563),
.B(n_4406),
.Y(n_4725)
);

NAND2x1_ASAP7_75t_L g4726 ( 
.A(n_4529),
.B(n_4468),
.Y(n_4726)
);

AND2x4_ASAP7_75t_L g4727 ( 
.A(n_4546),
.B(n_4501),
.Y(n_4727)
);

NAND2xp33_ASAP7_75t_SL g4728 ( 
.A(n_4525),
.B(n_4446),
.Y(n_4728)
);

OAI22xp5_ASAP7_75t_L g4729 ( 
.A1(n_4533),
.A2(n_4452),
.B1(n_4367),
.B2(n_4384),
.Y(n_4729)
);

CKINVDCx16_ASAP7_75t_R g4730 ( 
.A(n_4520),
.Y(n_4730)
);

INVx2_ASAP7_75t_SL g4731 ( 
.A(n_4528),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4549),
.Y(n_4732)
);

NOR2xp67_ASAP7_75t_L g4733 ( 
.A(n_4700),
.B(n_4567),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4535),
.B(n_4494),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4527),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4545),
.B(n_4318),
.Y(n_4736)
);

A2O1A1Ixp33_ASAP7_75t_L g4737 ( 
.A1(n_4567),
.A2(n_4386),
.B(n_4267),
.C(n_4314),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4668),
.B(n_4320),
.Y(n_4738)
);

OR2x6_ASAP7_75t_SL g4739 ( 
.A(n_4534),
.B(n_4225),
.Y(n_4739)
);

BUFx3_ASAP7_75t_L g4740 ( 
.A(n_4571),
.Y(n_4740)
);

OR2x6_ASAP7_75t_SL g4741 ( 
.A(n_4626),
.B(n_4225),
.Y(n_4741)
);

A2O1A1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_4627),
.A2(n_4301),
.B(n_4428),
.C(n_4419),
.Y(n_4742)
);

NOR2xp67_ASAP7_75t_L g4743 ( 
.A(n_4700),
.B(n_4509),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4556),
.Y(n_4744)
);

OR2x2_ASAP7_75t_L g4745 ( 
.A(n_4538),
.B(n_4381),
.Y(n_4745)
);

INVx1_ASAP7_75t_SL g4746 ( 
.A(n_4517),
.Y(n_4746)
);

AND2x4_ASAP7_75t_L g4747 ( 
.A(n_4546),
.B(n_4501),
.Y(n_4747)
);

BUFx2_ASAP7_75t_L g4748 ( 
.A(n_4536),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4565),
.Y(n_4749)
);

INVx2_ASAP7_75t_SL g4750 ( 
.A(n_4561),
.Y(n_4750)
);

HB1xp67_ASAP7_75t_L g4751 ( 
.A(n_4636),
.Y(n_4751)
);

O2A1O1Ixp33_ASAP7_75t_L g4752 ( 
.A1(n_4547),
.A2(n_4266),
.B(n_4500),
.C(n_4474),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4676),
.B(n_4332),
.Y(n_4753)
);

NOR2x1_ASAP7_75t_SL g4754 ( 
.A(n_4579),
.B(n_4257),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4558),
.Y(n_4755)
);

NOR2x2_ASAP7_75t_L g4756 ( 
.A(n_4579),
.B(n_4447),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4573),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4566),
.Y(n_4758)
);

BUFx4f_ASAP7_75t_SL g4759 ( 
.A(n_4539),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4574),
.Y(n_4760)
);

AND2x4_ASAP7_75t_L g4761 ( 
.A(n_4531),
.B(n_4485),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4582),
.Y(n_4762)
);

AOI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4633),
.A2(n_4248),
.B(n_4235),
.Y(n_4763)
);

BUFx3_ASAP7_75t_L g4764 ( 
.A(n_4519),
.Y(n_4764)
);

AND2x4_ASAP7_75t_L g4765 ( 
.A(n_4637),
.B(n_4485),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_4594),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4682),
.B(n_4317),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_4602),
.Y(n_4768)
);

INVx1_ASAP7_75t_SL g4769 ( 
.A(n_4605),
.Y(n_4769)
);

AND2x4_ASAP7_75t_L g4770 ( 
.A(n_4553),
.B(n_4298),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4657),
.B(n_4413),
.Y(n_4771)
);

OR2x6_ASAP7_75t_SL g4772 ( 
.A(n_4684),
.B(n_4507),
.Y(n_4772)
);

AND2x4_ASAP7_75t_L g4773 ( 
.A(n_4595),
.B(n_4482),
.Y(n_4773)
);

BUFx6f_ASAP7_75t_L g4774 ( 
.A(n_4576),
.Y(n_4774)
);

HB1xp67_ASAP7_75t_L g4775 ( 
.A(n_4568),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4690),
.B(n_4317),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4704),
.B(n_4393),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4583),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4623),
.B(n_4482),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4540),
.A2(n_4355),
.B(n_4299),
.Y(n_4780)
);

OR2x6_ASAP7_75t_L g4781 ( 
.A(n_4650),
.B(n_4392),
.Y(n_4781)
);

O2A1O1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4593),
.A2(n_4378),
.B(n_4387),
.C(n_4429),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4584),
.Y(n_4783)
);

NOR2xp67_ASAP7_75t_L g4784 ( 
.A(n_4659),
.B(n_558),
.Y(n_4784)
);

HB1xp67_ASAP7_75t_L g4785 ( 
.A(n_4524),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4518),
.Y(n_4786)
);

A2O1A1Ixp33_ASAP7_75t_L g4787 ( 
.A1(n_4559),
.A2(n_4437),
.B(n_4480),
.C(n_4481),
.Y(n_4787)
);

NOR2xp67_ASAP7_75t_L g4788 ( 
.A(n_4659),
.B(n_558),
.Y(n_4788)
);

BUFx2_ASAP7_75t_L g4789 ( 
.A(n_4589),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4621),
.Y(n_4790)
);

INVx3_ASAP7_75t_L g4791 ( 
.A(n_4578),
.Y(n_4791)
);

OR2x6_ASAP7_75t_L g4792 ( 
.A(n_4650),
.B(n_4487),
.Y(n_4792)
);

CKINVDCx12_ASAP7_75t_R g4793 ( 
.A(n_4551),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4640),
.Y(n_4794)
);

AND2x4_ASAP7_75t_L g4795 ( 
.A(n_4614),
.B(n_4348),
.Y(n_4795)
);

OR2x2_ASAP7_75t_L g4796 ( 
.A(n_4708),
.B(n_4436),
.Y(n_4796)
);

AOI21x1_ASAP7_75t_SL g4797 ( 
.A1(n_4680),
.A2(n_4438),
.B(n_4362),
.Y(n_4797)
);

AND2x2_ASAP7_75t_SL g4798 ( 
.A(n_4683),
.B(n_4399),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_SL g4799 ( 
.A1(n_4677),
.A2(n_4399),
.B(n_4390),
.Y(n_4799)
);

OAI22xp5_ASAP7_75t_L g4800 ( 
.A1(n_4616),
.A2(n_4356),
.B1(n_4376),
.B2(n_4327),
.Y(n_4800)
);

BUFx3_ASAP7_75t_L g4801 ( 
.A(n_4555),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4643),
.B(n_4379),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4653),
.Y(n_4803)
);

OAI22xp5_ASAP7_75t_SL g4804 ( 
.A1(n_4629),
.A2(n_4240),
.B1(n_4405),
.B2(n_4404),
.Y(n_4804)
);

AND2x4_ASAP7_75t_L g4805 ( 
.A(n_4570),
.B(n_4364),
.Y(n_4805)
);

O2A1O1Ixp33_ASAP7_75t_L g4806 ( 
.A1(n_4646),
.A2(n_4705),
.B(n_4654),
.C(n_4667),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4613),
.B(n_4548),
.Y(n_4807)
);

AOI21xp5_ASAP7_75t_L g4808 ( 
.A1(n_4611),
.A2(n_4264),
.B(n_4282),
.Y(n_4808)
);

OAI31xp33_ASAP7_75t_L g4809 ( 
.A1(n_4599),
.A2(n_4410),
.A3(n_561),
.B(n_559),
.Y(n_4809)
);

INVx2_ASAP7_75t_L g4810 ( 
.A(n_4651),
.Y(n_4810)
);

INVxp67_ASAP7_75t_L g4811 ( 
.A(n_4557),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4596),
.Y(n_4812)
);

INVx1_ASAP7_75t_SL g4813 ( 
.A(n_4555),
.Y(n_4813)
);

AOI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4638),
.A2(n_4343),
.B(n_4339),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4648),
.B(n_4240),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4699),
.B(n_4530),
.Y(n_4816)
);

OR2x2_ASAP7_75t_L g4817 ( 
.A(n_4572),
.B(n_560),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4554),
.B(n_4407),
.Y(n_4818)
);

A2O1A1Ixp33_ASAP7_75t_L g4819 ( 
.A1(n_4698),
.A2(n_4435),
.B(n_4424),
.C(n_563),
.Y(n_4819)
);

A2O1A1Ixp33_ASAP7_75t_SL g4820 ( 
.A1(n_4695),
.A2(n_563),
.B(n_560),
.C(n_562),
.Y(n_4820)
);

A2O1A1Ixp33_ASAP7_75t_SL g4821 ( 
.A1(n_4585),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4661),
.B(n_564),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4665),
.B(n_4569),
.Y(n_4823)
);

NOR2xp67_ASAP7_75t_L g4824 ( 
.A(n_4522),
.B(n_565),
.Y(n_4824)
);

A2O1A1Ixp33_ASAP7_75t_L g4825 ( 
.A1(n_4543),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_4825)
);

AOI21xp5_ASAP7_75t_SL g4826 ( 
.A1(n_4662),
.A2(n_569),
.B(n_570),
.Y(n_4826)
);

O2A1O1Ixp5_ASAP7_75t_L g4827 ( 
.A1(n_4537),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_4827)
);

CKINVDCx5p33_ASAP7_75t_R g4828 ( 
.A(n_4606),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4735),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4749),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4757),
.Y(n_4831)
);

OAI21x1_ASAP7_75t_L g4832 ( 
.A1(n_4763),
.A2(n_4587),
.B(n_4625),
.Y(n_4832)
);

HB1xp67_ASAP7_75t_L g4833 ( 
.A(n_4751),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4789),
.Y(n_4834)
);

INVx2_ASAP7_75t_SL g4835 ( 
.A(n_4740),
.Y(n_4835)
);

OR2x6_ASAP7_75t_L g4836 ( 
.A(n_4733),
.B(n_4672),
.Y(n_4836)
);

INVx2_ASAP7_75t_L g4837 ( 
.A(n_4714),
.Y(n_4837)
);

NAND2x1p5_ASAP7_75t_L g4838 ( 
.A(n_4731),
.B(n_4576),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4762),
.Y(n_4839)
);

OAI21x1_ASAP7_75t_L g4840 ( 
.A1(n_4814),
.A2(n_4652),
.B(n_4694),
.Y(n_4840)
);

INVx2_ASAP7_75t_L g4841 ( 
.A(n_4719),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4778),
.Y(n_4842)
);

CKINVDCx20_ASAP7_75t_R g4843 ( 
.A(n_4730),
.Y(n_4843)
);

HB1xp67_ASAP7_75t_L g4844 ( 
.A(n_4775),
.Y(n_4844)
);

INVx3_ASAP7_75t_L g4845 ( 
.A(n_4761),
.Y(n_4845)
);

INVx2_ASAP7_75t_L g4846 ( 
.A(n_4744),
.Y(n_4846)
);

OAI22xp5_ASAP7_75t_L g4847 ( 
.A1(n_4739),
.A2(n_4741),
.B1(n_4772),
.B2(n_4824),
.Y(n_4847)
);

NOR2xp67_ASAP7_75t_L g4848 ( 
.A(n_4791),
.B(n_4560),
.Y(n_4848)
);

BUFx2_ASAP7_75t_L g4849 ( 
.A(n_4748),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4783),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4755),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4758),
.Y(n_4852)
);

AOI22xp33_ASAP7_75t_L g4853 ( 
.A1(n_4713),
.A2(n_4673),
.B1(n_4552),
.B2(n_4655),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4812),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4750),
.Y(n_4855)
);

OR2x2_ASAP7_75t_L g4856 ( 
.A(n_4785),
.B(n_4736),
.Y(n_4856)
);

INVx3_ASAP7_75t_L g4857 ( 
.A(n_4770),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4794),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4810),
.Y(n_4859)
);

BUFx2_ASAP7_75t_L g4860 ( 
.A(n_4764),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4760),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4745),
.Y(n_4862)
);

AOI21xp5_ASAP7_75t_L g4863 ( 
.A1(n_4754),
.A2(n_4550),
.B(n_4588),
.Y(n_4863)
);

OAI21x1_ASAP7_75t_L g4864 ( 
.A1(n_4721),
.A2(n_4642),
.B(n_4600),
.Y(n_4864)
);

BUFx3_ASAP7_75t_L g4865 ( 
.A(n_4828),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4732),
.Y(n_4866)
);

AOI21x1_ASAP7_75t_L g4867 ( 
.A1(n_4780),
.A2(n_4672),
.B(n_4580),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4766),
.Y(n_4868)
);

BUFx3_ASAP7_75t_L g4869 ( 
.A(n_4759),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4773),
.Y(n_4870)
);

AND2x4_ASAP7_75t_L g4871 ( 
.A(n_4765),
.B(n_4692),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4790),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4786),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_4802),
.B(n_4663),
.Y(n_4874)
);

INVx1_ASAP7_75t_SL g4875 ( 
.A(n_4769),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4753),
.Y(n_4876)
);

BUFx3_ASAP7_75t_L g4877 ( 
.A(n_4801),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4767),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4793),
.B(n_4608),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4776),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4823),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4724),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4803),
.Y(n_4883)
);

OR2x2_ASAP7_75t_L g4884 ( 
.A(n_4816),
.B(n_4815),
.Y(n_4884)
);

AOI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_4800),
.A2(n_4673),
.B1(n_4516),
.B2(n_4707),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4738),
.Y(n_4886)
);

BUFx2_ASAP7_75t_L g4887 ( 
.A(n_4774),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4734),
.B(n_4590),
.Y(n_4888)
);

AND2x2_ASAP7_75t_L g4889 ( 
.A(n_4807),
.B(n_4631),
.Y(n_4889)
);

OAI21x1_ASAP7_75t_L g4890 ( 
.A1(n_4808),
.A2(n_4688),
.B(n_4617),
.Y(n_4890)
);

AO21x2_ASAP7_75t_L g4891 ( 
.A1(n_4777),
.A2(n_4696),
.B(n_4689),
.Y(n_4891)
);

OR2x6_ASAP7_75t_L g4892 ( 
.A(n_4781),
.B(n_4598),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4796),
.Y(n_4893)
);

AO21x2_ASAP7_75t_L g4894 ( 
.A1(n_4784),
.A2(n_4706),
.B(n_4664),
.Y(n_4894)
);

OAI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_4737),
.A2(n_4685),
.B1(n_4641),
.B2(n_4701),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4771),
.Y(n_4896)
);

INVxp67_ASAP7_75t_L g4897 ( 
.A(n_4746),
.Y(n_4897)
);

OAI21xp5_ASAP7_75t_L g4898 ( 
.A1(n_4715),
.A2(n_4678),
.B(n_4679),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4798),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4712),
.Y(n_4900)
);

BUFx2_ASAP7_75t_L g4901 ( 
.A(n_4774),
.Y(n_4901)
);

OAI21xp5_ASAP7_75t_L g4902 ( 
.A1(n_4825),
.A2(n_4687),
.B(n_4701),
.Y(n_4902)
);

HB1xp67_ASAP7_75t_SL g4903 ( 
.A(n_4727),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4779),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4718),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4718),
.Y(n_4906)
);

BUFx3_ASAP7_75t_L g4907 ( 
.A(n_4768),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_SL g4908 ( 
.A(n_4747),
.B(n_4615),
.Y(n_4908)
);

INVxp67_ASAP7_75t_L g4909 ( 
.A(n_4725),
.Y(n_4909)
);

INVx3_ASAP7_75t_L g4910 ( 
.A(n_4781),
.Y(n_4910)
);

OAI21x1_ASAP7_75t_L g4911 ( 
.A1(n_4726),
.A2(n_4797),
.B(n_4711),
.Y(n_4911)
);

AOI22xp33_ASAP7_75t_L g4912 ( 
.A1(n_4792),
.A2(n_4703),
.B1(n_4656),
.B2(n_4686),
.Y(n_4912)
);

OR2x2_ASAP7_75t_L g4913 ( 
.A(n_4716),
.B(n_4635),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4818),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4805),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4817),
.Y(n_4916)
);

BUFx3_ASAP7_75t_L g4917 ( 
.A(n_4813),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4795),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4756),
.Y(n_4919)
);

INVx2_ASAP7_75t_L g4920 ( 
.A(n_4720),
.Y(n_4920)
);

AO21x2_ASAP7_75t_L g4921 ( 
.A1(n_4788),
.A2(n_4709),
.B(n_4634),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4878),
.Y(n_4922)
);

OAI21xp33_ASAP7_75t_L g4923 ( 
.A1(n_4919),
.A2(n_4717),
.B(n_4722),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4880),
.B(n_4884),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4849),
.Y(n_4925)
);

HB1xp67_ASAP7_75t_L g4926 ( 
.A(n_4833),
.Y(n_4926)
);

NOR2x1_ASAP7_75t_SL g4927 ( 
.A(n_4836),
.B(n_4792),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4874),
.B(n_4811),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4844),
.Y(n_4929)
);

INVx3_ASAP7_75t_L g4930 ( 
.A(n_4836),
.Y(n_4930)
);

BUFx8_ASAP7_75t_L g4931 ( 
.A(n_4860),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4854),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4866),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4900),
.B(n_4619),
.Y(n_4934)
);

INVx2_ASAP7_75t_SL g4935 ( 
.A(n_4835),
.Y(n_4935)
);

BUFx6f_ASAP7_75t_L g4936 ( 
.A(n_4865),
.Y(n_4936)
);

OR2x2_ASAP7_75t_L g4937 ( 
.A(n_4856),
.B(n_4592),
.Y(n_4937)
);

INVx2_ASAP7_75t_L g4938 ( 
.A(n_4837),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4900),
.B(n_4597),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4914),
.B(n_4743),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4889),
.B(n_4601),
.Y(n_4941)
);

OAI211xp5_ASAP7_75t_SL g4942 ( 
.A1(n_4853),
.A2(n_4885),
.B(n_4912),
.C(n_4847),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4873),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4881),
.B(n_4729),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4904),
.B(n_4564),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4841),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4845),
.B(n_4615),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4845),
.B(n_4630),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4882),
.B(n_4544),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4834),
.B(n_4577),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4829),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4859),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4846),
.Y(n_4953)
);

OAI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4903),
.A2(n_4826),
.B1(n_4723),
.B2(n_4591),
.Y(n_4954)
);

INVx2_ASAP7_75t_L g4955 ( 
.A(n_4851),
.Y(n_4955)
);

AND2x2_ASAP7_75t_L g4956 ( 
.A(n_4909),
.B(n_4644),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4886),
.B(n_4782),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4871),
.B(n_4624),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4852),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4861),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4871),
.B(n_4870),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4870),
.B(n_4857),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4868),
.Y(n_4963)
);

INVx2_ASAP7_75t_L g4964 ( 
.A(n_4872),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4857),
.B(n_4575),
.Y(n_4965)
);

INVx2_ASAP7_75t_L g4966 ( 
.A(n_4883),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4862),
.B(n_4822),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4830),
.Y(n_4968)
);

BUFx2_ASAP7_75t_L g4969 ( 
.A(n_4855),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_L g4970 ( 
.A(n_4876),
.B(n_4541),
.Y(n_4970)
);

NOR2x1p5_ASAP7_75t_L g4971 ( 
.A(n_4910),
.B(n_4899),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4831),
.Y(n_4972)
);

HB1xp67_ASAP7_75t_L g4973 ( 
.A(n_4848),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4839),
.Y(n_4974)
);

HB1xp67_ASAP7_75t_L g4975 ( 
.A(n_4907),
.Y(n_4975)
);

AND2x2_ASAP7_75t_L g4976 ( 
.A(n_4910),
.B(n_4632),
.Y(n_4976)
);

HB1xp67_ASAP7_75t_L g4977 ( 
.A(n_4875),
.Y(n_4977)
);

AOI22xp33_ASAP7_75t_L g4978 ( 
.A1(n_4898),
.A2(n_4728),
.B1(n_4804),
.B2(n_4809),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4918),
.B(n_4675),
.Y(n_4979)
);

INVxp33_ASAP7_75t_L g4980 ( 
.A(n_4879),
.Y(n_4980)
);

INVx3_ASAP7_75t_L g4981 ( 
.A(n_4892),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4842),
.Y(n_4982)
);

BUFx3_ASAP7_75t_L g4983 ( 
.A(n_4843),
.Y(n_4983)
);

INVxp67_ASAP7_75t_L g4984 ( 
.A(n_4917),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4850),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4893),
.B(n_4609),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4915),
.B(n_4647),
.Y(n_4987)
);

INVx2_ASAP7_75t_L g4988 ( 
.A(n_4905),
.Y(n_4988)
);

BUFx6f_ASAP7_75t_L g4989 ( 
.A(n_4869),
.Y(n_4989)
);

INVx5_ASAP7_75t_L g4990 ( 
.A(n_4892),
.Y(n_4990)
);

INVxp67_ASAP7_75t_SL g4991 ( 
.A(n_4897),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4915),
.B(n_4671),
.Y(n_4992)
);

INVxp67_ASAP7_75t_L g4993 ( 
.A(n_4877),
.Y(n_4993)
);

AND2x4_ASAP7_75t_L g4994 ( 
.A(n_4920),
.B(n_4581),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4896),
.B(n_4628),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_4905),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4888),
.B(n_4658),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4913),
.B(n_4658),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4858),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4906),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4916),
.B(n_4787),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4906),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4890),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4864),
.Y(n_5004)
);

AND2x4_ASAP7_75t_L g5005 ( 
.A(n_4927),
.B(n_4899),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4969),
.Y(n_5006)
);

INVx4_ASAP7_75t_L g5007 ( 
.A(n_4989),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4932),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4932),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4926),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4922),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4922),
.B(n_4891),
.Y(n_5012)
);

INVx2_ASAP7_75t_SL g5013 ( 
.A(n_4931),
.Y(n_5013)
);

HB1xp67_ASAP7_75t_L g5014 ( 
.A(n_4988),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4972),
.Y(n_5015)
);

INVx3_ASAP7_75t_L g5016 ( 
.A(n_4931),
.Y(n_5016)
);

AOI22xp33_ASAP7_75t_L g5017 ( 
.A1(n_4942),
.A2(n_4895),
.B1(n_4894),
.B2(n_4921),
.Y(n_5017)
);

AND2x2_ASAP7_75t_L g5018 ( 
.A(n_4961),
.B(n_4887),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4962),
.B(n_4901),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_5001),
.B(n_4911),
.Y(n_5020)
);

INVx2_ASAP7_75t_SL g5021 ( 
.A(n_4936),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4972),
.Y(n_5022)
);

OAI211xp5_ASAP7_75t_L g5023 ( 
.A1(n_4978),
.A2(n_4902),
.B(n_4752),
.C(n_4867),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4930),
.B(n_4908),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4930),
.B(n_4867),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4985),
.Y(n_5026)
);

BUFx2_ASAP7_75t_L g5027 ( 
.A(n_4975),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4985),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_4996),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4999),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4999),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4957),
.B(n_4863),
.Y(n_5032)
);

INVx2_ASAP7_75t_L g5033 ( 
.A(n_4953),
.Y(n_5033)
);

BUFx3_ASAP7_75t_L g5034 ( 
.A(n_4983),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_4953),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_4960),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_4973),
.B(n_4838),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4924),
.Y(n_5038)
);

INVx2_ASAP7_75t_L g5039 ( 
.A(n_4960),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_4963),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4965),
.B(n_4840),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4952),
.B(n_4951),
.Y(n_5042)
);

OR2x2_ASAP7_75t_L g5043 ( 
.A(n_4937),
.B(n_4832),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4952),
.B(n_4799),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4940),
.B(n_4622),
.Y(n_5045)
);

OR2x2_ASAP7_75t_L g5046 ( 
.A(n_4949),
.B(n_4645),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4971),
.B(n_4977),
.Y(n_5047)
);

AOI22xp33_ASAP7_75t_L g5048 ( 
.A1(n_4923),
.A2(n_4649),
.B1(n_4670),
.B2(n_4639),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4963),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_5000),
.B(n_4819),
.Y(n_5050)
);

OAI221xp5_ASAP7_75t_L g5051 ( 
.A1(n_4954),
.A2(n_4991),
.B1(n_4944),
.B2(n_4981),
.C(n_4984),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4947),
.B(n_4976),
.Y(n_5052)
);

OAI31xp33_ASAP7_75t_L g5053 ( 
.A1(n_4981),
.A2(n_4710),
.A3(n_4821),
.B(n_4820),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_4997),
.B(n_4581),
.Y(n_5054)
);

HB1xp67_ASAP7_75t_L g5055 ( 
.A(n_5000),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4948),
.B(n_4742),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_5005),
.B(n_4980),
.Y(n_5057)
);

OR2x2_ASAP7_75t_L g5058 ( 
.A(n_5050),
.B(n_4929),
.Y(n_5058)
);

AND2x4_ASAP7_75t_L g5059 ( 
.A(n_5005),
.B(n_4990),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_5047),
.B(n_4956),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_5050),
.B(n_4933),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_5037),
.B(n_5024),
.Y(n_5062)
);

INVx2_ASAP7_75t_SL g5063 ( 
.A(n_5016),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5027),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_5032),
.B(n_4943),
.Y(n_5065)
);

BUFx3_ASAP7_75t_L g5066 ( 
.A(n_5016),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_5056),
.B(n_4993),
.Y(n_5067)
);

AND2x4_ASAP7_75t_L g5068 ( 
.A(n_5007),
.B(n_4990),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_5014),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_5041),
.B(n_4925),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_5032),
.B(n_4968),
.Y(n_5071)
);

INVxp67_ASAP7_75t_L g5072 ( 
.A(n_5034),
.Y(n_5072)
);

AND2x4_ASAP7_75t_L g5073 ( 
.A(n_5007),
.B(n_4990),
.Y(n_5073)
);

HB1xp67_ASAP7_75t_L g5074 ( 
.A(n_5010),
.Y(n_5074)
);

AOI22xp33_ASAP7_75t_L g5075 ( 
.A1(n_5051),
.A2(n_4989),
.B1(n_4934),
.B2(n_4939),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_5006),
.B(n_4935),
.Y(n_5076)
);

OR2x2_ASAP7_75t_L g5077 ( 
.A(n_5038),
.B(n_5002),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_5042),
.Y(n_5078)
);

BUFx3_ASAP7_75t_L g5079 ( 
.A(n_5013),
.Y(n_5079)
);

AND2x2_ASAP7_75t_L g5080 ( 
.A(n_5021),
.B(n_4998),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_5025),
.B(n_4958),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_5042),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5011),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5055),
.Y(n_5084)
);

BUFx2_ASAP7_75t_L g5085 ( 
.A(n_5054),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_5017),
.B(n_4974),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_5055),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_5019),
.B(n_4941),
.Y(n_5088)
);

AND2x4_ASAP7_75t_L g5089 ( 
.A(n_5045),
.B(n_4989),
.Y(n_5089)
);

OR2x2_ASAP7_75t_L g5090 ( 
.A(n_5012),
.B(n_5002),
.Y(n_5090)
);

HB1xp67_ASAP7_75t_L g5091 ( 
.A(n_5014),
.Y(n_5091)
);

INVx4_ASAP7_75t_L g5092 ( 
.A(n_5018),
.Y(n_5092)
);

NOR2xp67_ASAP7_75t_L g5093 ( 
.A(n_5023),
.B(n_5004),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_5015),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_5029),
.Y(n_5095)
);

AND2x2_ASAP7_75t_L g5096 ( 
.A(n_5052),
.B(n_5043),
.Y(n_5096)
);

AND2x2_ASAP7_75t_L g5097 ( 
.A(n_5020),
.B(n_4994),
.Y(n_5097)
);

NOR2xp33_ASAP7_75t_SL g5098 ( 
.A(n_5051),
.B(n_4936),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5022),
.Y(n_5099)
);

AND2x4_ASAP7_75t_L g5100 ( 
.A(n_5044),
.B(n_4936),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5026),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_5020),
.B(n_4994),
.Y(n_5102)
);

NOR2xp33_ASAP7_75t_L g5103 ( 
.A(n_5023),
.B(n_4967),
.Y(n_5103)
);

AND2x4_ASAP7_75t_L g5104 ( 
.A(n_5044),
.B(n_4928),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5028),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_5012),
.B(n_4982),
.Y(n_5106)
);

AND2x4_ASAP7_75t_L g5107 ( 
.A(n_5030),
.B(n_5003),
.Y(n_5107)
);

HB1xp67_ASAP7_75t_L g5108 ( 
.A(n_5008),
.Y(n_5108)
);

INVx3_ASAP7_75t_L g5109 ( 
.A(n_5033),
.Y(n_5109)
);

BUFx2_ASAP7_75t_L g5110 ( 
.A(n_5035),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5031),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_5009),
.B(n_4950),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_5046),
.B(n_4995),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_5036),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_5039),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_5071),
.Y(n_5116)
);

OAI33xp33_ASAP7_75t_L g5117 ( 
.A1(n_5064),
.A2(n_4970),
.A3(n_4986),
.B1(n_4806),
.B2(n_4660),
.B3(n_4562),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5065),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_5066),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_5079),
.B(n_4604),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_5063),
.Y(n_5121)
);

INVxp33_ASAP7_75t_L g5122 ( 
.A(n_5098),
.Y(n_5122)
);

AND2x2_ASAP7_75t_L g5123 ( 
.A(n_5057),
.B(n_4945),
.Y(n_5123)
);

INVx2_ASAP7_75t_L g5124 ( 
.A(n_5109),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_5058),
.Y(n_5125)
);

BUFx2_ASAP7_75t_L g5126 ( 
.A(n_5100),
.Y(n_5126)
);

OAI211xp5_ASAP7_75t_L g5127 ( 
.A1(n_5103),
.A2(n_5053),
.B(n_5048),
.C(n_4674),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5074),
.Y(n_5128)
);

AO21x2_ASAP7_75t_L g5129 ( 
.A1(n_5093),
.A2(n_5049),
.B(n_5040),
.Y(n_5129)
);

HB1xp67_ASAP7_75t_L g5130 ( 
.A(n_5091),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_5077),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_5110),
.Y(n_5132)
);

AND2x4_ASAP7_75t_L g5133 ( 
.A(n_5072),
.B(n_4979),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_5061),
.B(n_5053),
.Y(n_5134)
);

INVx2_ASAP7_75t_L g5135 ( 
.A(n_5069),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5108),
.Y(n_5136)
);

AOI211xp5_ASAP7_75t_L g5137 ( 
.A1(n_5059),
.A2(n_5073),
.B(n_5068),
.C(n_5100),
.Y(n_5137)
);

BUFx6f_ASAP7_75t_L g5138 ( 
.A(n_5068),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_5113),
.Y(n_5139)
);

HB1xp67_ASAP7_75t_L g5140 ( 
.A(n_5084),
.Y(n_5140)
);

OAI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_5075),
.A2(n_4987),
.B1(n_4992),
.B2(n_4966),
.Y(n_5141)
);

OAI21x1_ASAP7_75t_SL g5142 ( 
.A1(n_5092),
.A2(n_4618),
.B(n_4938),
.Y(n_5142)
);

INVx4_ASAP7_75t_L g5143 ( 
.A(n_5089),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_5078),
.B(n_4946),
.Y(n_5144)
);

AOI31xp67_ASAP7_75t_L g5145 ( 
.A1(n_5086),
.A2(n_4959),
.A3(n_4964),
.B(n_4955),
.Y(n_5145)
);

OAI22xp5_ASAP7_75t_L g5146 ( 
.A1(n_5059),
.A2(n_5062),
.B1(n_5104),
.B2(n_5085),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_5087),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_5082),
.B(n_5104),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_5095),
.Y(n_5149)
);

INVx2_ASAP7_75t_L g5150 ( 
.A(n_5076),
.Y(n_5150)
);

AND2x2_ASAP7_75t_L g5151 ( 
.A(n_5089),
.B(n_5097),
.Y(n_5151)
);

AND2x2_ASAP7_75t_L g5152 ( 
.A(n_5102),
.B(n_4697),
.Y(n_5152)
);

AOI222xp33_ASAP7_75t_L g5153 ( 
.A1(n_5067),
.A2(n_4827),
.B1(n_4691),
.B2(n_4702),
.C1(n_4681),
.C2(n_4693),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_5112),
.Y(n_5154)
);

INVxp67_ASAP7_75t_L g5155 ( 
.A(n_5073),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_5114),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5083),
.Y(n_5157)
);

NOR2xp33_ASAP7_75t_L g5158 ( 
.A(n_5088),
.B(n_571),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5094),
.Y(n_5159)
);

NAND3xp33_ASAP7_75t_L g5160 ( 
.A(n_5090),
.B(n_573),
.C(n_574),
.Y(n_5160)
);

NOR3xp33_ASAP7_75t_L g5161 ( 
.A(n_5106),
.B(n_5096),
.C(n_5099),
.Y(n_5161)
);

OR2x2_ASAP7_75t_L g5162 ( 
.A(n_5101),
.B(n_573),
.Y(n_5162)
);

HB1xp67_ASAP7_75t_L g5163 ( 
.A(n_5105),
.Y(n_5163)
);

BUFx3_ASAP7_75t_L g5164 ( 
.A(n_5080),
.Y(n_5164)
);

AOI222xp33_ASAP7_75t_L g5165 ( 
.A1(n_5111),
.A2(n_579),
.B1(n_581),
.B2(n_575),
.C1(n_577),
.C2(n_580),
.Y(n_5165)
);

INVx4_ASAP7_75t_L g5166 ( 
.A(n_5070),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_5081),
.A2(n_580),
.B1(n_575),
.B2(n_579),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5115),
.Y(n_5168)
);

BUFx3_ASAP7_75t_L g5169 ( 
.A(n_5107),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5060),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_SL g5171 ( 
.A1(n_5107),
.A2(n_581),
.B(n_583),
.Y(n_5171)
);

INVx3_ASAP7_75t_L g5172 ( 
.A(n_5079),
.Y(n_5172)
);

AO21x2_ASAP7_75t_L g5173 ( 
.A1(n_5093),
.A2(n_583),
.B(n_584),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_5071),
.Y(n_5174)
);

OR2x2_ASAP7_75t_L g5175 ( 
.A(n_5061),
.B(n_584),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_5071),
.Y(n_5176)
);

OA21x2_ASAP7_75t_L g5177 ( 
.A1(n_5072),
.A2(n_585),
.B(n_586),
.Y(n_5177)
);

AND2x2_ASAP7_75t_L g5178 ( 
.A(n_5057),
.B(n_587),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_5075),
.A2(n_590),
.B1(n_587),
.B2(n_588),
.Y(n_5179)
);

AOI21x1_ASAP7_75t_L g5180 ( 
.A1(n_5059),
.A2(n_964),
.B(n_590),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_5066),
.Y(n_5181)
);

OAI21x1_ASAP7_75t_L g5182 ( 
.A1(n_5091),
.A2(n_591),
.B(n_593),
.Y(n_5182)
);

INVx2_ASAP7_75t_L g5183 ( 
.A(n_5066),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_5057),
.B(n_591),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_5071),
.Y(n_5185)
);

O2A1O1Ixp33_ASAP7_75t_SL g5186 ( 
.A1(n_5063),
.A2(n_595),
.B(n_593),
.C(n_594),
.Y(n_5186)
);

AND2x6_ASAP7_75t_L g5187 ( 
.A(n_5066),
.B(n_594),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_5172),
.B(n_964),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5130),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_5128),
.Y(n_5190)
);

HB1xp67_ASAP7_75t_L g5191 ( 
.A(n_5135),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5119),
.B(n_5181),
.Y(n_5192)
);

OR2x2_ASAP7_75t_L g5193 ( 
.A(n_5139),
.B(n_595),
.Y(n_5193)
);

INVx2_ASAP7_75t_SL g5194 ( 
.A(n_5183),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5125),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_5140),
.Y(n_5196)
);

AND2x2_ASAP7_75t_L g5197 ( 
.A(n_5151),
.B(n_5122),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_5121),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5148),
.Y(n_5199)
);

OR2x2_ASAP7_75t_L g5200 ( 
.A(n_5116),
.B(n_962),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5163),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_5164),
.B(n_596),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5136),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5174),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_5176),
.B(n_596),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5185),
.Y(n_5206)
);

CKINVDCx16_ASAP7_75t_R g5207 ( 
.A(n_5120),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5118),
.B(n_5170),
.Y(n_5208)
);

NAND2x1p5_ASAP7_75t_L g5209 ( 
.A(n_5177),
.B(n_597),
.Y(n_5209)
);

AOI22xp33_ASAP7_75t_L g5210 ( 
.A1(n_5161),
.A2(n_601),
.B1(n_598),
.B2(n_599),
.Y(n_5210)
);

INVx2_ASAP7_75t_SL g5211 ( 
.A(n_5138),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_5134),
.B(n_598),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_5127),
.B(n_957),
.Y(n_5213)
);

NAND2xp5_ASAP7_75t_L g5214 ( 
.A(n_5131),
.B(n_957),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_5180),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_5132),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5126),
.Y(n_5217)
);

BUFx3_ASAP7_75t_L g5218 ( 
.A(n_5138),
.Y(n_5218)
);

NAND2x1_ASAP7_75t_L g5219 ( 
.A(n_5142),
.B(n_599),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5126),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5177),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_5155),
.B(n_955),
.Y(n_5222)
);

INVx1_ASAP7_75t_SL g5223 ( 
.A(n_5178),
.Y(n_5223)
);

AND2x2_ASAP7_75t_L g5224 ( 
.A(n_5143),
.B(n_601),
.Y(n_5224)
);

OR2x2_ASAP7_75t_L g5225 ( 
.A(n_5144),
.B(n_952),
.Y(n_5225)
);

AND2x2_ASAP7_75t_L g5226 ( 
.A(n_5166),
.B(n_602),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_5123),
.B(n_602),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5182),
.Y(n_5228)
);

OR2x6_ASAP7_75t_L g5229 ( 
.A(n_5142),
.B(n_603),
.Y(n_5229)
);

HB1xp67_ASAP7_75t_L g5230 ( 
.A(n_5149),
.Y(n_5230)
);

INVxp67_ASAP7_75t_SL g5231 ( 
.A(n_5184),
.Y(n_5231)
);

OR2x2_ASAP7_75t_L g5232 ( 
.A(n_5147),
.B(n_604),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5157),
.Y(n_5233)
);

AND2x4_ASAP7_75t_L g5234 ( 
.A(n_5150),
.B(n_604),
.Y(n_5234)
);

AND2x2_ASAP7_75t_L g5235 ( 
.A(n_5137),
.B(n_605),
.Y(n_5235)
);

AND2x2_ASAP7_75t_L g5236 ( 
.A(n_5152),
.B(n_605),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5159),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5168),
.Y(n_5238)
);

AND2x2_ASAP7_75t_L g5239 ( 
.A(n_5154),
.B(n_607),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_5133),
.Y(n_5240)
);

NOR2x1_ASAP7_75t_L g5241 ( 
.A(n_5173),
.B(n_608),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5187),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5217),
.Y(n_5243)
);

OR2x2_ASAP7_75t_L g5244 ( 
.A(n_5220),
.B(n_5216),
.Y(n_5244)
);

NAND2x1p5_ASAP7_75t_L g5245 ( 
.A(n_5219),
.B(n_5175),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_5191),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_5194),
.B(n_5187),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5222),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_5192),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_5235),
.B(n_5187),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_5224),
.Y(n_5251)
);

AND2x2_ASAP7_75t_L g5252 ( 
.A(n_5207),
.B(n_5146),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_5189),
.B(n_5179),
.Y(n_5253)
);

INVx1_ASAP7_75t_SL g5254 ( 
.A(n_5218),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5189),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_5197),
.B(n_5124),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5230),
.Y(n_5257)
);

HB1xp67_ASAP7_75t_L g5258 ( 
.A(n_5196),
.Y(n_5258)
);

OR2x2_ASAP7_75t_L g5259 ( 
.A(n_5199),
.B(n_5156),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_5231),
.B(n_5158),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_5198),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5226),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5221),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_5228),
.B(n_5162),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5201),
.Y(n_5265)
);

AND2x2_ASAP7_75t_L g5266 ( 
.A(n_5229),
.B(n_5141),
.Y(n_5266)
);

AOI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_5219),
.A2(n_5117),
.B(n_5171),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_5223),
.B(n_5165),
.Y(n_5268)
);

INVx3_ASAP7_75t_L g5269 ( 
.A(n_5229),
.Y(n_5269)
);

AND2x2_ASAP7_75t_L g5270 ( 
.A(n_5240),
.B(n_5169),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_5215),
.B(n_5160),
.Y(n_5271)
);

AND2x2_ASAP7_75t_L g5272 ( 
.A(n_5211),
.B(n_5129),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_5202),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_5213),
.B(n_5167),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_5234),
.Y(n_5275)
);

INVx3_ASAP7_75t_L g5276 ( 
.A(n_5234),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5242),
.B(n_5153),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_5212),
.B(n_5204),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5188),
.Y(n_5279)
);

OR2x2_ASAP7_75t_L g5280 ( 
.A(n_5208),
.B(n_609),
.Y(n_5280)
);

INVx2_ASAP7_75t_SL g5281 ( 
.A(n_5227),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_5239),
.B(n_5145),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_5190),
.Y(n_5283)
);

OR2x2_ASAP7_75t_L g5284 ( 
.A(n_5195),
.B(n_609),
.Y(n_5284)
);

AND2x2_ASAP7_75t_L g5285 ( 
.A(n_5236),
.B(n_5186),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5203),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_5225),
.B(n_610),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5209),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5205),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5206),
.B(n_5210),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5238),
.B(n_610),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_5214),
.B(n_611),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5232),
.Y(n_5293)
);

OR2x6_ASAP7_75t_L g5294 ( 
.A(n_5200),
.B(n_611),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5193),
.B(n_612),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5233),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_5237),
.B(n_613),
.Y(n_5297)
);

AND2x2_ASAP7_75t_L g5298 ( 
.A(n_5241),
.B(n_614),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_5217),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5217),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_5217),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_5194),
.B(n_615),
.Y(n_5302)
);

OR2x2_ASAP7_75t_L g5303 ( 
.A(n_5244),
.B(n_616),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5254),
.B(n_616),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5249),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5246),
.B(n_617),
.Y(n_5306)
);

NAND2x1p5_ASAP7_75t_L g5307 ( 
.A(n_5269),
.B(n_617),
.Y(n_5307)
);

OAI21xp33_ASAP7_75t_L g5308 ( 
.A1(n_5252),
.A2(n_951),
.B(n_618),
.Y(n_5308)
);

INVx1_ASAP7_75t_SL g5309 ( 
.A(n_5270),
.Y(n_5309)
);

OR2x2_ASAP7_75t_L g5310 ( 
.A(n_5257),
.B(n_618),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_5256),
.Y(n_5311)
);

AOI22xp33_ASAP7_75t_L g5312 ( 
.A1(n_5266),
.A2(n_623),
.B1(n_619),
.B2(n_621),
.Y(n_5312)
);

OR3x2_ASAP7_75t_L g5313 ( 
.A(n_5248),
.B(n_621),
.C(n_624),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_5277),
.B(n_624),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5263),
.B(n_625),
.Y(n_5315)
);

NOR2x1_ASAP7_75t_L g5316 ( 
.A(n_5269),
.B(n_5302),
.Y(n_5316)
);

NOR2xp33_ASAP7_75t_L g5317 ( 
.A(n_5245),
.B(n_5276),
.Y(n_5317)
);

HB1xp67_ASAP7_75t_L g5318 ( 
.A(n_5258),
.Y(n_5318)
);

INVx2_ASAP7_75t_SL g5319 ( 
.A(n_5272),
.Y(n_5319)
);

OR2x2_ASAP7_75t_L g5320 ( 
.A(n_5259),
.B(n_626),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_5261),
.Y(n_5321)
);

AND2x4_ASAP7_75t_L g5322 ( 
.A(n_5288),
.B(n_626),
.Y(n_5322)
);

NOR2xp33_ASAP7_75t_L g5323 ( 
.A(n_5276),
.B(n_627),
.Y(n_5323)
);

INVx2_ASAP7_75t_L g5324 ( 
.A(n_5275),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5243),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_5299),
.Y(n_5326)
);

OR2x2_ASAP7_75t_L g5327 ( 
.A(n_5264),
.B(n_627),
.Y(n_5327)
);

INVxp67_ASAP7_75t_L g5328 ( 
.A(n_5247),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_5300),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_5281),
.B(n_628),
.Y(n_5330)
);

AOI22xp33_ASAP7_75t_L g5331 ( 
.A1(n_5282),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5298),
.B(n_630),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_5285),
.B(n_631),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_5297),
.B(n_632),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5251),
.B(n_5262),
.Y(n_5335)
);

HB1xp67_ASAP7_75t_L g5336 ( 
.A(n_5301),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5297),
.B(n_632),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_5273),
.B(n_633),
.Y(n_5338)
);

AND2x2_ASAP7_75t_L g5339 ( 
.A(n_5250),
.B(n_633),
.Y(n_5339)
);

INVx1_ASAP7_75t_SL g5340 ( 
.A(n_5287),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_5289),
.B(n_5279),
.Y(n_5341)
);

AND2x2_ASAP7_75t_L g5342 ( 
.A(n_5294),
.B(n_634),
.Y(n_5342)
);

INVx2_ASAP7_75t_L g5343 ( 
.A(n_5283),
.Y(n_5343)
);

INVx2_ASAP7_75t_SL g5344 ( 
.A(n_5280),
.Y(n_5344)
);

NOR4xp25_ASAP7_75t_SL g5345 ( 
.A(n_5265),
.B(n_637),
.C(n_635),
.D(n_636),
.Y(n_5345)
);

INVx2_ASAP7_75t_L g5346 ( 
.A(n_5255),
.Y(n_5346)
);

NAND4xp25_ASAP7_75t_L g5347 ( 
.A(n_5268),
.B(n_639),
.C(n_636),
.D(n_637),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5295),
.Y(n_5348)
);

AND2x2_ASAP7_75t_L g5349 ( 
.A(n_5294),
.B(n_639),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5286),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_5267),
.B(n_640),
.Y(n_5351)
);

OAI221xp5_ASAP7_75t_L g5352 ( 
.A1(n_5253),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.C(n_644),
.Y(n_5352)
);

NAND2xp5_ASAP7_75t_L g5353 ( 
.A(n_5293),
.B(n_641),
.Y(n_5353)
);

OR2x2_ASAP7_75t_L g5354 ( 
.A(n_5284),
.B(n_643),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_5292),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5274),
.B(n_645),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_5309),
.B(n_5260),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5304),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5311),
.B(n_5271),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5319),
.B(n_5296),
.Y(n_5360)
);

OR2x2_ASAP7_75t_L g5361 ( 
.A(n_5315),
.B(n_5291),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5318),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5339),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_5333),
.B(n_5290),
.Y(n_5364)
);

INVxp67_ASAP7_75t_L g5365 ( 
.A(n_5317),
.Y(n_5365)
);

NAND5xp2_ASAP7_75t_SL g5366 ( 
.A(n_5331),
.B(n_5278),
.C(n_647),
.D(n_645),
.E(n_646),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_5324),
.B(n_646),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5321),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_5322),
.B(n_647),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_5322),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_SL g5371 ( 
.A(n_5351),
.B(n_648),
.Y(n_5371)
);

AND2x2_ASAP7_75t_L g5372 ( 
.A(n_5335),
.B(n_648),
.Y(n_5372)
);

INVx2_ASAP7_75t_L g5373 ( 
.A(n_5307),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5310),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_5340),
.B(n_650),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_5323),
.B(n_650),
.Y(n_5376)
);

AND2x2_ASAP7_75t_L g5377 ( 
.A(n_5355),
.B(n_651),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_5305),
.B(n_651),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5312),
.B(n_652),
.Y(n_5379)
);

NAND2xp67_ASAP7_75t_L g5380 ( 
.A(n_5343),
.B(n_653),
.Y(n_5380)
);

AND2x2_ASAP7_75t_L g5381 ( 
.A(n_5328),
.B(n_653),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_5334),
.Y(n_5382)
);

NAND2x1p5_ASAP7_75t_L g5383 ( 
.A(n_5342),
.B(n_951),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5337),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5349),
.Y(n_5385)
);

INVxp67_ASAP7_75t_SL g5386 ( 
.A(n_5306),
.Y(n_5386)
);

AND2x2_ASAP7_75t_L g5387 ( 
.A(n_5341),
.B(n_5344),
.Y(n_5387)
);

HB1xp67_ASAP7_75t_L g5388 ( 
.A(n_5330),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_5336),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_5308),
.B(n_654),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5316),
.B(n_949),
.Y(n_5391)
);

AND2x2_ASAP7_75t_L g5392 ( 
.A(n_5314),
.B(n_655),
.Y(n_5392)
);

INVx3_ASAP7_75t_L g5393 ( 
.A(n_5303),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_5345),
.B(n_655),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5354),
.Y(n_5395)
);

OR2x6_ASAP7_75t_L g5396 ( 
.A(n_5356),
.B(n_656),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_L g5397 ( 
.A(n_5348),
.B(n_656),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_5320),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_5332),
.Y(n_5399)
);

NOR2xp33_ASAP7_75t_L g5400 ( 
.A(n_5347),
.B(n_657),
.Y(n_5400)
);

CKINVDCx16_ASAP7_75t_R g5401 ( 
.A(n_5327),
.Y(n_5401)
);

AND2x4_ASAP7_75t_L g5402 ( 
.A(n_5346),
.B(n_657),
.Y(n_5402)
);

HB1xp67_ASAP7_75t_L g5403 ( 
.A(n_5325),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5338),
.Y(n_5404)
);

OR2x2_ASAP7_75t_L g5405 ( 
.A(n_5353),
.B(n_658),
.Y(n_5405)
);

AND2x2_ASAP7_75t_L g5406 ( 
.A(n_5326),
.B(n_948),
.Y(n_5406)
);

OR2x2_ASAP7_75t_L g5407 ( 
.A(n_5352),
.B(n_658),
.Y(n_5407)
);

INVx1_ASAP7_75t_SL g5408 ( 
.A(n_5367),
.Y(n_5408)
);

OR2x2_ASAP7_75t_L g5409 ( 
.A(n_5394),
.B(n_5407),
.Y(n_5409)
);

AND2x2_ASAP7_75t_SL g5410 ( 
.A(n_5357),
.B(n_5329),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5369),
.Y(n_5411)
);

AOI211x1_ASAP7_75t_L g5412 ( 
.A1(n_5359),
.A2(n_5350),
.B(n_5313),
.C(n_661),
.Y(n_5412)
);

AOI322xp5_ASAP7_75t_L g5413 ( 
.A1(n_5387),
.A2(n_5350),
.A3(n_667),
.B1(n_662),
.B2(n_666),
.C1(n_659),
.C2(n_660),
.Y(n_5413)
);

OAI21xp5_ASAP7_75t_L g5414 ( 
.A1(n_5365),
.A2(n_659),
.B(n_664),
.Y(n_5414)
);

OAI221xp5_ASAP7_75t_L g5415 ( 
.A1(n_5362),
.A2(n_668),
.B1(n_664),
.B2(n_666),
.C(n_669),
.Y(n_5415)
);

OAI22xp5_ASAP7_75t_L g5416 ( 
.A1(n_5373),
.A2(n_673),
.B1(n_670),
.B2(n_672),
.Y(n_5416)
);

AOI22xp5_ASAP7_75t_L g5417 ( 
.A1(n_5400),
.A2(n_676),
.B1(n_672),
.B2(n_674),
.Y(n_5417)
);

INVx4_ASAP7_75t_L g5418 ( 
.A(n_5402),
.Y(n_5418)
);

AND2x2_ASAP7_75t_L g5419 ( 
.A(n_5372),
.B(n_5381),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_5370),
.Y(n_5420)
);

AND2x2_ASAP7_75t_L g5421 ( 
.A(n_5377),
.B(n_674),
.Y(n_5421)
);

AND2x4_ASAP7_75t_L g5422 ( 
.A(n_5368),
.B(n_676),
.Y(n_5422)
);

INVx1_ASAP7_75t_SL g5423 ( 
.A(n_5402),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5391),
.Y(n_5424)
);

OAI211xp5_ASAP7_75t_SL g5425 ( 
.A1(n_5360),
.A2(n_679),
.B(n_677),
.C(n_678),
.Y(n_5425)
);

AOI211x1_ASAP7_75t_L g5426 ( 
.A1(n_5364),
.A2(n_679),
.B(n_677),
.C(n_678),
.Y(n_5426)
);

NOR2xp33_ASAP7_75t_L g5427 ( 
.A(n_5401),
.B(n_680),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_5378),
.Y(n_5428)
);

NAND2x1_ASAP7_75t_L g5429 ( 
.A(n_5389),
.B(n_681),
.Y(n_5429)
);

INVx1_ASAP7_75t_SL g5430 ( 
.A(n_5405),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5392),
.B(n_681),
.Y(n_5431)
);

NAND4xp75_ASAP7_75t_SL g5432 ( 
.A(n_5406),
.B(n_685),
.C(n_682),
.D(n_683),
.Y(n_5432)
);

NAND2x1_ASAP7_75t_L g5433 ( 
.A(n_5393),
.B(n_682),
.Y(n_5433)
);

INVx2_ASAP7_75t_L g5434 ( 
.A(n_5383),
.Y(n_5434)
);

A2O1A1Ixp33_ASAP7_75t_L g5435 ( 
.A1(n_5363),
.A2(n_689),
.B(n_686),
.C(n_687),
.Y(n_5435)
);

NOR3xp33_ASAP7_75t_L g5436 ( 
.A(n_5397),
.B(n_686),
.C(n_689),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5375),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_5380),
.B(n_5399),
.Y(n_5438)
);

AOI21xp5_ASAP7_75t_L g5439 ( 
.A1(n_5371),
.A2(n_691),
.B(n_692),
.Y(n_5439)
);

AOI322xp5_ASAP7_75t_L g5440 ( 
.A1(n_5386),
.A2(n_697),
.A3(n_696),
.B1(n_694),
.B2(n_691),
.C1(n_693),
.C2(n_695),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_5398),
.Y(n_5441)
);

NOR2xp33_ASAP7_75t_L g5442 ( 
.A(n_5385),
.B(n_693),
.Y(n_5442)
);

OAI22xp33_ASAP7_75t_L g5443 ( 
.A1(n_5396),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_5443)
);

AOI22xp5_ASAP7_75t_L g5444 ( 
.A1(n_5374),
.A2(n_699),
.B1(n_697),
.B2(n_698),
.Y(n_5444)
);

OAI22xp5_ASAP7_75t_L g5445 ( 
.A1(n_5396),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.Y(n_5445)
);

HB1xp67_ASAP7_75t_L g5446 ( 
.A(n_5403),
.Y(n_5446)
);

INVxp67_ASAP7_75t_L g5447 ( 
.A(n_5376),
.Y(n_5447)
);

OAI21xp33_ASAP7_75t_L g5448 ( 
.A1(n_5395),
.A2(n_701),
.B(n_702),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_5382),
.B(n_701),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5390),
.Y(n_5450)
);

OA21x2_ASAP7_75t_SL g5451 ( 
.A1(n_5379),
.A2(n_703),
.B(n_704),
.Y(n_5451)
);

AOI22xp5_ASAP7_75t_L g5452 ( 
.A1(n_5358),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_5452)
);

NAND2x1p5_ASAP7_75t_L g5453 ( 
.A(n_5420),
.B(n_5384),
.Y(n_5453)
);

AND2x2_ASAP7_75t_L g5454 ( 
.A(n_5421),
.B(n_5388),
.Y(n_5454)
);

NAND2xp5_ASAP7_75t_SL g5455 ( 
.A(n_5422),
.B(n_5404),
.Y(n_5455)
);

NAND2xp5_ASAP7_75t_L g5456 ( 
.A(n_5413),
.B(n_5361),
.Y(n_5456)
);

OR2x2_ASAP7_75t_L g5457 ( 
.A(n_5433),
.B(n_5366),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5418),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5446),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5431),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5429),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5427),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_5410),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5422),
.Y(n_5464)
);

INVx1_ASAP7_75t_SL g5465 ( 
.A(n_5423),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5409),
.Y(n_5466)
);

INVxp67_ASAP7_75t_L g5467 ( 
.A(n_5442),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5441),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5419),
.B(n_707),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_5408),
.B(n_948),
.Y(n_5470)
);

NAND2x1_ASAP7_75t_SL g5471 ( 
.A(n_5418),
.B(n_708),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_5440),
.B(n_708),
.Y(n_5472)
);

OR2x2_ASAP7_75t_L g5473 ( 
.A(n_5445),
.B(n_5435),
.Y(n_5473)
);

NOR2xp33_ASAP7_75t_L g5474 ( 
.A(n_5424),
.B(n_5448),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5416),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5412),
.B(n_709),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_5426),
.B(n_709),
.Y(n_5477)
);

INVxp67_ASAP7_75t_L g5478 ( 
.A(n_5415),
.Y(n_5478)
);

INVxp67_ASAP7_75t_L g5479 ( 
.A(n_5449),
.Y(n_5479)
);

NOR2xp33_ASAP7_75t_L g5480 ( 
.A(n_5434),
.B(n_710),
.Y(n_5480)
);

INVx1_ASAP7_75t_SL g5481 ( 
.A(n_5430),
.Y(n_5481)
);

AND2x2_ASAP7_75t_L g5482 ( 
.A(n_5437),
.B(n_5411),
.Y(n_5482)
);

INVx1_ASAP7_75t_SL g5483 ( 
.A(n_5432),
.Y(n_5483)
);

NOR2xp33_ASAP7_75t_L g5484 ( 
.A(n_5438),
.B(n_710),
.Y(n_5484)
);

AND2x2_ASAP7_75t_L g5485 ( 
.A(n_5428),
.B(n_947),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5444),
.Y(n_5486)
);

AND2x2_ASAP7_75t_L g5487 ( 
.A(n_5447),
.B(n_712),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5450),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5452),
.Y(n_5489)
);

NAND4xp25_ASAP7_75t_L g5490 ( 
.A(n_5451),
.B(n_715),
.C(n_713),
.D(n_714),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5443),
.Y(n_5491)
);

OAI21xp5_ASAP7_75t_L g5492 ( 
.A1(n_5439),
.A2(n_715),
.B(n_717),
.Y(n_5492)
);

AND3x2_ASAP7_75t_L g5493 ( 
.A(n_5458),
.B(n_5436),
.C(n_5414),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5468),
.Y(n_5494)
);

NOR2xp33_ASAP7_75t_L g5495 ( 
.A(n_5490),
.B(n_5425),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5465),
.B(n_5417),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_5469),
.B(n_717),
.Y(n_5497)
);

BUFx2_ASAP7_75t_L g5498 ( 
.A(n_5471),
.Y(n_5498)
);

NOR4xp25_ASAP7_75t_SL g5499 ( 
.A(n_5463),
.B(n_720),
.C(n_718),
.D(n_719),
.Y(n_5499)
);

INVx2_ASAP7_75t_L g5500 ( 
.A(n_5453),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5481),
.B(n_719),
.Y(n_5501)
);

OAI21xp5_ASAP7_75t_SL g5502 ( 
.A1(n_5483),
.A2(n_5490),
.B(n_5478),
.Y(n_5502)
);

NAND2xp5_ASAP7_75t_L g5503 ( 
.A(n_5459),
.B(n_720),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_5470),
.Y(n_5504)
);

INVxp67_ASAP7_75t_L g5505 ( 
.A(n_5480),
.Y(n_5505)
);

INVx2_ASAP7_75t_L g5506 ( 
.A(n_5464),
.Y(n_5506)
);

INVx1_ASAP7_75t_SL g5507 ( 
.A(n_5457),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5487),
.Y(n_5508)
);

NOR2x1_ASAP7_75t_L g5509 ( 
.A(n_5476),
.B(n_721),
.Y(n_5509)
);

OAI22xp5_ASAP7_75t_L g5510 ( 
.A1(n_5491),
.A2(n_723),
.B1(n_721),
.B2(n_722),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5485),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_L g5512 ( 
.A(n_5461),
.B(n_722),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5488),
.Y(n_5513)
);

OAI32xp33_ASAP7_75t_L g5514 ( 
.A1(n_5473),
.A2(n_725),
.A3(n_723),
.B1(n_724),
.B2(n_726),
.Y(n_5514)
);

NOR3xp33_ASAP7_75t_SL g5515 ( 
.A(n_5484),
.B(n_724),
.C(n_725),
.Y(n_5515)
);

NOR2xp33_ASAP7_75t_L g5516 ( 
.A(n_5472),
.B(n_726),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_5454),
.B(n_727),
.Y(n_5517)
);

AND2x2_ASAP7_75t_L g5518 ( 
.A(n_5466),
.B(n_5475),
.Y(n_5518)
);

NOR2xp33_ASAP7_75t_L g5519 ( 
.A(n_5477),
.B(n_5486),
.Y(n_5519)
);

BUFx4f_ASAP7_75t_SL g5520 ( 
.A(n_5455),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5489),
.Y(n_5521)
);

INVx1_ASAP7_75t_SL g5522 ( 
.A(n_5482),
.Y(n_5522)
);

CKINVDCx14_ASAP7_75t_R g5523 ( 
.A(n_5462),
.Y(n_5523)
);

AOI21xp5_ASAP7_75t_L g5524 ( 
.A1(n_5502),
.A2(n_5456),
.B(n_5474),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_SL g5525 ( 
.A(n_5500),
.B(n_5467),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5494),
.Y(n_5526)
);

NAND4xp25_ASAP7_75t_L g5527 ( 
.A(n_5507),
.B(n_5492),
.C(n_5460),
.D(n_5479),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5513),
.Y(n_5528)
);

NOR2xp33_ASAP7_75t_L g5529 ( 
.A(n_5522),
.B(n_5510),
.Y(n_5529)
);

INVxp67_ASAP7_75t_L g5530 ( 
.A(n_5517),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5506),
.B(n_728),
.Y(n_5531)
);

NOR3x1_ASAP7_75t_L g5532 ( 
.A(n_5497),
.B(n_728),
.C(n_729),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_5520),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5512),
.Y(n_5534)
);

NOR3xp33_ASAP7_75t_L g5535 ( 
.A(n_5514),
.B(n_5521),
.C(n_5501),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5518),
.Y(n_5536)
);

NOR2xp33_ASAP7_75t_L g5537 ( 
.A(n_5495),
.B(n_730),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_L g5538 ( 
.A(n_5499),
.B(n_731),
.Y(n_5538)
);

NOR3xp33_ASAP7_75t_L g5539 ( 
.A(n_5523),
.B(n_731),
.C(n_732),
.Y(n_5539)
);

INVxp67_ASAP7_75t_L g5540 ( 
.A(n_5503),
.Y(n_5540)
);

AND2x4_ASAP7_75t_L g5541 ( 
.A(n_5498),
.B(n_732),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_5493),
.B(n_733),
.Y(n_5542)
);

NAND2xp5_ASAP7_75t_L g5543 ( 
.A(n_5516),
.B(n_734),
.Y(n_5543)
);

NAND5xp2_ASAP7_75t_L g5544 ( 
.A(n_5519),
.B(n_5515),
.C(n_5496),
.D(n_5504),
.E(n_5508),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_5505),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_5533),
.B(n_5528),
.Y(n_5546)
);

NOR2xp33_ASAP7_75t_L g5547 ( 
.A(n_5538),
.B(n_5511),
.Y(n_5547)
);

NOR2xp33_ASAP7_75t_L g5548 ( 
.A(n_5536),
.B(n_5509),
.Y(n_5548)
);

AOI21xp5_ASAP7_75t_L g5549 ( 
.A1(n_5524),
.A2(n_734),
.B(n_735),
.Y(n_5549)
);

NAND4xp25_ASAP7_75t_L g5550 ( 
.A(n_5544),
.B(n_737),
.C(n_735),
.D(n_736),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5541),
.B(n_737),
.Y(n_5551)
);

AND2x2_ASAP7_75t_L g5552 ( 
.A(n_5541),
.B(n_738),
.Y(n_5552)
);

AOI222xp33_ASAP7_75t_L g5553 ( 
.A1(n_5526),
.A2(n_741),
.B1(n_743),
.B2(n_738),
.C1(n_740),
.C2(n_742),
.Y(n_5553)
);

NAND2xp5_ASAP7_75t_L g5554 ( 
.A(n_5539),
.B(n_742),
.Y(n_5554)
);

NOR2x1_ASAP7_75t_L g5555 ( 
.A(n_5527),
.B(n_743),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5542),
.Y(n_5556)
);

NAND3xp33_ASAP7_75t_L g5557 ( 
.A(n_5535),
.B(n_744),
.C(n_746),
.Y(n_5557)
);

NAND4xp25_ASAP7_75t_L g5558 ( 
.A(n_5529),
.B(n_5537),
.C(n_5532),
.D(n_5525),
.Y(n_5558)
);

NOR3xp33_ASAP7_75t_L g5559 ( 
.A(n_5531),
.B(n_746),
.C(n_747),
.Y(n_5559)
);

NAND2xp5_ASAP7_75t_SL g5560 ( 
.A(n_5543),
.B(n_747),
.Y(n_5560)
);

OAI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_5530),
.A2(n_748),
.B(n_749),
.Y(n_5561)
);

AOI21xp5_ASAP7_75t_L g5562 ( 
.A1(n_5545),
.A2(n_748),
.B(n_749),
.Y(n_5562)
);

AND3x2_ASAP7_75t_L g5563 ( 
.A(n_5540),
.B(n_750),
.C(n_751),
.Y(n_5563)
);

NAND2xp5_ASAP7_75t_L g5564 ( 
.A(n_5534),
.B(n_750),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_5528),
.B(n_946),
.Y(n_5565)
);

OAI221xp5_ASAP7_75t_L g5566 ( 
.A1(n_5528),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.C(n_755),
.Y(n_5566)
);

NAND3xp33_ASAP7_75t_L g5567 ( 
.A(n_5539),
.B(n_752),
.C(n_753),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5546),
.Y(n_5568)
);

NAND2xp5_ASAP7_75t_L g5569 ( 
.A(n_5563),
.B(n_754),
.Y(n_5569)
);

AOI221xp5_ASAP7_75t_L g5570 ( 
.A1(n_5566),
.A2(n_759),
.B1(n_756),
.B2(n_757),
.C(n_760),
.Y(n_5570)
);

HB1xp67_ASAP7_75t_L g5571 ( 
.A(n_5552),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_SL g5572 ( 
.A(n_5549),
.B(n_757),
.Y(n_5572)
);

NOR2xp67_ASAP7_75t_L g5573 ( 
.A(n_5550),
.B(n_759),
.Y(n_5573)
);

AND2x4_ASAP7_75t_L g5574 ( 
.A(n_5557),
.B(n_760),
.Y(n_5574)
);

INVxp67_ASAP7_75t_L g5575 ( 
.A(n_5551),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5565),
.Y(n_5576)
);

AOI22xp33_ASAP7_75t_L g5577 ( 
.A1(n_5559),
.A2(n_764),
.B1(n_761),
.B2(n_762),
.Y(n_5577)
);

NAND2xp5_ASAP7_75t_L g5578 ( 
.A(n_5553),
.B(n_761),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5564),
.Y(n_5579)
);

AOI31xp33_ASAP7_75t_L g5580 ( 
.A1(n_5554),
.A2(n_946),
.A3(n_766),
.B(n_762),
.Y(n_5580)
);

OAI22xp5_ASAP7_75t_L g5581 ( 
.A1(n_5568),
.A2(n_5556),
.B1(n_5547),
.B2(n_5555),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5569),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5578),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_5571),
.Y(n_5584)
);

AOI211xp5_ASAP7_75t_SL g5585 ( 
.A1(n_5580),
.A2(n_5548),
.B(n_5562),
.C(n_5558),
.Y(n_5585)
);

NAND3xp33_ASAP7_75t_L g5586 ( 
.A(n_5570),
.B(n_5561),
.C(n_5567),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5573),
.Y(n_5587)
);

BUFx24_ASAP7_75t_SL g5588 ( 
.A(n_5577),
.Y(n_5588)
);

NOR2x1p5_ASAP7_75t_L g5589 ( 
.A(n_5576),
.B(n_5560),
.Y(n_5589)
);

NOR2x1_ASAP7_75t_L g5590 ( 
.A(n_5579),
.B(n_765),
.Y(n_5590)
);

NOR2x1_ASAP7_75t_L g5591 ( 
.A(n_5572),
.B(n_765),
.Y(n_5591)
);

NOR2x1_ASAP7_75t_L g5592 ( 
.A(n_5574),
.B(n_5575),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5574),
.Y(n_5593)
);

AND2x4_ASAP7_75t_L g5594 ( 
.A(n_5568),
.B(n_766),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5568),
.Y(n_5595)
);

INVx3_ASAP7_75t_L g5596 ( 
.A(n_5594),
.Y(n_5596)
);

NOR3xp33_ASAP7_75t_L g5597 ( 
.A(n_5581),
.B(n_943),
.C(n_767),
.Y(n_5597)
);

AND3x4_ASAP7_75t_L g5598 ( 
.A(n_5588),
.B(n_5592),
.C(n_5591),
.Y(n_5598)
);

NOR2x1_ASAP7_75t_L g5599 ( 
.A(n_5595),
.B(n_768),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_5594),
.B(n_769),
.Y(n_5600)
);

OAI221xp5_ASAP7_75t_SL g5601 ( 
.A1(n_5584),
.A2(n_772),
.B1(n_770),
.B2(n_771),
.C(n_774),
.Y(n_5601)
);

NOR2x1_ASAP7_75t_L g5602 ( 
.A(n_5586),
.B(n_770),
.Y(n_5602)
);

AND2x4_ASAP7_75t_L g5603 ( 
.A(n_5593),
.B(n_771),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5600),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_5603),
.Y(n_5605)
);

INVx2_ASAP7_75t_L g5606 ( 
.A(n_5596),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5599),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_SL g5608 ( 
.A(n_5597),
.B(n_5583),
.Y(n_5608)
);

XNOR2xp5_ASAP7_75t_L g5609 ( 
.A(n_5598),
.B(n_5589),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_5602),
.B(n_5590),
.Y(n_5610)
);

NOR2xp33_ASAP7_75t_L g5611 ( 
.A(n_5601),
.B(n_5587),
.Y(n_5611)
);

OAI22x1_ASAP7_75t_L g5612 ( 
.A1(n_5598),
.A2(n_5582),
.B1(n_5585),
.B2(n_775),
.Y(n_5612)
);

OR2x2_ASAP7_75t_L g5613 ( 
.A(n_5600),
.B(n_772),
.Y(n_5613)
);

HB1xp67_ASAP7_75t_L g5614 ( 
.A(n_5599),
.Y(n_5614)
);

INVx4_ASAP7_75t_L g5615 ( 
.A(n_5606),
.Y(n_5615)
);

INVx1_ASAP7_75t_SL g5616 ( 
.A(n_5613),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5609),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5612),
.Y(n_5618)
);

AOI22xp5_ASAP7_75t_L g5619 ( 
.A1(n_5611),
.A2(n_778),
.B1(n_774),
.B2(n_776),
.Y(n_5619)
);

AND2x2_ASAP7_75t_L g5620 ( 
.A(n_5605),
.B(n_776),
.Y(n_5620)
);

AOI221xp5_ASAP7_75t_L g5621 ( 
.A1(n_5608),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.C(n_782),
.Y(n_5621)
);

NOR2xp33_ASAP7_75t_L g5622 ( 
.A(n_5615),
.B(n_5604),
.Y(n_5622)
);

A2O1A1Ixp33_ASAP7_75t_L g5623 ( 
.A1(n_5618),
.A2(n_5607),
.B(n_5610),
.C(n_5614),
.Y(n_5623)
);

NAND4xp75_ASAP7_75t_L g5624 ( 
.A(n_5617),
.B(n_782),
.C(n_779),
.D(n_780),
.Y(n_5624)
);

AOI22xp5_ASAP7_75t_L g5625 ( 
.A1(n_5620),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_5625)
);

HB1xp67_ASAP7_75t_L g5626 ( 
.A(n_5616),
.Y(n_5626)
);

AOI211xp5_ASAP7_75t_SL g5627 ( 
.A1(n_5621),
.A2(n_786),
.B(n_783),
.C(n_785),
.Y(n_5627)
);

AOI21xp5_ASAP7_75t_L g5628 ( 
.A1(n_5619),
.A2(n_941),
.B(n_786),
.Y(n_5628)
);

AOI221xp5_ASAP7_75t_L g5629 ( 
.A1(n_5622),
.A2(n_5623),
.B1(n_5626),
.B2(n_5628),
.C(n_5625),
.Y(n_5629)
);

NAND4xp25_ASAP7_75t_L g5630 ( 
.A(n_5627),
.B(n_5624),
.C(n_790),
.D(n_788),
.Y(n_5630)
);

OR2x6_ASAP7_75t_L g5631 ( 
.A(n_5626),
.B(n_789),
.Y(n_5631)
);

NOR2xp33_ASAP7_75t_L g5632 ( 
.A(n_5622),
.B(n_789),
.Y(n_5632)
);

AOI21xp5_ASAP7_75t_L g5633 ( 
.A1(n_5629),
.A2(n_791),
.B(n_792),
.Y(n_5633)
);

AOI21xp5_ASAP7_75t_L g5634 ( 
.A1(n_5631),
.A2(n_792),
.B(n_793),
.Y(n_5634)
);

OR3x2_ASAP7_75t_L g5635 ( 
.A(n_5634),
.B(n_5630),
.C(n_5632),
.Y(n_5635)
);

OAI31xp33_ASAP7_75t_SL g5636 ( 
.A1(n_5635),
.A2(n_5633),
.A3(n_796),
.B(n_794),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5636),
.B(n_795),
.Y(n_5637)
);

NAND3xp33_ASAP7_75t_L g5638 ( 
.A(n_5637),
.B(n_795),
.C(n_796),
.Y(n_5638)
);

INVxp67_ASAP7_75t_L g5639 ( 
.A(n_5638),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5639),
.B(n_797),
.Y(n_5640)
);

AOI21xp33_ASAP7_75t_L g5641 ( 
.A1(n_5640),
.A2(n_797),
.B(n_798),
.Y(n_5641)
);

AOI211xp5_ASAP7_75t_L g5642 ( 
.A1(n_5641),
.A2(n_802),
.B(n_799),
.C(n_801),
.Y(n_5642)
);


endmodule