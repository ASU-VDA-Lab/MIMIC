module fake_jpeg_318_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.Y(n_58)
);

NAND2x1_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_41),
.B1(n_28),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_60),
.B1(n_38),
.B2(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_30),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_53),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_53),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_36),
.C(n_31),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_61),
.B1(n_60),
.B2(n_63),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_14),
.B1(n_26),
.B2(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_85),
.B(n_1),
.Y(n_86)
);

OR2x4_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_92),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_71),
.B(n_4),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_91),
.B(n_8),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_78),
.B1(n_79),
.B2(n_83),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_93),
.B1(n_95),
.B2(n_8),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_71),
.B(n_4),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_6),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_7),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_100),
.B1(n_88),
.B2(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_91),
.C(n_98),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_98),
.B(n_102),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_96),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_9),
.B(n_10),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_9),
.A3(n_11),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_22),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_24),
.Y(n_110)
);


endmodule