module fake_jpeg_7099_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_18),
.Y(n_55)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_27),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_45),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_35),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_29),
.C(n_20),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_65),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_26),
.B1(n_35),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_35),
.B1(n_26),
.B2(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_80),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_86),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_87),
.B1(n_33),
.B2(n_27),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_34),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_45),
.B1(n_38),
.B2(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_59),
.B1(n_66),
.B2(n_65),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_37),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_67),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_41),
.B1(n_45),
.B2(n_43),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_44),
.B(n_30),
.C(n_25),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_58),
.B(n_68),
.C(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_96),
.C(n_103),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_30),
.B(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_107),
.B1(n_115),
.B2(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_53),
.B1(n_66),
.B2(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_104),
.B1(n_110),
.B2(n_117),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_19),
.B(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_17),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_44),
.B1(n_32),
.B2(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_111),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_70),
.B1(n_77),
.B2(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_30),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_84),
.B1(n_83),
.B2(n_92),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_68),
.B(n_50),
.C(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_133),
.Y(n_145)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_110),
.B1(n_115),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_138),
.B1(n_83),
.B2(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_137),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_140),
.B(n_79),
.Y(n_157)
);

INVxp33_ASAP7_75t_SL g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_91),
.B1(n_92),
.B2(n_75),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_24),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_109),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_104),
.B1(n_113),
.B2(n_99),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_148),
.B1(n_164),
.B2(n_157),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_113),
.C(n_75),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_149),
.C(n_155),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_104),
.B1(n_113),
.B2(n_108),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_109),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_140),
.B1(n_122),
.B2(n_123),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_127),
.A3(n_124),
.B1(n_125),
.B2(n_120),
.C1(n_132),
.C2(n_134),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_137),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_161),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_165),
.B(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_131),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_89),
.B1(n_68),
.B2(n_71),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_73),
.B(n_32),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_151),
.B1(n_143),
.B2(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_146),
.B(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_184),
.B1(n_166),
.B2(n_143),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_181),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_160),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_142),
.C(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_182),
.C(n_172),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_24),
.C(n_15),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_24),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_71),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_72),
.Y(n_186)
);

AOI321xp33_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_148),
.A3(n_164),
.B1(n_25),
.B2(n_31),
.C(n_4),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_177),
.CI(n_182),
.CON(n_209),
.SN(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_196),
.B1(n_184),
.B2(n_179),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_168),
.B(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_145),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_199),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_145),
.B1(n_156),
.B2(n_146),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_144),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_178),
.B(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_31),
.B1(n_25),
.B2(n_2),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_203),
.B1(n_173),
.B2(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_209),
.C(n_216),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_167),
.B(n_171),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_214),
.B1(n_215),
.B2(n_3),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_189),
.B1(n_196),
.B2(n_201),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_215),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_3),
.B(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_222),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_195),
.C(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_193),
.C(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_192),
.C(n_187),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_190),
.Y(n_223)
);

OAI221xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_226),
.B1(n_214),
.B2(n_207),
.C(n_9),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_14),
.B(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_209),
.B1(n_8),
.B2(n_10),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_6),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_225),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_221),
.B1(n_220),
.B2(n_11),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_10),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_8),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_12),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_229),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_240),
.Y(n_245)
);

OAI21x1_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_240),
.B(n_12),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_246),
.B(n_12),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.Y(n_250)
);


endmodule