module fake_jpeg_21752_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_33),
.B(n_12),
.Y(n_48)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_29),
.B1(n_24),
.B2(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_20),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_68),
.B1(n_38),
.B2(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_61),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_32),
.B1(n_26),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_22),
.B1(n_21),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_22),
.B1(n_25),
.B2(n_19),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_38),
.B1(n_39),
.B2(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_79),
.B1(n_61),
.B2(n_53),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_35),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_27),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_41),
.B1(n_43),
.B2(n_34),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_88),
.B1(n_35),
.B2(n_14),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_21),
.B1(n_31),
.B2(n_12),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_49),
.B1(n_16),
.B2(n_17),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_50),
.B1(n_67),
.B2(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_94),
.B1(n_101),
.B2(n_107),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_73),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_63),
.C(n_51),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_18),
.C(n_15),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_55),
.B(n_12),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_103),
.B(n_83),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_59),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_56),
.B1(n_54),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_78),
.B1(n_84),
.B2(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_83),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_85),
.B(n_83),
.C(n_88),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_130),
.B1(n_77),
.B2(n_100),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_82),
.B(n_88),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_131),
.C(n_18),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_132),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_88),
.B(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_124),
.B(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_125),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_81),
.B(n_85),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_83),
.A3(n_86),
.B1(n_80),
.B2(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_23),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_13),
.B(n_19),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_78),
.B1(n_77),
.B2(n_16),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_107),
.B1(n_106),
.B2(n_95),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_140),
.B1(n_145),
.B2(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_107),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_156),
.B(n_110),
.Y(n_168)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_143),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_92),
.B1(n_108),
.B2(n_109),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_154),
.B1(n_150),
.B2(n_139),
.Y(n_160)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_97),
.B1(n_16),
.B2(n_17),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_23),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

OAI22x1_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_100),
.B1(n_18),
.B2(n_14),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_127),
.B(n_111),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_16),
.B1(n_17),
.B2(n_13),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_131),
.C(n_130),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_161),
.C(n_164),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_173),
.B1(n_183),
.B2(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_117),
.C(n_112),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_110),
.C(n_116),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_177),
.B(n_1),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_116),
.B1(n_118),
.B2(n_2),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_175),
.B1(n_144),
.B2(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_140),
.C(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_137),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_118),
.B1(n_19),
.B2(n_13),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_8),
.B(n_11),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_181),
.C(n_7),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_14),
.B(n_3),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_23),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_155),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_15),
.B1(n_14),
.B2(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_205),
.B1(n_175),
.B2(n_170),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_196),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_136),
.B1(n_143),
.B2(n_137),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_202),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_7),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_200),
.B1(n_177),
.B2(n_174),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_1),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_159),
.C(n_172),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_183),
.C(n_197),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_168),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_192),
.B1(n_202),
.B2(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_200),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_229),
.B1(n_3),
.B2(n_4),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_205),
.B(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_179),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_213),
.B1(n_219),
.B2(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_221),
.B1(n_204),
.B2(n_167),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_189),
.B1(n_172),
.B2(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_222),
.B1(n_227),
.B2(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_203),
.B1(n_167),
.B2(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_216),
.C(n_214),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_238),
.C(n_233),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_220),
.B1(n_208),
.B2(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_249),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_230),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_4),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_251),
.C(n_247),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_230),
.C(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_258),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_6),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_4),
.C(n_5),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_251),
.B1(n_6),
.B2(n_7),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_5),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_6),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_277),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_8),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_275),
.B(n_273),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_276),
.B(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_280),
.C(n_10),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_9),
.B(n_10),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_9),
.B(n_11),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_9),
.CI(n_11),
.CON(n_287),
.SN(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_11),
.Y(n_288)
);


endmodule