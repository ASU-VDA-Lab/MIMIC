module fake_netlist_1_2708_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_2), .B(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_6), .B(n_0), .Y(n_10) );
NOR3x1_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .C(n_7), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_9), .B(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
OA21x2_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_9), .B(n_11), .Y(n_14) );
endmodule