module fake_jpeg_17436_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_1),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_41),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_47),
.B1(n_57),
.B2(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_79),
.B1(n_80),
.B2(n_3),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_59),
.B1(n_56),
.B2(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_53),
.B1(n_50),
.B2(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_2),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_52),
.C(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_55),
.B1(n_49),
.B2(n_45),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_49),
.B1(n_45),
.B2(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_53),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_79),
.B(n_4),
.C(n_5),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_29),
.B1(n_40),
.B2(n_12),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_82),
.C(n_74),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_92),
.C(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_82),
.B1(n_87),
.B2(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_83),
.B1(n_78),
.B2(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_6),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_94),
.B(n_86),
.Y(n_103)
);

OAI321xp33_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_103),
.A3(n_97),
.B1(n_78),
.B2(n_7),
.C(n_19),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.C(n_7),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_13),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_18),
.C(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_21),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_28),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_30),
.B(n_33),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_34),
.B(n_36),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_38),
.Y(n_114)
);


endmodule