module real_aes_7543_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g446 ( .A(n_0), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_1), .A2(n_124), .B(n_128), .C(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_2), .A2(n_158), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g513 ( .A(n_3), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_4), .B(n_225), .Y(n_244) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_158), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g124 ( .A(n_6), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g199 ( .A(n_7), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_8), .B(n_41), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_9), .A2(n_157), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_10), .B(n_136), .Y(n_211) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_12), .B(n_239), .Y(n_537) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g549 ( .A(n_14), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_15), .A2(n_134), .B(n_221), .C(n_223), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_16), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_17), .B(n_501), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_18), .B(n_158), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_19), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_20), .A2(n_239), .B(n_254), .C(n_256), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_21), .B(n_225), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_22), .B(n_136), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_23), .A2(n_166), .B(n_223), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_24), .B(n_136), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_25), .Y(n_175) );
INVx1_ASAP7_75t_L g132 ( .A(n_26), .Y(n_132) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_27), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_28), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_29), .B(n_136), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_30), .A2(n_31), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_30), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_31), .Y(n_747) );
INVx1_ASAP7_75t_L g164 ( .A(n_32), .Y(n_164) );
INVx1_ASAP7_75t_L g492 ( .A(n_33), .Y(n_492) );
INVx2_ASAP7_75t_L g122 ( .A(n_34), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_35), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_36), .A2(n_239), .B(n_240), .C(n_242), .Y(n_238) );
INVxp67_ASAP7_75t_L g165 ( .A(n_37), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_38), .A2(n_128), .B(n_131), .C(n_139), .Y(n_127) );
CKINVDCx14_ASAP7_75t_R g237 ( .A(n_39), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_40), .A2(n_124), .B(n_128), .C(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g491 ( .A(n_42), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_43), .A2(n_183), .B(n_197), .C(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_44), .B(n_136), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_45), .A2(n_744), .B1(n_750), .B2(n_751), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_45), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_46), .A2(n_745), .B1(n_746), .B2(n_749), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_46), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_47), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_48), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_49), .B(n_440), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_50), .A2(n_444), .B1(n_463), .B2(n_752), .Y(n_462) );
INVx1_ASAP7_75t_L g252 ( .A(n_51), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_52), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_53), .B(n_158), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_54), .A2(n_128), .B1(n_256), .B2(n_490), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_55), .A2(n_104), .B1(n_449), .B2(n_458), .C1(n_461), .C2(n_753), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_55), .A2(n_70), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_55), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_56), .Y(n_510) );
CKINVDCx14_ASAP7_75t_R g195 ( .A(n_57), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_58), .A2(n_197), .B(n_242), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_59), .Y(n_565) );
INVx1_ASAP7_75t_L g480 ( .A(n_60), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_61), .A2(n_90), .B1(n_438), .B2(n_439), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_61), .Y(n_439) );
INVx1_ASAP7_75t_L g125 ( .A(n_62), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_63), .Y(n_143) );
INVx1_ASAP7_75t_SL g241 ( .A(n_64), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_65), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_66), .B(n_225), .Y(n_258) );
INVx1_ASAP7_75t_L g178 ( .A(n_67), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_68), .A2(n_242), .B(n_501), .C(n_502), .Y(n_500) );
INVxp67_ASAP7_75t_L g503 ( .A(n_69), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_L g457 ( .A(n_71), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_72), .A2(n_158), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_73), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_74), .A2(n_158), .B(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_75), .Y(n_495) );
INVx1_ASAP7_75t_L g559 ( .A(n_76), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_77), .A2(n_157), .B(n_159), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g219 ( .A(n_79), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_80), .A2(n_124), .B(n_128), .C(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_81), .A2(n_158), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g222 ( .A(n_82), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_83), .B(n_133), .Y(n_526) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx1_ASAP7_75t_L g210 ( .A(n_85), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_86), .B(n_501), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_87), .A2(n_124), .B(n_128), .C(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g443 ( .A(n_88), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g466 ( .A(n_88), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_89), .A2(n_128), .B(n_177), .C(n_185), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_90), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_91), .B(n_140), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_92), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_93), .A2(n_124), .B(n_128), .C(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_94), .Y(n_541) );
INVx1_ASAP7_75t_L g499 ( .A(n_95), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_96), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_97), .B(n_133), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_98), .B(n_148), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_99), .B(n_148), .Y(n_550) );
INVx2_ASAP7_75t_L g255 ( .A(n_100), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_101), .B(n_457), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_102), .A2(n_158), .B(n_498), .Y(n_497) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_440), .B(n_448), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B1(n_110), .B2(n_111), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_108), .B(n_147), .Y(n_528) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
XOR2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_437), .Y(n_111) );
INVx2_ASAP7_75t_L g467 ( .A(n_112), .Y(n_467) );
OR4x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_327), .C(n_374), .D(n_414), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_273), .C(n_302), .Y(n_113) );
AOI211xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_188), .B(n_226), .C(n_266), .Y(n_114) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_115), .A2(n_286), .B(n_303), .C(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_150), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_117), .B(n_265), .Y(n_264) );
INVx3_ASAP7_75t_SL g269 ( .A(n_117), .Y(n_269) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_117), .Y(n_281) );
AND2x4_ASAP7_75t_L g285 ( .A(n_117), .B(n_233), .Y(n_285) );
AND2x2_ASAP7_75t_L g296 ( .A(n_117), .B(n_173), .Y(n_296) );
OR2x2_ASAP7_75t_L g320 ( .A(n_117), .B(n_229), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_117), .B(n_234), .Y(n_333) );
AND2x2_ASAP7_75t_L g373 ( .A(n_117), .B(n_359), .Y(n_373) );
AND2x2_ASAP7_75t_L g380 ( .A(n_117), .B(n_343), .Y(n_380) );
AND2x2_ASAP7_75t_L g410 ( .A(n_117), .B(n_151), .Y(n_410) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_145), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_127), .C(n_140), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_119), .A2(n_175), .B(n_176), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_119), .A2(n_207), .B(n_208), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_119), .A2(n_168), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_119), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_119), .A2(n_559), .B(n_560), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
AND2x4_ASAP7_75t_L g158 ( .A(n_120), .B(n_124), .Y(n_158) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
INVx1_ASAP7_75t_L g257 ( .A(n_122), .Y(n_257) );
INVx1_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
INVx3_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_123), .Y(n_167) );
INVx1_ASAP7_75t_L g501 ( .A(n_123), .Y(n_501) );
BUFx3_ASAP7_75t_L g139 ( .A(n_124), .Y(n_139) );
INVx4_ASAP7_75t_SL g168 ( .A(n_124), .Y(n_168) );
INVx5_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx3_ASAP7_75t_L g184 ( .A(n_129), .Y(n_184) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_129), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_135), .C(n_137), .Y(n_131) );
OAI22xp33_ASAP7_75t_L g163 ( .A1(n_133), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_133), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_134), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_134), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_134), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx4_ASAP7_75t_L g239 ( .A(n_136), .Y(n_239) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_138), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_140), .A2(n_193), .B(n_200), .Y(n_192) );
INVx1_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_140), .A2(n_544), .B(n_550), .Y(n_543) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g149 ( .A(n_141), .B(n_142), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_147), .A2(n_174), .B(n_186), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_147), .B(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_148), .Y(n_216) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_148), .A2(n_497), .B(n_504), .Y(n_496) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_150), .B(n_337), .Y(n_349) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_172), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_151), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g287 ( .A(n_151), .B(n_172), .Y(n_287) );
BUFx3_ASAP7_75t_L g295 ( .A(n_151), .Y(n_295) );
OR2x2_ASAP7_75t_L g316 ( .A(n_151), .B(n_191), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_151), .B(n_337), .Y(n_427) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B(n_169), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_153), .A2(n_230), .B(n_231), .Y(n_229) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_153), .A2(n_558), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_154), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_155), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_155), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_155), .A2(n_509), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g230 ( .A(n_156), .Y(n_230) );
BUFx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_SL g159 ( .A1(n_160), .A2(n_161), .B(n_162), .C(n_168), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_161), .A2(n_168), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_SL g218 ( .A1(n_161), .A2(n_168), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_168), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_161), .A2(n_168), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_161), .A2(n_168), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_161), .A2(n_168), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_161), .A2(n_168), .B(n_546), .C(n_547), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_166), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_166), .B(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_166), .B(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_167), .A2(n_180), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
INVx1_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_171), .B(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_171), .A2(n_533), .B(n_540), .Y(n_532) );
AND2x2_ASAP7_75t_L g232 ( .A(n_172), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g280 ( .A(n_172), .Y(n_280) );
AND2x2_ASAP7_75t_L g343 ( .A(n_172), .B(n_234), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_172), .A2(n_346), .B1(n_348), .B2(n_350), .C(n_351), .Y(n_345) );
AND2x2_ASAP7_75t_L g359 ( .A(n_172), .B(n_229), .Y(n_359) );
AND2x2_ASAP7_75t_L g385 ( .A(n_172), .B(n_269), .Y(n_385) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g265 ( .A(n_173), .B(n_234), .Y(n_265) );
BUFx2_ASAP7_75t_L g399 ( .A(n_173), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_181), .C(n_182), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_179), .A2(n_182), .B(n_210), .C(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_182), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_182), .A2(n_562), .B(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g223 ( .A(n_184), .Y(n_223) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI32xp33_ASAP7_75t_L g365 ( .A1(n_189), .A2(n_326), .A3(n_340), .B1(n_366), .B2(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_201), .Y(n_189) );
AND2x2_ASAP7_75t_L g306 ( .A(n_190), .B(n_248), .Y(n_306) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g288 ( .A(n_191), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_191), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g360 ( .A(n_191), .B(n_248), .Y(n_360) );
AND2x2_ASAP7_75t_L g371 ( .A(n_191), .B(n_263), .Y(n_371) );
BUFx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g272 ( .A(n_192), .B(n_249), .Y(n_272) );
AND2x2_ASAP7_75t_L g276 ( .A(n_192), .B(n_249), .Y(n_276) );
AND2x2_ASAP7_75t_L g311 ( .A(n_192), .B(n_262), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_192), .B(n_214), .Y(n_318) );
OAI211xp5_ASAP7_75t_L g323 ( .A1(n_192), .A2(n_269), .B(n_280), .C(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g377 ( .A(n_192), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_192), .B(n_203), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_201), .B(n_260), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_201), .B(n_276), .Y(n_366) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g271 ( .A(n_202), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_214), .Y(n_202) );
AND2x2_ASAP7_75t_L g263 ( .A(n_203), .B(n_215), .Y(n_263) );
OR2x2_ASAP7_75t_L g278 ( .A(n_203), .B(n_215), .Y(n_278) );
AND2x2_ASAP7_75t_L g301 ( .A(n_203), .B(n_262), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_203), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_203), .B(n_261), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_203), .A2(n_289), .B1(n_335), .B2(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_203), .B(n_377), .Y(n_401) );
AND2x2_ASAP7_75t_L g416 ( .A(n_203), .B(n_276), .Y(n_416) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx3_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
AND2x2_ASAP7_75t_L g290 ( .A(n_204), .B(n_215), .Y(n_290) );
AND2x2_ASAP7_75t_L g292 ( .A(n_204), .B(n_248), .Y(n_292) );
AND3x2_ASAP7_75t_L g354 ( .A(n_204), .B(n_318), .C(n_355), .Y(n_354) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_212), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_205), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_205), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_205), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g389 ( .A(n_214), .B(n_261), .Y(n_389) );
INVx1_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g248 ( .A(n_215), .B(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_215), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_215), .B(n_260), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_215), .B(n_301), .C(n_377), .Y(n_429) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_224), .Y(n_215) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_216), .A2(n_235), .B(n_244), .Y(n_234) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_216), .A2(n_250), .B(n_258), .Y(n_249) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_225), .A2(n_478), .B(n_484), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_245), .B1(n_259), .B2(n_264), .Y(n_226) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_232), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_229), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g341 ( .A(n_229), .Y(n_341) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_232), .A2(n_358), .A3(n_359), .B(n_360), .Y(n_357) );
AND2x2_ASAP7_75t_L g382 ( .A(n_232), .B(n_269), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_232), .B(n_295), .Y(n_428) );
AND2x2_ASAP7_75t_L g337 ( .A(n_233), .B(n_269), .Y(n_337) );
AND2x2_ASAP7_75t_L g398 ( .A(n_233), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g268 ( .A(n_234), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g326 ( .A(n_234), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_239), .B(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_243), .Y(n_538) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_246), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_247), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AOI221x1_ASAP7_75t_SL g314 ( .A1(n_248), .A2(n_315), .B1(n_317), .B2(n_319), .C(n_321), .Y(n_314) );
INVx2_ASAP7_75t_L g262 ( .A(n_249), .Y(n_262) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_249), .Y(n_356) );
INVx2_ASAP7_75t_L g515 ( .A(n_256), .Y(n_515) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g344 ( .A(n_259), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_260), .B(n_277), .Y(n_369) );
INVx1_ASAP7_75t_SL g432 ( .A(n_260), .Y(n_432) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g350 ( .A(n_263), .B(n_276), .Y(n_350) );
INVx1_ASAP7_75t_L g418 ( .A(n_264), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_264), .B(n_347), .Y(n_431) );
INVx2_ASAP7_75t_SL g270 ( .A(n_265), .Y(n_270) );
AND2x2_ASAP7_75t_L g313 ( .A(n_265), .B(n_269), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_265), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_265), .B(n_340), .Y(n_367) );
AOI21xp33_ASAP7_75t_SL g266 ( .A1(n_267), .A2(n_270), .B(n_271), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_268), .B(n_340), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_268), .B(n_295), .Y(n_436) );
OR2x2_ASAP7_75t_L g308 ( .A(n_269), .B(n_287), .Y(n_308) );
AND2x2_ASAP7_75t_L g407 ( .A(n_269), .B(n_398), .Y(n_407) );
OAI22xp5_ASAP7_75t_SL g282 ( .A1(n_270), .A2(n_283), .B1(n_288), .B2(n_291), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_270), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g330 ( .A(n_272), .B(n_278), .Y(n_330) );
INVx1_ASAP7_75t_L g394 ( .A(n_272), .Y(n_394) );
AOI311xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_279), .A3(n_281), .B(n_282), .C(n_293), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_277), .A2(n_409), .B1(n_421), .B2(n_424), .C(n_426), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_277), .B(n_432), .Y(n_434) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
AOI211xp5_ASAP7_75t_L g321 ( .A1(n_280), .A2(n_322), .B(n_323), .C(n_325), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_SL g390 ( .A1(n_284), .A2(n_286), .B(n_391), .C(n_392), .Y(n_390) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_285), .B(n_359), .Y(n_425) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_288), .A2(n_308), .B1(n_309), .B2(n_312), .C(n_314), .Y(n_307) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g393 ( .A(n_290), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_294), .A2(n_352), .B(n_353), .C(n_357), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_295), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_295), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g317 ( .A(n_301), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_305), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g419 ( .A(n_308), .Y(n_419) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_311), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g346 ( .A(n_311), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g423 ( .A(n_311), .Y(n_423) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_340), .Y(n_364) );
INVx1_ASAP7_75t_SL g358 ( .A(n_320), .Y(n_358) );
INVx1_ASAP7_75t_L g335 ( .A(n_326), .Y(n_335) );
NAND3xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_345), .C(n_361), .Y(n_327) );
AOI322xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .A3(n_332), .B1(n_334), .B2(n_338), .C1(n_342), .C2(n_344), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_382), .B(n_383), .C(n_390), .Y(n_381) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_332), .A2(n_353), .B1(n_384), .B2(n_386), .Y(n_383) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g342 ( .A(n_340), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g379 ( .A(n_340), .B(n_380), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g430 ( .A1(n_340), .A2(n_431), .A3(n_432), .B1(n_433), .B2(n_435), .Y(n_430) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g352 ( .A(n_343), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_343), .A2(n_396), .B1(n_400), .B2(n_402), .C(n_405), .Y(n_395) );
AND2x2_ASAP7_75t_L g409 ( .A(n_343), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g412 ( .A(n_347), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g422 ( .A(n_347), .B(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g413 ( .A(n_356), .B(n_377), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B(n_365), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_378), .B(n_381), .C(n_395), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_389), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g404 ( .A(n_401), .Y(n_404) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_411), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_417), .B(n_420), .C(n_430), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp33_ASAP7_75t_L g754 ( .A(n_441), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g460 ( .A(n_443), .Y(n_460) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_444), .B(n_466), .Y(n_752) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
CKINVDCx6p67_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_454), .A2(n_455), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g755 ( .A(n_454), .B(n_456), .Y(n_755) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_743), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B1(n_468), .B2(n_470), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_466), .Y(n_469) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_665), .C(n_710), .Y(n_472) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_588), .C(n_629), .D(n_646), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_505), .B(n_519), .C(n_551), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_476), .B(n_506), .Y(n_505) );
NOR4xp25_ASAP7_75t_L g612 ( .A(n_476), .B(n_606), .C(n_613), .D(n_619), .Y(n_612) );
AND2x2_ASAP7_75t_L g685 ( .A(n_476), .B(n_574), .Y(n_685) );
AND2x2_ASAP7_75t_L g704 ( .A(n_476), .B(n_650), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_476), .B(n_699), .Y(n_713) );
AND2x2_ASAP7_75t_L g726 ( .A(n_476), .B(n_518), .Y(n_726) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g571 ( .A(n_477), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_477), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g628 ( .A(n_477), .B(n_486), .Y(n_628) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_477), .B(n_574), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_477), .B(n_486), .Y(n_643) );
AND2x2_ASAP7_75t_L g652 ( .A(n_477), .B(n_577), .Y(n_652) );
BUFx2_ASAP7_75t_L g675 ( .A(n_477), .Y(n_675) );
AND2x2_ASAP7_75t_L g679 ( .A(n_477), .B(n_496), .Y(n_679) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_496), .Y(n_518) );
BUFx2_ASAP7_75t_L g581 ( .A(n_486), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_486), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_613) );
OR2x2_ASAP7_75t_L g635 ( .A(n_486), .B(n_508), .Y(n_635) );
AND2x2_ASAP7_75t_L g699 ( .A(n_486), .B(n_577), .Y(n_699) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_508), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_487), .B(n_496), .Y(n_574) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_487), .Y(n_616) );
OR2x2_ASAP7_75t_L g651 ( .A(n_487), .B(n_507), .Y(n_651) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx3_ASAP7_75t_L g579 ( .A(n_496), .Y(n_579) );
BUFx2_ASAP7_75t_L g603 ( .A(n_496), .Y(n_603) );
AND2x2_ASAP7_75t_L g636 ( .A(n_496), .B(n_571), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_505), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_507), .B(n_579), .Y(n_583) );
INVx1_ASAP7_75t_L g611 ( .A(n_507), .Y(n_611) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g577 ( .A(n_508), .Y(n_577) );
INVx1_ASAP7_75t_L g589 ( .A(n_518), .Y(n_589) );
NAND2x1_ASAP7_75t_SL g519 ( .A(n_520), .B(n_529), .Y(n_519) );
AND2x2_ASAP7_75t_L g587 ( .A(n_520), .B(n_542), .Y(n_587) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_520), .Y(n_661) );
AND2x2_ASAP7_75t_L g688 ( .A(n_520), .B(n_608), .Y(n_688) );
AND2x2_ASAP7_75t_L g696 ( .A(n_520), .B(n_658), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_520), .B(n_554), .Y(n_723) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g555 ( .A(n_521), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_521), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
INVx1_ASAP7_75t_L g599 ( .A(n_521), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_521), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g632 ( .A(n_521), .B(n_557), .Y(n_632) );
OR2x2_ASAP7_75t_L g670 ( .A(n_521), .B(n_625), .Y(n_670) );
AOI32xp33_ASAP7_75t_L g682 ( .A1(n_521), .A2(n_683), .A3(n_686), .B1(n_687), .B2(n_688), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_521), .B(n_658), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_521), .B(n_618), .Y(n_733) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g644 ( .A(n_530), .B(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
INVx1_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
AND2x2_ASAP7_75t_L g608 ( .A(n_531), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_531), .B(n_556), .Y(n_625) );
AND2x2_ASAP7_75t_L g658 ( .A(n_531), .B(n_634), .Y(n_658) );
AND2x2_ASAP7_75t_L g695 ( .A(n_531), .B(n_557), .Y(n_695) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g554 ( .A(n_532), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_532), .B(n_556), .Y(n_585) );
AND2x2_ASAP7_75t_L g592 ( .A(n_532), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g633 ( .A(n_532), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B(n_538), .Y(n_535) );
INVx2_ASAP7_75t_L g609 ( .A(n_542), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_542), .B(n_556), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_542), .B(n_600), .Y(n_681) );
INVx1_ASAP7_75t_L g703 ( .A(n_542), .Y(n_703) );
INVx1_ASAP7_75t_L g720 ( .A(n_542), .Y(n_720) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g573 ( .A(n_543), .B(n_556), .Y(n_573) );
AND2x2_ASAP7_75t_L g595 ( .A(n_543), .B(n_557), .Y(n_595) );
INVx1_ASAP7_75t_L g634 ( .A(n_543), .Y(n_634) );
AOI221x1_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_566), .B1(n_572), .B2(n_574), .C(n_575), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_552), .A2(n_639), .B1(n_706), .B2(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g597 ( .A(n_553), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g692 ( .A(n_553), .B(n_572), .Y(n_692) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g648 ( .A(n_554), .B(n_573), .Y(n_648) );
INVx1_ASAP7_75t_L g660 ( .A(n_555), .Y(n_660) );
AND2x2_ASAP7_75t_L g671 ( .A(n_555), .B(n_658), .Y(n_671) );
AND2x2_ASAP7_75t_L g738 ( .A(n_555), .B(n_633), .Y(n_738) );
INVx2_ASAP7_75t_L g600 ( .A(n_556), .Y(n_600) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_567), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g690 ( .A(n_567), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_568), .B(n_651), .Y(n_654) );
INVx3_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_569), .A2(n_690), .B(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_572), .B(n_598), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_573), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g664 ( .A(n_573), .B(n_592), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_573), .B(n_599), .Y(n_741) );
AND2x2_ASAP7_75t_L g610 ( .A(n_574), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g677 ( .A(n_574), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_580), .B(n_584), .Y(n_575) );
NAND2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_577), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g626 ( .A(n_577), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g638 ( .A(n_577), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_577), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g662 ( .A(n_578), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_578), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_578), .B(n_581), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_581), .A2(n_620), .B(n_650), .C(n_652), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_581), .A2(n_668), .B1(n_671), .B2(n_672), .C(n_676), .Y(n_667) );
AND2x2_ASAP7_75t_L g663 ( .A(n_582), .B(n_616), .Y(n_663) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g623 ( .A(n_587), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g694 ( .A(n_587), .B(n_695), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_596), .C(n_621), .Y(n_588) );
NAND3xp33_ASAP7_75t_SL g707 ( .A(n_589), .B(n_708), .C(n_709), .Y(n_707) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
OR2x2_ASAP7_75t_L g680 ( .A(n_591), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B1(n_604), .B2(n_610), .C(n_612), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_598), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g620 ( .A(n_603), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_603), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
OR2x2_ASAP7_75t_L g740 ( .A(n_603), .B(n_651), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVxp67_ASAP7_75t_L g714 ( .A(n_606), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_608), .B(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g615 ( .A(n_609), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_611), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_611), .B(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_611), .B(n_678), .Y(n_717) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_615), .Y(n_641) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g731 ( .A(n_620), .B(n_651), .Y(n_731) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g709 ( .A(n_626), .Y(n_709) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI322xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_635), .A3(n_636), .B1(n_637), .B2(n_640), .C1(n_642), .C2(n_644), .Y(n_629) );
OAI322xp33_ASAP7_75t_L g711 ( .A1(n_630), .A2(n_712), .A3(n_713), .B1(n_714), .B2(n_715), .C1(n_716), .C2(n_718), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx4_ASAP7_75t_L g645 ( .A(n_632), .Y(n_645) );
AND2x2_ASAP7_75t_L g706 ( .A(n_632), .B(n_658), .Y(n_706) );
AND2x2_ASAP7_75t_L g719 ( .A(n_632), .B(n_720), .Y(n_719) );
CKINVDCx16_ASAP7_75t_R g730 ( .A(n_635), .Y(n_730) );
INVx1_ASAP7_75t_L g708 ( .A(n_636), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g642 ( .A(n_638), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g725 ( .A(n_638), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_638), .B(n_679), .Y(n_736) );
OR2x2_ASAP7_75t_L g669 ( .A(n_641), .B(n_670), .Y(n_669) );
INVxp33_ASAP7_75t_L g686 ( .A(n_641), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_653), .C(n_655), .Y(n_646) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_645), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g729 ( .A(n_645), .Y(n_729) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_677), .A3(n_694), .B1(n_696), .B2(n_697), .C1(n_700), .C2(n_704), .Y(n_693) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_663), .B2(n_664), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_689), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_682), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_670), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp33_ASAP7_75t_SL g687 ( .A(n_673), .B(n_684), .Y(n_687) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI322xp33_ASAP7_75t_L g727 ( .A1(n_675), .A2(n_728), .A3(n_730), .B1(n_731), .B2(n_732), .C1(n_734), .C2(n_737), .Y(n_727) );
AOI21xp33_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_685), .B(n_733), .Y(n_742) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_691), .B(n_693), .C(n_705), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR4xp25_ASAP7_75t_L g710 ( .A(n_711), .B(n_721), .C(n_727), .D(n_739), .Y(n_710) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx14_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_744), .Y(n_751) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
endmodule