module fake_jpeg_9562_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_10),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_36),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_33),
.B(n_28),
.C(n_26),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_27),
.CON(n_56),
.SN(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_32),
.B1(n_35),
.B2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_23),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_18),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_26),
.C(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_67),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_40),
.C(n_42),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_74),
.C(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_32),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_40),
.C(n_51),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_16),
.B1(n_19),
.B2(n_27),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_0),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_40),
.C(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_16),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_38),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_40),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_83),
.B1(n_73),
.B2(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_38),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_1),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_88),
.B(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_109),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_79),
.C(n_65),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_111),
.C(n_121),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_35),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_77),
.B(n_69),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_120),
.B(n_24),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_90),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.C(n_11),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_122),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_30),
.B(n_2),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_30),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_30),
.C(n_8),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_104),
.C(n_86),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_134),
.C(n_135),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_104),
.B(n_3),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_83),
.B1(n_70),
.B2(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_112),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_112),
.B(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_116),
.B1(n_114),
.B2(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_15),
.A3(n_14),
.B1(n_12),
.B2(n_4),
.C(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_12),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_131),
.C(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_131),
.C(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_132),
.B(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_169),
.C(n_75),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_153),
.B(n_143),
.Y(n_167)
);

AOI311xp33_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_159),
.A3(n_125),
.B(n_118),
.C(n_15),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_149),
.C(n_143),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_160),
.B(n_161),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_172),
.C(n_174),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_170),
.C(n_100),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_95),
.B(n_4),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule