module fake_netlist_6_3292_n_888 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_888);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_888;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_41),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_60),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_136),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_53),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_108),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_77),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_71),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_28),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_98),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_37),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_147),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_26),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_5),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_54),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_55),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_69),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_82),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_63),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_66),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_111),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_176),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_130),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_75),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_106),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_165),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_116),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_172),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_89),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_195),
.B(n_22),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_23),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_0),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_189),
.B(n_24),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_0),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_204),
.B(n_1),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_229),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_215),
.A2(n_2),
.B(n_3),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_245),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_233),
.A2(n_234),
.B(n_187),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_193),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_197),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_232),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_205),
.B(n_208),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_191),
.B(n_6),
.Y(n_303)
);

CKINVDCx6p67_ASAP7_75t_R g304 ( 
.A(n_200),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

NOR2x1p5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_190),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_252),
.B1(n_199),
.B2(n_251),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_7),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_269),
.B(n_202),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_207),
.C(n_206),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_291),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_211),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_288),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_270),
.B(n_219),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_216),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_261),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_261),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_270),
.B(n_220),
.Y(n_341)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_264),
.A2(n_221),
.B(n_217),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_270),
.B(n_222),
.Y(n_343)
);

AO21x2_ASAP7_75t_L g344 ( 
.A1(n_276),
.A2(n_231),
.B(n_225),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_288),
.Y(n_345)
);

AO22x2_ASAP7_75t_L g346 ( 
.A1(n_256),
.A2(n_253),
.B1(n_246),
.B2(n_243),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_256),
.B(n_224),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_267),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_304),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_260),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_L g357 ( 
.A(n_275),
.B(n_226),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_256),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_356),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_356),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_268),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_311),
.B(n_303),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_292),
.B(n_305),
.C(n_300),
.Y(n_367)
);

NAND2x1_ASAP7_75t_L g368 ( 
.A(n_319),
.B(n_268),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_268),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_298),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_302),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_257),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_302),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_302),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_257),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_257),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_265),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_265),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_344),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_315),
.B(n_265),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_322),
.B(n_331),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_266),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_321),
.A2(n_305),
.B1(n_258),
.B2(n_259),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_266),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_312),
.B(n_235),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_314),
.B(n_266),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_299),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_316),
.B(n_236),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_338),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_299),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_299),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_299),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_306),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_313),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_306),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_299),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_342),
.B(n_238),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_349),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_287),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_307),
.A2(n_227),
.B1(n_230),
.B2(n_237),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_292),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_353),
.B(n_267),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_L g424 ( 
.A(n_325),
.B(n_239),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_325),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_282),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_326),
.B(n_278),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_373),
.A2(n_351),
.B(n_335),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_329),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_281),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_358),
.A2(n_242),
.B1(n_281),
.B2(n_241),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_351),
.B(n_335),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_367),
.B(n_412),
.C(n_391),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_370),
.A2(n_259),
.B(n_258),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_329),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_392),
.B(n_352),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_362),
.B(n_360),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_374),
.B(n_412),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_363),
.B(n_287),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_287),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_384),
.B(n_287),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_393),
.B(n_304),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_351),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_397),
.B(n_262),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_351),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_383),
.A2(n_280),
.B(n_278),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_418),
.A2(n_264),
.B(n_274),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_366),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_274),
.B(n_240),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_416),
.A2(n_248),
.B(n_249),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_250),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_290),
.B(n_280),
.Y(n_465)
);

BUFx8_ASAP7_75t_SL g466 ( 
.A(n_402),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_369),
.B(n_272),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

O2A1O1Ixp5_ASAP7_75t_L g469 ( 
.A1(n_416),
.A2(n_279),
.B(n_272),
.C(n_283),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_406),
.A2(n_279),
.B(n_272),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_389),
.A2(n_278),
.B(n_290),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_395),
.B(n_277),
.C(n_345),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_390),
.A2(n_280),
.B(n_278),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_367),
.A2(n_262),
.B(n_263),
.C(n_279),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_397),
.B(n_283),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_399),
.B(n_283),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_404),
.B(n_263),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_393),
.A2(n_345),
.B(n_328),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_365),
.A2(n_290),
.B(n_280),
.C(n_278),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_417),
.A2(n_328),
.B(n_290),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_371),
.B(n_280),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_420),
.B(n_286),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_395),
.B(n_286),
.Y(n_486)
);

NOR2x1_ASAP7_75t_SL g487 ( 
.A(n_378),
.B(n_409),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_375),
.A2(n_290),
.B1(n_96),
.B2(n_100),
.Y(n_488)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_400),
.A2(n_10),
.B(n_11),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_407),
.A2(n_94),
.B(n_184),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_408),
.A2(n_93),
.B(n_183),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_25),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_414),
.A2(n_95),
.B(n_182),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_398),
.B(n_10),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_401),
.B(n_11),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_422),
.A2(n_101),
.B(n_181),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_27),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_413),
.B(n_29),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_372),
.A2(n_102),
.B(n_178),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_439),
.A2(n_423),
.B(n_400),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_436),
.A2(n_386),
.B(n_385),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_458),
.A2(n_409),
.B(n_380),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_447),
.A2(n_409),
.B(n_377),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_448),
.A2(n_403),
.B(n_427),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_429),
.A2(n_403),
.B(n_409),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_30),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_450),
.A2(n_185),
.B(n_92),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_452),
.A2(n_456),
.B(n_443),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_455),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_514)
);

AOI21x1_ASAP7_75t_L g515 ( 
.A1(n_430),
.A2(n_103),
.B(n_174),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_500),
.A2(n_90),
.B(n_173),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_31),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_499),
.A2(n_88),
.B(n_169),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_449),
.A2(n_177),
.B(n_87),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_12),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_14),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_449),
.A2(n_167),
.B(n_105),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_460),
.A2(n_163),
.B(n_86),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_454),
.B(n_15),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_487),
.A2(n_83),
.B(n_161),
.Y(n_526)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_32),
.Y(n_527)
);

AOI21xp33_ASAP7_75t_L g528 ( 
.A1(n_461),
.A2(n_15),
.B(n_16),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_460),
.A2(n_162),
.B(n_107),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_33),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_34),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_466),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_475),
.A2(n_160),
.B(n_109),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_464),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_468),
.A2(n_81),
.B(n_153),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_486),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_468),
.A2(n_110),
.B(n_152),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_453),
.A2(n_79),
.B(n_151),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_479),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_459),
.B(n_78),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_475),
.A2(n_112),
.B(n_149),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_470),
.A2(n_76),
.B(n_148),
.Y(n_542)
);

CKINVDCx8_ASAP7_75t_R g543 ( 
.A(n_432),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_454),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_494),
.B(n_74),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_455),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_469),
.A2(n_72),
.B(n_146),
.Y(n_547)
);

OAI21x1_ASAP7_75t_SL g548 ( 
.A1(n_489),
.A2(n_70),
.B(n_145),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_453),
.A2(n_68),
.B(n_144),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_434),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_65),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_17),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_453),
.A2(n_113),
.B(n_143),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_455),
.A2(n_64),
.B(n_142),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_498),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_442),
.B(n_62),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_457),
.A2(n_115),
.B(n_141),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_484),
.A2(n_473),
.B(n_471),
.Y(n_560)
);

AO31x2_ASAP7_75t_L g561 ( 
.A1(n_482),
.A2(n_19),
.A3(n_20),
.B(n_36),
.Y(n_561)
);

BUFx2_ASAP7_75t_SL g562 ( 
.A(n_544),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_433),
.Y(n_563)
);

OAI211xp5_ASAP7_75t_L g564 ( 
.A1(n_528),
.A2(n_485),
.B(n_496),
.C(n_495),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_505),
.A2(n_492),
.B(n_493),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_503),
.A2(n_462),
.B(n_478),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_444),
.Y(n_568)
);

AO222x2_ASAP7_75t_L g569 ( 
.A1(n_552),
.A2(n_19),
.B1(n_20),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_476),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_519),
.Y(n_571)
);

AO21x2_ASAP7_75t_L g572 ( 
.A1(n_503),
.A2(n_491),
.B(n_490),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

AOI21xp33_ASAP7_75t_L g574 ( 
.A1(n_528),
.A2(n_488),
.B(n_463),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_480),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_513),
.B(n_546),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_525),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_508),
.A2(n_465),
.B(n_501),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_522),
.A2(n_480),
.B1(n_476),
.B2(n_497),
.Y(n_579)
);

OAI21x1_ASAP7_75t_SL g580 ( 
.A1(n_548),
.A2(n_480),
.B(n_45),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_553),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_536),
.B(n_476),
.C(n_480),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_531),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_546),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_508),
.A2(n_42),
.B(n_46),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_512),
.B(n_47),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_546),
.B(n_48),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_556),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_504),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_534),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_49),
.Y(n_593)
);

OAI21x1_ASAP7_75t_SL g594 ( 
.A1(n_510),
.A2(n_51),
.B(n_52),
.Y(n_594)
);

OAI21x1_ASAP7_75t_SL g595 ( 
.A1(n_510),
.A2(n_57),
.B(n_58),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_540),
.Y(n_596)
);

AO21x1_ASAP7_75t_L g597 ( 
.A1(n_530),
.A2(n_59),
.B(n_61),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_532),
.B(n_117),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_517),
.A2(n_119),
.B(n_120),
.Y(n_599)
);

BUFx2_ASAP7_75t_SL g600 ( 
.A(n_526),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_540),
.Y(n_601)
);

INVx3_ASAP7_75t_SL g602 ( 
.A(n_514),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_560),
.A2(n_121),
.B(n_122),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_506),
.A2(n_123),
.B(n_125),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_507),
.A2(n_126),
.B(n_128),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_545),
.B(n_154),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_530),
.A2(n_129),
.B(n_131),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_545),
.B(n_135),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_557),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_610)
);

OAI21x1_ASAP7_75t_SL g611 ( 
.A1(n_542),
.A2(n_547),
.B(n_517),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

OAI21x1_ASAP7_75t_SL g614 ( 
.A1(n_542),
.A2(n_547),
.B(n_551),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_585),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_571),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_590),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_589),
.Y(n_619)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_613),
.A2(n_551),
.B(n_515),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_602),
.B(n_561),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

BUFx2_ASAP7_75t_SL g623 ( 
.A(n_585),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_577),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_585),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_514),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_612),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_566),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

AO21x1_ASAP7_75t_SL g632 ( 
.A1(n_574),
.A2(n_561),
.B(n_541),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_611),
.A2(n_523),
.B(n_533),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_592),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_586),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_581),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_568),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_602),
.B(n_561),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_565),
.A2(n_529),
.B(n_524),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_583),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_593),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_586),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_563),
.A2(n_554),
.B1(n_549),
.B2(n_538),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_563),
.A2(n_535),
.B1(n_537),
.B2(n_555),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_587),
.A2(n_518),
.B(n_511),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_574),
.A2(n_520),
.B1(n_558),
.B2(n_516),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_584),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_576),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_596),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_570),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_570),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_567),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_576),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_596),
.A2(n_582),
.B1(n_564),
.B2(n_607),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_626),
.B(n_599),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_656),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_599),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_619),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_588),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_564),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_640),
.B(n_588),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_640),
.B(n_607),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_614),
.B1(n_610),
.B2(n_569),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_656),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_617),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_619),
.B(n_567),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_659),
.B(n_609),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_659),
.B(n_572),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_639),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_653),
.B(n_562),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_618),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_627),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_639),
.A2(n_610),
.B1(n_569),
.B2(n_597),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_624),
.B(n_598),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_645),
.B(n_608),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_638),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_628),
.B(n_608),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_654),
.B(n_616),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_658),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_646),
.B(n_604),
.C(n_579),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_645),
.B(n_572),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_652),
.B(n_604),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_652),
.B(n_594),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_654),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_637),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_635),
.B(n_578),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_637),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_627),
.Y(n_697)
);

OAI222xp33_ASAP7_75t_L g698 ( 
.A1(n_618),
.A2(n_630),
.B1(n_634),
.B2(n_642),
.C1(n_629),
.C2(n_647),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_630),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_655),
.B(n_578),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_644),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_636),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_627),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_650),
.B(n_600),
.Y(n_705)
);

OAI21xp33_ASAP7_75t_L g706 ( 
.A1(n_629),
.A2(n_580),
.B(n_595),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_578),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_627),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_615),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_651),
.A2(n_623),
.B1(n_660),
.B2(n_657),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_657),
.B(n_651),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_651),
.B(n_615),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_632),
.A2(n_631),
.B1(n_633),
.B2(n_649),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_625),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_665),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_701),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_665),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_676),
.B(n_625),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_670),
.A2(n_632),
.B1(n_631),
.B2(n_633),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_676),
.B(n_631),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_672),
.B(n_623),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_681),
.A2(n_622),
.B1(n_636),
.B2(n_633),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_669),
.B(n_633),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_667),
.B(n_622),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_701),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_669),
.B(n_622),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_711),
.B(n_641),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_666),
.B(n_620),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_648),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_694),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_699),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_679),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_663),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_711),
.B(n_641),
.Y(n_737)
);

INVxp33_ASAP7_75t_L g738 ( 
.A(n_682),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_663),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_671),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_666),
.B(n_620),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_671),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_687),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_668),
.B(n_648),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_687),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_668),
.B(n_712),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_684),
.B(n_677),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_709),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_712),
.B(n_715),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_678),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_705),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_700),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_708),
.B(n_713),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_680),
.B(n_708),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_694),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_700),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_688),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_674),
.B(n_685),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_713),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_680),
.B(n_697),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_730),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_755),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_751),
.B(n_683),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_751),
.B(n_698),
.C(n_706),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_736),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_746),
.B(n_664),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_739),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_749),
.B(n_664),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_738),
.A2(n_689),
.B1(n_706),
.B2(n_683),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_728),
.B(n_673),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_724),
.B(n_675),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_716),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_759),
.B(n_674),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_740),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_742),
.Y(n_778)
);

NOR2x1p5_ASAP7_75t_L g779 ( 
.A(n_747),
.B(n_725),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_728),
.B(n_673),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_728),
.B(n_707),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_738),
.B(n_690),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_754),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_752),
.B(n_675),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_743),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_737),
.B(n_707),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_753),
.B(n_690),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_745),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_753),
.B(n_662),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_757),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_734),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_748),
.B(n_662),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_719),
.B(n_691),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_733),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_737),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_766),
.B(n_752),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_763),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_793),
.B(n_756),
.Y(n_800)
);

NAND2xp67_ASAP7_75t_SL g801 ( 
.A(n_795),
.B(n_741),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_764),
.Y(n_802)
);

NAND2x1p5_ASAP7_75t_L g803 ( 
.A(n_796),
.B(n_721),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_792),
.B(n_756),
.Y(n_804)
);

OAI21xp33_ASAP7_75t_L g805 ( 
.A1(n_767),
.A2(n_720),
.B(n_744),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_767),
.B(n_722),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_775),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_789),
.B(n_731),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_797),
.B(n_737),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_782),
.B(n_733),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_779),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_772),
.B(n_748),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_775),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_794),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_774),
.B(n_727),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_768),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_770),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_794),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_776),
.B(n_732),
.Y(n_819)
);

OAI211xp5_ASAP7_75t_SL g820 ( 
.A1(n_806),
.A2(n_772),
.B(n_720),
.C(n_783),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_808),
.B(n_773),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_815),
.B(n_798),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_819),
.B(n_783),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_819),
.B(n_771),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_812),
.A2(n_710),
.B1(n_689),
.B2(n_692),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_807),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_813),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_803),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_799),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_802),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_816),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_809),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_798),
.B(n_769),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_800),
.B(n_785),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_825),
.A2(n_805),
.B(n_811),
.Y(n_835)
);

XOR2x2_ASAP7_75t_L g836 ( 
.A(n_824),
.B(n_750),
.Y(n_836)
);

AOI32xp33_ASAP7_75t_L g837 ( 
.A1(n_820),
.A2(n_809),
.A3(n_817),
.B1(n_800),
.B2(n_797),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_828),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_823),
.B(n_803),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_L g840 ( 
.A(n_822),
.B(n_810),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_829),
.Y(n_841)
);

AOI211xp5_ASAP7_75t_SL g842 ( 
.A1(n_835),
.A2(n_825),
.B(n_723),
.C(n_834),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_837),
.A2(n_834),
.B(n_810),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_SL g844 ( 
.A1(n_838),
.A2(n_828),
.B(n_832),
.C(n_831),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_839),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_833),
.B1(n_830),
.B2(n_773),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_841),
.B(n_821),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_843),
.A2(n_836),
.B1(n_786),
.B2(n_781),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_842),
.A2(n_804),
.B(n_827),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_844),
.A2(n_804),
.B(n_826),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_846),
.B(n_773),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_845),
.B(n_818),
.Y(n_852)
);

NOR2x1_ASAP7_75t_L g853 ( 
.A(n_851),
.B(n_847),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_848),
.B(n_788),
.C(n_777),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_849),
.B(n_791),
.C(n_790),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_852),
.C(n_850),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_855),
.Y(n_857)
);

NOR2x1_ASAP7_75t_L g858 ( 
.A(n_854),
.B(n_801),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_857),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

XNOR2x1_ASAP7_75t_L g861 ( 
.A(n_858),
.B(n_692),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_857),
.Y(n_862)
);

NAND4xp75_ASAP7_75t_L g863 ( 
.A(n_857),
.B(n_691),
.C(n_778),
.D(n_761),
.Y(n_863)
);

XNOR2xp5_ASAP7_75t_L g864 ( 
.A(n_860),
.B(n_862),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_863),
.A2(n_780),
.B1(n_814),
.B2(n_786),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_861),
.B(n_762),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_861),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_864),
.Y(n_869)
);

OAI22x1_ASAP7_75t_L g870 ( 
.A1(n_868),
.A2(n_760),
.B1(n_679),
.B2(n_704),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_865),
.Y(n_871)
);

AOI21x1_ASAP7_75t_L g872 ( 
.A1(n_867),
.A2(n_692),
.B(n_762),
.Y(n_872)
);

OA22x2_ASAP7_75t_L g873 ( 
.A1(n_869),
.A2(n_866),
.B1(n_760),
.B2(n_692),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_871),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_870),
.B(n_679),
.C(n_704),
.Y(n_875)
);

AOI22x1_ASAP7_75t_L g876 ( 
.A1(n_872),
.A2(n_697),
.B1(n_704),
.B2(n_765),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_SL g877 ( 
.A1(n_869),
.A2(n_697),
.B1(n_781),
.B2(n_786),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_874),
.B(n_735),
.Y(n_878)
);

AO22x2_ASAP7_75t_L g879 ( 
.A1(n_875),
.A2(n_735),
.B1(n_765),
.B2(n_780),
.Y(n_879)
);

INVx5_ASAP7_75t_SL g880 ( 
.A(n_877),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_873),
.B(n_780),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_880),
.A2(n_876),
.B1(n_781),
.B2(n_787),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_878),
.A2(n_703),
.B(n_714),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_881),
.B(n_784),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_882),
.A2(n_879),
.B(n_703),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_885),
.Y(n_886)
);

AOI221xp5_ASAP7_75t_L g887 ( 
.A1(n_886),
.A2(n_884),
.B1(n_883),
.B2(n_717),
.C(n_726),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_887),
.A2(n_696),
.B1(n_702),
.B2(n_695),
.Y(n_888)
);


endmodule