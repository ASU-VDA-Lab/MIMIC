module real_jpeg_25614_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_60),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_38),
.C(n_79),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_2),
.A2(n_61),
.B1(n_65),
.B2(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_123),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_2),
.A2(n_38),
.B1(n_40),
.B2(n_197),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_2),
.B(n_26),
.C(n_43),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_2),
.A2(n_25),
.B(n_258),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_56),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_61),
.B1(n_65),
.B2(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_5),
.A2(n_38),
.B1(n_40),
.B2(n_107),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_107),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_61),
.B1(n_65),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_38),
.B1(n_40),
.B2(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_54),
.B1(n_57),
.B2(n_83),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_83),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_54),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_61),
.B1(n_65),
.B2(n_70),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_8),
.A2(n_38),
.B1(n_40),
.B2(n_70),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_70),
.Y(n_228)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_37),
.B1(n_61),
.B2(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_38),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_47),
.B1(n_61),
.B2(n_65),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_12),
.A2(n_38),
.B1(n_40),
.B2(n_58),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_58),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_71),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_14),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_61),
.B1(n_65),
.B2(n_145),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_38),
.B1(n_40),
.B2(n_145),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_145),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_21),
.B(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_22),
.A2(n_74),
.B1(n_75),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_22),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_51),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_24),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_25),
.A2(n_31),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_25),
.A2(n_28),
.B1(n_95),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_27),
.B1(n_170),
.B2(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_25),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_29),
.B(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_30),
.B(n_197),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_32),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_41),
.B1(n_48),
.B2(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_40),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_38),
.B(n_265),
.Y(n_264)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_48),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_41),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_41),
.A2(n_48),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_45),
.A2(n_86),
.B1(n_101),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_45),
.A2(n_156),
.B(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_45),
.A2(n_193),
.B(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_45),
.B(n_197),
.Y(n_277)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_48),
.B(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_59),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_66),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_55),
.A2(n_63),
.A3(n_65),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_69),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_59),
.A2(n_67),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_72),
.B1(n_106),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_65),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_61),
.B(n_66),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_61),
.B(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_71),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_72),
.A2(n_111),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_85),
.B(n_89),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_77),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_77),
.A2(n_165),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_103),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_78),
.A2(n_149),
.B(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_86),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_86),
.A2(n_246),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_88),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_90),
.A2(n_91),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.C(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_92),
.A2(n_93),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_97),
.A2(n_154),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_102),
.B(n_104),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_122),
.A2(n_123),
.B1(n_164),
.B2(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_150),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_307),
.B(n_313),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_182),
.B(n_306),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_175),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_138),
.B(n_175),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_157),
.C(n_159),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_139),
.A2(n_140),
.B1(n_157),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_147),
.C(n_151),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_155),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_159),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_162),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_171),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_168),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_177),
.B(n_178),
.C(n_181),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_213),
.B(n_300),
.C(n_305),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_207),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_199),
.C(n_200),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_185),
.A2(n_186),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_199),
.B(n_200),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_294),
.B(n_299),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_247),
.B(n_293),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_236),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_218),
.B(n_236),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.C(n_233),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B(n_227),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_270),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_229),
.A2(n_233),
.B1(n_234),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_243),
.C(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_287),
.B(n_292),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_266),
.B(n_286),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_260),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_275),
.B(n_285),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_273),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_280),
.B(n_284),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_291),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_298),
.Y(n_299)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);


endmodule