module fake_jpeg_31399_n_447 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_49),
.Y(n_135)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_51),
.B(n_71),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_78),
.Y(n_105)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_0),
.CON(n_63),
.SN(n_63)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_16),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_14),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_90),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_22),
.B(n_0),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_77),
.B1(n_53),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_92),
.A2(n_102),
.B1(n_118),
.B2(n_126),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_93),
.B(n_104),
.Y(n_187)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_94),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_24),
.B(n_33),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_24),
.B1(n_17),
.B2(n_18),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_43),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_124),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_35),
.C(n_40),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_99),
.C(n_116),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_132),
.B1(n_27),
.B2(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_69),
.B(n_43),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_136),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_46),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_54),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_62),
.B1(n_61),
.B2(n_59),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_25),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_85),
.B(n_26),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_33),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_26),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_142),
.B(n_4),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_130),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_147),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_74),
.B1(n_40),
.B2(n_35),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_149),
.A2(n_193),
.B1(n_131),
.B2(n_91),
.Y(n_219)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_155),
.B(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_17),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_157),
.B(n_184),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_159),
.A2(n_176),
.B1(n_185),
.B2(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_36),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_100),
.C(n_128),
.Y(n_213)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

OA22x2_ASAP7_75t_SL g164 ( 
.A1(n_92),
.A2(n_139),
.B1(n_135),
.B2(n_132),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_178),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_111),
.A2(n_57),
.B1(n_55),
.B2(n_32),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_197),
.B(n_113),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_23),
.B1(n_22),
.B2(n_36),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_105),
.A2(n_23),
.B(n_32),
.C(n_2),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_118),
.B(n_32),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_179),
.A2(n_109),
.B1(n_108),
.B2(n_13),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_188),
.Y(n_231)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_189),
.B(n_7),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_32),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_123),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_123),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_96),
.A2(n_0),
.B(n_4),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_192),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_140),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_6),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_140),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_121),
.B(n_6),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_125),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_159),
.B1(n_172),
.B2(n_196),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_201),
.A2(n_234),
.B(n_238),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_214),
.B1(n_222),
.B2(n_236),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_189),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_128),
.B1(n_131),
.B2(n_91),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_157),
.B(n_100),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_215),
.B(n_226),
.C(n_166),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_227),
.B1(n_202),
.B2(n_212),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_164),
.A2(n_138),
.B1(n_127),
.B2(n_144),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_109),
.B(n_144),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_150),
.B(n_188),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_109),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_175),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_170),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_164),
.A2(n_127),
.B1(n_138),
.B2(n_108),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_155),
.A2(n_108),
.B1(n_10),
.B2(n_11),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_165),
.B1(n_146),
.B2(n_197),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_161),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_246),
.A2(n_264),
.B1(n_202),
.B2(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_208),
.B(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_248),
.B(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_184),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_255),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_175),
.B(n_149),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_270),
.B1(n_277),
.B2(n_252),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_253),
.B(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_187),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_167),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_217),
.B(n_177),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_280),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_268),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_209),
.A2(n_191),
.B(n_180),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_263),
.A2(n_264),
.B(n_273),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_204),
.A2(n_158),
.B(n_195),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_169),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_272),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_201),
.A2(n_175),
.B1(n_162),
.B2(n_152),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_274),
.B1(n_278),
.B2(n_244),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_207),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_194),
.Y(n_268)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_204),
.A2(n_181),
.B(n_168),
.C(n_171),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_232),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_223),
.A2(n_151),
.B(n_153),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_227),
.A2(n_215),
.B1(n_236),
.B2(n_206),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_239),
.A2(n_182),
.B1(n_228),
.B2(n_232),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_217),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_228),
.A2(n_230),
.B(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_205),
.B(n_231),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_284),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_215),
.A2(n_230),
.B1(n_214),
.B2(n_226),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_200),
.B1(n_211),
.B2(n_225),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_218),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_242),
.Y(n_311)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_234),
.C(n_211),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_295),
.Y(n_324)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_312),
.B1(n_266),
.B2(n_278),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_303),
.A2(n_263),
.B(n_262),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_200),
.C(n_243),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_307),
.C(n_315),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_242),
.Y(n_307)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_311),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_252),
.A2(n_244),
.B1(n_233),
.B2(n_221),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_283),
.B1(n_277),
.B2(n_250),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_229),
.C(n_216),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_279),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_249),
.B(n_207),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_343),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_281),
.C(n_257),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_331),
.C(n_335),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_247),
.B(n_274),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_329),
.A2(n_310),
.B(n_295),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_268),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_350),
.B1(n_299),
.B2(n_316),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_279),
.B(n_268),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_310),
.B(n_289),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_255),
.C(n_267),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_318),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_345),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_247),
.C(n_262),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_341),
.C(n_348),
.Y(n_356)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_250),
.A3(n_248),
.B1(n_286),
.B2(n_270),
.Y(n_339)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_250),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_295),
.A2(n_254),
.B1(n_269),
.B2(n_221),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_297),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_347),
.B(n_349),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_216),
.C(n_254),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_304),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_300),
.A2(n_269),
.B1(n_256),
.B2(n_271),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_289),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_360),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_352),
.A2(n_361),
.B1(n_367),
.B2(n_368),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_353),
.A2(n_363),
.B(n_328),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_275),
.C(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_359),
.A2(n_372),
.B(n_334),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_315),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_324),
.A2(n_295),
.B1(n_321),
.B2(n_301),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_310),
.B(n_308),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_290),
.C(n_312),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_369),
.C(n_371),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_324),
.A2(n_291),
.B1(n_293),
.B2(n_298),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_332),
.A2(n_340),
.B1(n_337),
.B2(n_336),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_290),
.C(n_292),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_293),
.C(n_298),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_294),
.B(n_319),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_294),
.Y(n_373)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_287),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_325),
.C(n_343),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_365),
.A2(n_340),
.B1(n_339),
.B2(n_322),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_379),
.B1(n_393),
.B2(n_361),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_347),
.Y(n_377)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_346),
.B1(n_342),
.B2(n_330),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_382),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_348),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_390),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_330),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_388),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_275),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_353),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_364),
.A2(n_328),
.B1(n_338),
.B2(n_345),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_389),
.A2(n_373),
.B1(n_363),
.B2(n_357),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_338),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_333),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_359),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_365),
.A2(n_344),
.B1(n_305),
.B2(n_319),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_305),
.C(n_296),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_366),
.C(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_398),
.C(n_403),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_355),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_404),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_371),
.C(n_355),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_357),
.B1(n_354),
.B2(n_367),
.Y(n_405)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_383),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_408),
.C(n_384),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_364),
.C(n_372),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_397),
.B(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_418),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_421),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_399),
.A2(n_380),
.B(n_388),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_416),
.A2(n_408),
.B(n_373),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_410),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_383),
.C(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_422),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_400),
.C(n_396),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_416),
.B(n_400),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_423),
.B(n_425),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_391),
.B1(n_378),
.B2(n_370),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_424),
.A2(n_385),
.B1(n_393),
.B2(n_419),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_420),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_427),
.B(n_429),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_389),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_385),
.B1(n_415),
.B2(n_421),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_407),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_411),
.C(n_422),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_433),
.B(n_437),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_396),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_435),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_440),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_433),
.A2(n_411),
.B(n_426),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_441),
.A2(n_434),
.B(n_436),
.C(n_398),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_438),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_439),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_442),
.B(n_309),
.Y(n_446)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_446),
.Y(n_447)
);


endmodule