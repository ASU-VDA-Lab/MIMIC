module fake_jpeg_13772_n_46 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_32;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_22),
.B(n_23),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_22),
.B(n_24),
.Y(n_35)
);

XNOR2x1_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_31),
.B(n_1),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

MAJx2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_0),
.C(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_40),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_41),
.B(n_37),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_2),
.C(n_3),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_4),
.C(n_5),
.Y(n_46)
);


endmodule