module fake_jpeg_3959_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_29),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_25),
.B1(n_16),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_29),
.B1(n_36),
.B2(n_33),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_32),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_44),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_35),
.B1(n_20),
.B2(n_31),
.Y(n_61)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_63),
.B1(n_30),
.B2(n_20),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_35),
.B1(n_20),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_44),
.B1(n_49),
.B2(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_76),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_41),
.B1(n_46),
.B2(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_77),
.B1(n_68),
.B2(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_54),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_59),
.C(n_69),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.C(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_100),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_67),
.C(n_57),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_78),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_62),
.B1(n_60),
.B2(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_86),
.B1(n_84),
.B2(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_105),
.B1(n_83),
.B2(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_101),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_56),
.B1(n_68),
.B2(n_58),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_114),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_112),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_74),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_97),
.B(n_30),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_73),
.B1(n_84),
.B2(n_58),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_58),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_65),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_73),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_90),
.A3(n_92),
.B1(n_97),
.B2(n_96),
.C1(n_93),
.C2(n_95),
.Y(n_126)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_81),
.B(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_93),
.B(n_106),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_129),
.B(n_131),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_121),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_134),
.B1(n_22),
.B2(n_26),
.Y(n_144)
);

AOI21x1_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_30),
.B(n_20),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_22),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_141),
.C(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_114),
.B1(n_111),
.B2(n_107),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_134),
.B1(n_129),
.B2(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_108),
.C(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_145),
.B(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_117),
.B1(n_122),
.B2(n_19),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_144),
.B1(n_22),
.B2(n_14),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_123),
.B(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_151),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_2),
.CI(n_3),
.CON(n_159),
.SN(n_159)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_141),
.B1(n_140),
.B2(n_136),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_132),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_14),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_3),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_14),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_156),
.CI(n_158),
.CON(n_166),
.SN(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_154),
.C(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_12),
.Y(n_161)
);

AOI31xp67_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_12),
.A3(n_4),
.B(n_5),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_150),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_166),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_167),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_152),
.C(n_4),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_159),
.B1(n_166),
.B2(n_6),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_7),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_3),
.B(n_5),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_7),
.B(n_8),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_164),
.B1(n_9),
.B2(n_11),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_172),
.C(n_169),
.Y(n_177)
);

AOI31xp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_7),
.A3(n_9),
.B(n_11),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.C(n_9),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_11),
.Y(n_180)
);


endmodule