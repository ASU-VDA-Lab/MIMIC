module fake_jpeg_30430_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_2),
.Y(n_67)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_20),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_40),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_47),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_16),
.B1(n_21),
.B2(n_15),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_58),
.B1(n_59),
.B2(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_27),
.B1(n_30),
.B2(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_50),
.B1(n_57),
.B2(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_75),
.Y(n_108)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_63),
.B1(n_64),
.B2(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_87),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_42),
.CI(n_57),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_39),
.C(n_22),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_93),
.C(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_82),
.B1(n_73),
.B2(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_110),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_112),
.B1(n_84),
.B2(n_42),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_13),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_88),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_109),
.C(n_105),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_98),
.B1(n_95),
.B2(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_122),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_110),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_85),
.B(n_89),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_108),
.B(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_74),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_126),
.B(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_76),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_102),
.C(n_101),
.D(n_9),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_136),
.B1(n_95),
.B2(n_119),
.C(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_115),
.B1(n_121),
.B2(n_104),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_114),
.C(n_116),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_135),
.C(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_116),
.B1(n_126),
.B2(n_113),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_149),
.B(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_150),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_134),
.C(n_129),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_R g159 ( 
.A(n_152),
.B(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_141),
.B(n_147),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_152),
.B(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_156),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_100),
.B(n_75),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_120),
.B1(n_156),
.B2(n_108),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_167),
.B(n_80),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_3),
.B(n_7),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.C(n_7),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_11),
.B(n_13),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_3),
.Y(n_175)
);


endmodule