module fake_netlist_5_1033_n_2226 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2226);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2226;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2193;
wire n_2052;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2111;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_75),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_39),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_23),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_164),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_107),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_163),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_84),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_204),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_77),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_37),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_145),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_23),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_188),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_50),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_71),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_152),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_35),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_190),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_66),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_192),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_64),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_133),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_19),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_161),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_225),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_138),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_63),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_154),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_203),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_92),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_52),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_185),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_72),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_169),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_149),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_28),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_122),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_69),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_112),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_165),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_230),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_123),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_98),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_216),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_38),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_47),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_0),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_132),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_182),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_79),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_175),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_39),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_97),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_19),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_113),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_134),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_3),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_32),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_136),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_61),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_110),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_196),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_77),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_45),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_153),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_197),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_181),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_99),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_27),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_24),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_174),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_80),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_70),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_96),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_115),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_8),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_78),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_49),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_69),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_90),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_63),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_119),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_137),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_116),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_0),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_44),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_212),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_12),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_127),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_45),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_125),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_34),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_109),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_189),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_193),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_210),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_150),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_186),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_5),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_2),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_13),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_15),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_48),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_67),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_217),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_24),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_100),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_223),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_130),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_170),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_31),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_214),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_44),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_162),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_57),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_207),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_61),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_168),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_105),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_46),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_215),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_2),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_148),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_87),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_21),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_36),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_28),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_144),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_108),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_179),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_9),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_33),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_59),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_76),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_213),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_200),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_74),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_219),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_41),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_81),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_201),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_57),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_151),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_139),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_34),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_53),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_158),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_155),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_120),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_114),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_6),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_50),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_208),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_12),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_54),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_177),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_166),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_17),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_20),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_56),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_48),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_167),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_118),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_4),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_173),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_103),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_56),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_1),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_29),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_221),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_15),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_30),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_104),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_121),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_205),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_94),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_209),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_40),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_72),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_124),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_178),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_229),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_234),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_82),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_106),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_67),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_128),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_85),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_75),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_59),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_143),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_62),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_117),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_88),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_461),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_294),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_316),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_301),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_248),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_339),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_301),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_301),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_301),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_351),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_358),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_331),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_301),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_349),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_301),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_352),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_301),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_237),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_301),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_241),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_260),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_260),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_330),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_260),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_279),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_260),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_236),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_260),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_264),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_278),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_424),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_259),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_280),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_241),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_365),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_283),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_283),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_267),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_381),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_442),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_286),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_453),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_281),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_281),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_292),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_413),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_295),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_314),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_288),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_288),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_237),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_406),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_406),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_319),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_418),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_321),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_274),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_325),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_277),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_299),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_238),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_251),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_256),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_261),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_326),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_289),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_264),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_298),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_328),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_268),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_282),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_250),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_303),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_313),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_323),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_356),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_332),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_359),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_361),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_271),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_400),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_363),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_333),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_371),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_375),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_304),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_271),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_300),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_387),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_306),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_342),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_299),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_348),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_348),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_240),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_398),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_357),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_240),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_398),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_409),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_423),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_309),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_315),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_414),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_370),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_373),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_439),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_374),
.Y(n_584)
);

INVxp33_ASAP7_75t_SL g585 ( 
.A(n_258),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_440),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_376),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_423),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_378),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_450),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_451),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_383),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_300),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_311),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_385),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_235),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_389),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_317),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_487),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_338),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_530),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_476),
.B(n_311),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_495),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_496),
.B(n_369),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_502),
.A2(n_265),
.B1(n_269),
.B2(n_258),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_496),
.B(n_540),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_532),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_468),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_477),
.B(n_369),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_287),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_469),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_492),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_540),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_492),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_491),
.A2(n_394),
.B1(n_403),
.B2(n_392),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_553),
.B(n_434),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_494),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_472),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

CKINVDCx6p67_ASAP7_75t_R g629 ( 
.A(n_516),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_553),
.B(n_434),
.Y(n_632)
);

NOR2x1_ASAP7_75t_L g633 ( 
.A(n_539),
.B(n_244),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_500),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_472),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_501),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_508),
.A2(n_554),
.B1(n_471),
.B2(n_489),
.Y(n_638)
);

XNOR2x1_ASAP7_75t_L g639 ( 
.A(n_545),
.B(n_265),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_493),
.B(n_287),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_475),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_541),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_475),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_593),
.B(n_338),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_562),
.B(n_337),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_562),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_594),
.B(n_337),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_535),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_473),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_474),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_482),
.A2(n_417),
.B1(n_426),
.B2(n_404),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_536),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_467),
.B(n_420),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_484),
.A2(n_430),
.B1(n_431),
.B2(n_269),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_480),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_479),
.Y(n_658)
);

INVxp33_ASAP7_75t_SL g659 ( 
.A(n_493),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_572),
.A2(n_432),
.B1(n_433),
.B2(n_431),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_537),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_486),
.B(n_420),
.Y(n_662)
);

BUFx8_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_498),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_481),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_498),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_483),
.Y(n_669)
);

OA21x2_ASAP7_75t_L g670 ( 
.A1(n_485),
.A2(n_290),
.B(n_270),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_556),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_503),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_556),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_590),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_560),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_503),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_590),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_506),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_513),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_564),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_507),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_514),
.B(n_270),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_507),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_533),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_519),
.B(n_290),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_585),
.A2(n_432),
.B1(n_433),
.B2(n_464),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_533),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_504),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_566),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_576),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_291),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_511),
.B(n_320),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_619),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_655),
.B(n_578),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_671),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_641),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_671),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_612),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_641),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_607),
.B(n_598),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_602),
.B(n_583),
.C(n_574),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_673),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_602),
.B(n_521),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_673),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_619),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_651),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_605),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_615),
.B(n_511),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_671),
.Y(n_714)
);

NOR2x1p5_ASAP7_75t_L g715 ( 
.A(n_676),
.B(n_436),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_651),
.Y(n_716)
);

CKINVDCx6p67_ASAP7_75t_R g717 ( 
.A(n_629),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_669),
.Y(n_718)
);

CKINVDCx11_ASAP7_75t_R g719 ( 
.A(n_614),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_640),
.B(n_515),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_669),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_605),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_647),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_648),
.B(n_515),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_648),
.B(n_517),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_647),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_608),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_608),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_611),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_611),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_618),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_618),
.Y(n_732)
);

XNOR2xp5_ASAP7_75t_L g733 ( 
.A(n_639),
.B(n_478),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_649),
.A2(n_372),
.B1(n_296),
.B2(n_307),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_644),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_612),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_517),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_691),
.B(n_518),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_691),
.B(n_518),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_671),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_647),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_644),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_652),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_609),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_599),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_676),
.B(n_526),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_671),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_633),
.B(n_372),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_683),
.B(n_548),
.C(n_547),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_652),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_658),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_686),
.B(n_551),
.C(n_549),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_652),
.B(n_526),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_696),
.B(n_555),
.C(n_552),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_634),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_697),
.B(n_528),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_666),
.B(n_528),
.Y(n_759)
);

XOR2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_505),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_658),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_600),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_666),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_676),
.B(n_531),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_666),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_601),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_649),
.A2(n_296),
.B1(n_307),
.B2(n_291),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_601),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_606),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_636),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_658),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_620),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_658),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_603),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_657),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_620),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_621),
.B(n_531),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_616),
.B(n_538),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_659),
.B(n_538),
.Y(n_780)
);

INVxp33_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_609),
.B(n_542),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_658),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_659),
.B(n_542),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_609),
.Y(n_785)
);

AND3x1_ASAP7_75t_L g786 ( 
.A(n_660),
.B(n_569),
.C(n_524),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_622),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_637),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_623),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_634),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_623),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_622),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_622),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_632),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_624),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_645),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_653),
.B(n_550),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_624),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_638),
.B(n_550),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_646),
.B(n_625),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_663),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_625),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_664),
.B(n_557),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_664),
.B(n_557),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_627),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_627),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_628),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_628),
.B(n_565),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_670),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_630),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_630),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_631),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_631),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_656),
.A2(n_687),
.B1(n_397),
.B2(n_312),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_674),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_678),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_678),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_663),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_649),
.B(n_645),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_678),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_SL g824 ( 
.A(n_688),
.B(n_565),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_678),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_603),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_571),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_670),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_678),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_684),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_670),
.Y(n_831)
);

INVx8_ASAP7_75t_L g832 ( 
.A(n_684),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_674),
.Y(n_833)
);

BUFx4f_ASAP7_75t_L g834 ( 
.A(n_670),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_684),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_684),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_677),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_684),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_685),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_685),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_662),
.A2(n_308),
.B(n_273),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_680),
.B(n_522),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_685),
.B(n_571),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_685),
.B(n_580),
.Y(n_844)
);

BUFx10_ASAP7_75t_L g845 ( 
.A(n_626),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_685),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_692),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_617),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_692),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_677),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_692),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_692),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_692),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_693),
.B(n_580),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_L g855 ( 
.A(n_642),
.B(n_252),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_693),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_693),
.B(n_582),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_693),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_672),
.B(n_582),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_680),
.B(n_584),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_693),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_613),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_818),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_834),
.B(n_252),
.Y(n_864)
);

OAI221xp5_ASAP7_75t_L g865 ( 
.A1(n_734),
.A2(n_610),
.B1(n_654),
.B2(n_689),
.C(n_650),
.Y(n_865)
);

BUFx12f_ASAP7_75t_SL g866 ( 
.A(n_749),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_796),
.B(n_635),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_SL g868 ( 
.A(n_803),
.B(n_613),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_818),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_745),
.B(n_396),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_794),
.B(n_587),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_801),
.B(n_587),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_745),
.B(n_589),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_779),
.B(n_589),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_833),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_834),
.B(n_252),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_719),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_833),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_785),
.B(n_592),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_796),
.B(n_635),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_756),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_756),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_758),
.B(n_713),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_762),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_803),
.B(n_821),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_762),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_785),
.B(n_592),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_776),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_787),
.B(n_595),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_706),
.B(n_597),
.C(n_595),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_766),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_837),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_698),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_776),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_766),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_736),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_775),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_787),
.B(n_597),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_792),
.B(n_661),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_800),
.A2(n_308),
.B1(n_275),
.B2(n_284),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_850),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_769),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_792),
.A2(n_510),
.B1(n_512),
.B2(n_509),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_782),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_706),
.B(n_663),
.C(n_665),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_842),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_703),
.B(n_667),
.Y(n_907)
);

BUFx6f_ASAP7_75t_SL g908 ( 
.A(n_862),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_703),
.B(n_768),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_827),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_754),
.B(n_396),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_700),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_775),
.B(n_643),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_811),
.B(n_285),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_842),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_793),
.B(n_239),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_736),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_793),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_698),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_821),
.B(n_525),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_822),
.A2(n_335),
.B1(n_297),
.B2(n_302),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_780),
.B(n_643),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_768),
.B(n_254),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_812),
.A2(n_276),
.B1(n_293),
.B2(n_266),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_305),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_789),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_770),
.B(n_310),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_759),
.B(n_239),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_834),
.B(n_252),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_737),
.B(n_242),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_773),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_773),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_708),
.B(n_675),
.Y(n_934)
);

NAND2x1_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_252),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_789),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_860),
.B(n_529),
.C(n_527),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_699),
.A2(n_334),
.B1(n_318),
.B2(n_322),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_708),
.A2(n_559),
.B(n_558),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_724),
.B(n_242),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_793),
.B(n_243),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_771),
.B(n_329),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_771),
.B(n_336),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_784),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_777),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_L g946 ( 
.A(n_843),
.B(n_396),
.Y(n_946)
);

XOR2xp5_ASAP7_75t_L g947 ( 
.A(n_760),
.B(n_617),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_723),
.A2(n_448),
.B(n_344),
.C(n_353),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_777),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_710),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_760),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_725),
.B(n_243),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_705),
.B(n_675),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_738),
.B(n_245),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_710),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_720),
.B(n_245),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_SL g957 ( 
.A1(n_749),
.A2(n_694),
.B1(n_681),
.B2(n_458),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_810),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_810),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_788),
.B(n_343),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_788),
.B(n_355),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_813),
.B(n_364),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_761),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_749),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_739),
.B(n_845),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_824),
.B(n_798),
.C(n_778),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_844),
.B(n_246),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_813),
.B(n_812),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_812),
.B(n_384),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_828),
.B(n_386),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_L g971 ( 
.A(n_854),
.B(n_396),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_857),
.B(n_246),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_712),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_767),
.A2(n_390),
.B1(n_391),
.B2(n_395),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_828),
.B(n_422),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_845),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_749),
.B(n_247),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_826),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_SL g979 ( 
.A(n_828),
.B(n_255),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_817),
.B(n_247),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_786),
.A2(n_408),
.B1(n_324),
.B2(n_327),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_723),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_726),
.B(n_255),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_726),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_761),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_786),
.B(n_255),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_805),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_807),
.B(n_694),
.C(n_681),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_845),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_859),
.B(n_577),
.C(n_563),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_733),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_831),
.B(n_425),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_715),
.B(n_629),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_741),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_741),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_747),
.B(n_581),
.C(n_579),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_764),
.B(n_249),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_743),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_831),
.B(n_249),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_743),
.B(n_255),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_791),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_715),
.B(n_586),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_791),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_751),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_862),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_831),
.B(n_428),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_751),
.B(n_255),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_848),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_795),
.Y(n_1009)
);

OAI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_781),
.A2(n_463),
.B1(n_455),
.B2(n_456),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_763),
.B(n_437),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_795),
.B(n_253),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_763),
.B(n_262),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_765),
.A2(n_416),
.B1(n_340),
.B2(n_341),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_799),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_799),
.B(n_253),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_804),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_765),
.B(n_804),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_862),
.B(n_591),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_808),
.B(n_460),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_808),
.B(n_690),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_809),
.B(n_690),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_809),
.B(n_679),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_814),
.B(n_679),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_814),
.B(n_682),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_700),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_815),
.B(n_816),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_816),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_712),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_750),
.B(n_257),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_826),
.B(n_695),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_722),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_883),
.A2(n_716),
.B1(n_718),
.B2(n_711),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_918),
.B(n_772),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_914),
.B(n_716),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1029),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1031),
.B(n_733),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_893),
.B(n_750),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_888),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_881),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_894),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_918),
.B(n_772),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_914),
.B(n_718),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_972),
.B(n_721),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_972),
.B(n_929),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_929),
.B(n_721),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_918),
.B(n_761),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1029),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1032),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_900),
.A2(n_345),
.B1(n_399),
.B2(n_701),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_874),
.B(n_748),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_944),
.B(n_755),
.C(n_753),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_874),
.B(n_863),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1032),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_SL g1055 ( 
.A1(n_957),
.A2(n_436),
.B1(n_441),
.B2(n_443),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_917),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_934),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_893),
.B(n_753),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1008),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_1019),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_882),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_910),
.B(n_755),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_919),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_882),
.Y(n_1064)
);

INVxp33_ASAP7_75t_L g1065 ( 
.A(n_913),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_963),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_884),
.Y(n_1068)
);

NAND2xp33_ASAP7_75t_SL g1069 ( 
.A(n_918),
.B(n_262),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_966),
.A2(n_861),
.B1(n_858),
.B2(n_851),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_869),
.B(n_748),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_875),
.B(n_748),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_884),
.Y(n_1073)
);

AND2x6_ASAP7_75t_L g1074 ( 
.A(n_968),
.B(n_819),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_917),
.B(n_761),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_917),
.B(n_761),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_872),
.B(n_740),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_904),
.A2(n_861),
.B1(n_858),
.B2(n_851),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_885),
.B(n_717),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_886),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_878),
.B(n_701),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_917),
.B(n_783),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_886),
.Y(n_1083)
);

AND2x6_ASAP7_75t_SL g1084 ( 
.A(n_980),
.B(n_567),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_891),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_987),
.B(n_740),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_891),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_892),
.B(n_704),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_895),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_901),
.B(n_707),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1002),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_979),
.A2(n_853),
.B(n_820),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_919),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_902),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_927),
.B(n_936),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_902),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_896),
.B(n_871),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_913),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_871),
.B(n_717),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_958),
.B(n_709),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_867),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_924),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_959),
.B(n_709),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_909),
.B(n_783),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_897),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_940),
.B(n_830),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_900),
.A2(n_396),
.B1(n_435),
.B2(n_731),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_924),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_940),
.B(n_830),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_932),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_952),
.B(n_830),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_978),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_932),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_877),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_906),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_933),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_952),
.B(n_835),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_950),
.B(n_695),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_915),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_933),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_931),
.B(n_835),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_931),
.B(n_835),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_945),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_880),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_945),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_955),
.B(n_819),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1005),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_964),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_980),
.B(n_890),
.Y(n_1129)
);

NAND2x1p5_ASAP7_75t_L g1130 ( 
.A(n_963),
.B(n_985),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_949),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1005),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_949),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_866),
.B(n_841),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_903),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_965),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1001),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1003),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_963),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_963),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_999),
.B(n_838),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_885),
.B(n_832),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_982),
.B(n_838),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_997),
.A2(n_853),
.B1(n_836),
.B2(n_820),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1009),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_984),
.B(n_838),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_864),
.A2(n_832),
.B(n_876),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_996),
.B(n_825),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_953),
.B(n_568),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_985),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_925),
.B(n_954),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_981),
.A2(n_443),
.B1(n_462),
.B2(n_444),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_985),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_985),
.B(n_772),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1015),
.Y(n_1155)
);

OR2x6_ASAP7_75t_SL g1156 ( 
.A(n_905),
.B(n_441),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_920),
.B(n_832),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_973),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_921),
.A2(n_731),
.B(n_732),
.C(n_855),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_976),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_997),
.A2(n_839),
.B1(n_825),
.B2(n_849),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_908),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1017),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_994),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_986),
.B(n_774),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_995),
.B(n_840),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_998),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1004),
.B(n_840),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_976),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_989),
.B(n_829),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_925),
.B(n_568),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_900),
.A2(n_435),
.B1(n_396),
.B2(n_732),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1028),
.B(n_840),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_907),
.B(n_846),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1027),
.Y(n_1175)
);

OR2x2_ASAP7_75t_SL g1176 ( 
.A(n_873),
.B(n_262),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_947),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_954),
.A2(n_444),
.B(n_462),
.C(n_464),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1018),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1021),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1022),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_991),
.B(n_570),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_935),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_899),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_864),
.A2(n_832),
.B(n_774),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1023),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_986),
.B(n_783),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1024),
.B(n_846),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1025),
.B(n_846),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_879),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_887),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_969),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_962),
.B(n_757),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1011),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_923),
.B(n_757),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_970),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_926),
.B(n_757),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_920),
.B(n_832),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_876),
.A2(n_774),
.B(n_702),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_993),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_920),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_928),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_942),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_943),
.B(n_797),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_975),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1010),
.B(n_263),
.C(n_257),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_960),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_922),
.B(n_570),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_992),
.Y(n_1209)
);

NOR2x2_ASAP7_75t_L g1210 ( 
.A(n_868),
.B(n_829),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_961),
.B(n_1006),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_898),
.B(n_700),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_977),
.B(n_700),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1147),
.A2(n_930),
.B(n_912),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_930),
.B(n_1026),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1045),
.B(n_951),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_SL g1218 ( 
.A(n_1152),
.B(n_1178),
.C(n_1129),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1151),
.A2(n_977),
.B1(n_1030),
.B2(n_865),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1067),
.A2(n_870),
.B(n_856),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1092),
.A2(n_839),
.B(n_836),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1129),
.A2(n_1178),
.B(n_1152),
.C(n_1053),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1108),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1149),
.B(n_990),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_967),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1202),
.B(n_938),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1186),
.B(n_939),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1062),
.A2(n_911),
.B(n_889),
.C(n_956),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1062),
.B(n_916),
.Y(n_1229)
);

BUFx4f_ASAP7_75t_L g1230 ( 
.A(n_1079),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1199),
.A2(n_849),
.B(n_847),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1203),
.A2(n_941),
.B(n_971),
.C(n_946),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1067),
.A2(n_856),
.B(n_852),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_SL g1234 ( 
.A(n_1067),
.B(n_983),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1105),
.B(n_908),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_1112),
.B(n_841),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1115),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1060),
.B(n_988),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1207),
.A2(n_1014),
.B(n_1016),
.C(n_1012),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1052),
.A2(n_1171),
.B1(n_1058),
.B2(n_1038),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1177),
.B(n_937),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1059),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_R g1243 ( 
.A(n_1098),
.B(n_263),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1056),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1108),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1115),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1119),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1099),
.B(n_320),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1190),
.B(n_783),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1119),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_SL g1251 ( 
.A(n_1165),
.B(n_320),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1035),
.B(n_974),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1056),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1186),
.B(n_847),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_SL g1255 ( 
.A(n_1050),
.B(n_346),
.C(n_272),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1056),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1067),
.A2(n_1209),
.B(n_1185),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1043),
.B(n_735),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1040),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1209),
.A2(n_856),
.B(n_852),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1191),
.B(n_783),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1039),
.B(n_272),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1056),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1116),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1116),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1187),
.A2(n_948),
.B(n_1013),
.C(n_1000),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1097),
.A2(n_1007),
.B(n_1000),
.C(n_855),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1141),
.A2(n_852),
.B(n_702),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1192),
.A2(n_702),
.B(n_700),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1194),
.A2(n_802),
.B(n_797),
.C(n_742),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1169),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1131),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1041),
.B(n_346),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1169),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1091),
.A2(n_377),
.B1(n_380),
.B2(n_382),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1175),
.B(n_744),
.Y(n_1276)
);

O2A1O1Ixp5_ASAP7_75t_L g1277 ( 
.A1(n_1077),
.A2(n_802),
.B(n_797),
.C(n_790),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1139),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1121),
.A2(n_702),
.B(n_714),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1122),
.A2(n_714),
.B(n_790),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1050),
.A2(n_447),
.B1(n_347),
.B2(n_438),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1131),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1139),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1142),
.B(n_790),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_714),
.B(n_752),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1063),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1140),
.B(n_714),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1182),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1061),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1046),
.A2(n_722),
.B(n_727),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1163),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1163),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1063),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1064),
.Y(n_1294)
);

NOR3xp33_ASAP7_75t_L g1295 ( 
.A(n_1037),
.B(n_438),
.C(n_465),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1057),
.B(n_573),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1139),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1184),
.B(n_728),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1055),
.A2(n_454),
.B1(n_447),
.B2(n_449),
.C(n_465),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1109),
.A2(n_1117),
.B(n_1111),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1139),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1140),
.B(n_823),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1093),
.Y(n_1303)
);

CKINVDCx10_ASAP7_75t_R g1304 ( 
.A(n_1079),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1080),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1135),
.B(n_573),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1184),
.B(n_1180),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1093),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1038),
.A2(n_368),
.B1(n_354),
.B2(n_360),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1051),
.A2(n_752),
.B(n_823),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1101),
.A2(n_746),
.B(n_729),
.C(n_730),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1184),
.B(n_347),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1154),
.A2(n_1193),
.B(n_1195),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1180),
.B(n_730),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1181),
.B(n_445),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1047),
.A2(n_588),
.B(n_575),
.C(n_396),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1101),
.A2(n_1095),
.B(n_1044),
.C(n_1136),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1127),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1127),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1154),
.A2(n_1072),
.B(n_1071),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1165),
.A2(n_445),
.B1(n_449),
.B2(n_452),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1058),
.B(n_452),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1107),
.A2(n_457),
.B1(n_459),
.B2(n_454),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1098),
.A2(n_457),
.B1(n_459),
.B2(n_362),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1181),
.B(n_366),
.Y(n_1325)
);

OAI22x1_ASAP7_75t_L g1326 ( 
.A1(n_1201),
.A2(n_367),
.B1(n_466),
.B2(n_388),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1150),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1068),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1107),
.A2(n_588),
.B1(n_575),
.B2(n_419),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1065),
.B(n_393),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1172),
.A2(n_1164),
.B1(n_1167),
.B2(n_1213),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1083),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1150),
.Y(n_1333)
);

O2A1O1Ixp5_ASAP7_75t_SL g1334 ( 
.A1(n_1104),
.A2(n_379),
.B(n_446),
.C(n_435),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1132),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1065),
.B(n_401),
.Y(n_1336)
);

AOI221xp5_ASAP7_75t_L g1337 ( 
.A1(n_1206),
.A2(n_412),
.B1(n_429),
.B2(n_421),
.C(n_402),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1153),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1196),
.A2(n_415),
.B(n_407),
.C(n_410),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1086),
.B(n_262),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1124),
.B(n_379),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1086),
.B(n_379),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1200),
.B(n_83),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1114),
.B(n_86),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1196),
.B(n_262),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1068),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1205),
.B(n_350),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_446),
.B1(n_435),
.B2(n_419),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1197),
.A2(n_752),
.B(n_823),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1160),
.B(n_446),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1104),
.A2(n_752),
.B(n_823),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1204),
.A2(n_752),
.B(n_823),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1128),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1085),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1087),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1205),
.A2(n_419),
.B(n_350),
.C(n_435),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1075),
.A2(n_752),
.B(n_823),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1118),
.B(n_350),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1212),
.A2(n_806),
.B(n_350),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1212),
.A2(n_419),
.B(n_350),
.C(n_435),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1066),
.B(n_419),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1188),
.A2(n_1189),
.B(n_1042),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1066),
.A2(n_435),
.B1(n_3),
.B2(n_4),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1033),
.A2(n_1),
.B(n_5),
.C(n_7),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1156),
.Y(n_1365)
);

NOR2x1_ASAP7_75t_SL g1366 ( 
.A(n_1153),
.B(n_806),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1118),
.B(n_7),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1132),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1084),
.B(n_10),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1034),
.A2(n_806),
.B(n_233),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_13),
.B2(n_14),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1331),
.A2(n_1042),
.B(n_1034),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1240),
.B(n_1214),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1368),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1360),
.A2(n_1174),
.A3(n_1073),
.B(n_1113),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1231),
.A2(n_1221),
.B(n_1320),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1300),
.A2(n_1144),
.B(n_1161),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1216),
.A2(n_1158),
.B(n_1076),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_R g1380 ( 
.A(n_1243),
.B(n_1218),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1229),
.A2(n_1206),
.B(n_1159),
.C(n_1078),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1328),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1357),
.A2(n_1173),
.B(n_1143),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1259),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1217),
.B(n_1288),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1288),
.B(n_1200),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1241),
.B(n_1208),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1368),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1215),
.A2(n_1214),
.B(n_1076),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1270),
.A2(n_1073),
.A3(n_1138),
.B(n_1145),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1356),
.A2(n_1138),
.A3(n_1145),
.B(n_1120),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1318),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_SL g1393 ( 
.A1(n_1228),
.A2(n_1082),
.B(n_1166),
.C(n_1146),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1335),
.B(n_1142),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1368),
.Y(n_1395)
);

AND2x6_ASAP7_75t_SL g1396 ( 
.A(n_1369),
.B(n_1142),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1242),
.B(n_1208),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1351),
.A2(n_1168),
.B(n_1082),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1344),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1331),
.A2(n_1214),
.B(n_1130),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_SL g1401 ( 
.A(n_1327),
.B(n_1162),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1327),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1340),
.A2(n_1120),
.A3(n_1102),
.B(n_1123),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1307),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1219),
.A2(n_1176),
.B1(n_1157),
.B2(n_1198),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1289),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1255),
.A2(n_1148),
.B(n_1210),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1319),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1364),
.A2(n_1100),
.B(n_1081),
.C(n_1088),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1257),
.A2(n_1070),
.B(n_1094),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1279),
.A2(n_1133),
.B(n_1096),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1362),
.A2(n_1158),
.B(n_1214),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1313),
.A2(n_1074),
.B(n_1103),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1252),
.B(n_1090),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_R g1415 ( 
.A(n_1236),
.B(n_1134),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1268),
.A2(n_1137),
.B(n_1089),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1303),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1157),
.C(n_1148),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1304),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_SL g1420 ( 
.A(n_1251),
.B(n_1134),
.C(n_1069),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1371),
.A2(n_1157),
.B1(n_1198),
.B2(n_1158),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1317),
.A2(n_1170),
.B(n_1069),
.C(n_1126),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1308),
.B(n_1126),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1280),
.A2(n_1125),
.B(n_1110),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1327),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1285),
.A2(n_1155),
.B(n_1130),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1371),
.A2(n_1054),
.B(n_1036),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1226),
.B(n_1048),
.Y(n_1428)
);

NOR4xp25_ASAP7_75t_L g1429 ( 
.A(n_1281),
.B(n_1049),
.C(n_1210),
.D(n_1183),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1294),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_SL g1431 ( 
.A(n_1327),
.B(n_1158),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1239),
.A2(n_1074),
.B(n_806),
.C(n_16),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1305),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1346),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1332),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1269),
.A2(n_1074),
.B(n_228),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1224),
.A2(n_1367),
.B(n_1347),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1263),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1308),
.B(n_1074),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1232),
.A2(n_227),
.B(n_224),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1354),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1355),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1341),
.A2(n_11),
.B(n_14),
.C(n_17),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1234),
.A2(n_195),
.B(n_194),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1310),
.A2(n_187),
.B(n_183),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1334),
.A2(n_176),
.B(n_172),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1306),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1227),
.B(n_11),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1281),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_1449)
);

AOI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1359),
.A2(n_160),
.B(n_147),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1248),
.B(n_18),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1345),
.A2(n_146),
.B(n_142),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1290),
.A2(n_140),
.B(n_131),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1295),
.A2(n_1238),
.B1(n_1330),
.B2(n_1336),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1290),
.A2(n_129),
.B(n_126),
.Y(n_1455)
);

AO31x2_ASAP7_75t_L g1456 ( 
.A1(n_1329),
.A2(n_22),
.A3(n_25),
.B(n_26),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1248),
.B(n_25),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1329),
.A2(n_27),
.A3(n_29),
.B(n_30),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_SL g1459 ( 
.A(n_1353),
.B(n_31),
.Y(n_1459)
);

AO21x1_ASAP7_75t_L g1460 ( 
.A1(n_1342),
.A2(n_32),
.B(n_36),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1303),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1237),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1246),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_SL g1464 ( 
.A1(n_1312),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1220),
.A2(n_1260),
.B(n_1258),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1247),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1278),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1235),
.B(n_42),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1225),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1250),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1299),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1363),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1223),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1296),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1235),
.B(n_55),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1349),
.A2(n_58),
.A3(n_60),
.B(n_62),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1266),
.A2(n_58),
.B(n_64),
.C(n_65),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1350),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1352),
.A2(n_101),
.B(n_95),
.Y(n_1479)
);

AOI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1249),
.A2(n_91),
.B(n_89),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1277),
.A2(n_68),
.B(n_70),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1254),
.B(n_76),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1298),
.A2(n_71),
.B(n_73),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1262),
.B(n_73),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1273),
.B(n_1293),
.Y(n_1485)
);

NAND2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1333),
.B(n_1338),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1267),
.A2(n_1254),
.B(n_1314),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1245),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1263),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1324),
.B(n_1286),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1284),
.A2(n_1343),
.B(n_1370),
.Y(n_1491)
);

NOR2x1_ASAP7_75t_L g1492 ( 
.A(n_1338),
.B(n_1256),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1358),
.A2(n_1276),
.B(n_1339),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1264),
.Y(n_1494)
);

O2A1O1Ixp5_ASAP7_75t_L g1495 ( 
.A1(n_1261),
.A2(n_1321),
.B(n_1315),
.C(n_1323),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1348),
.A2(n_1337),
.B(n_1361),
.C(n_1315),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1233),
.A2(n_1311),
.B(n_1287),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1325),
.A2(n_1292),
.B(n_1291),
.Y(n_1498)
);

CKINVDCx6p67_ASAP7_75t_R g1499 ( 
.A(n_1326),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1265),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1343),
.B(n_1365),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1309),
.B(n_1321),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1302),
.A2(n_1244),
.B(n_1256),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1230),
.B(n_1323),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1253),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1272),
.A2(n_1282),
.B(n_1283),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_1253),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1283),
.B(n_1253),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1284),
.B(n_1278),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1278),
.B(n_1297),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1275),
.A2(n_1230),
.B(n_1297),
.C(n_1301),
.Y(n_1511)
);

CKINVDCx6p67_ASAP7_75t_R g1512 ( 
.A(n_1297),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1366),
.A2(n_1316),
.B(n_1301),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1301),
.A2(n_1045),
.B(n_1331),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1216),
.A2(n_1211),
.B(n_1300),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1259),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1328),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_SL g1518 ( 
.A1(n_1340),
.A2(n_1151),
.B(n_1045),
.Y(n_1518)
);

BUFx4f_ASAP7_75t_SL g1519 ( 
.A(n_1271),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1229),
.B(n_1217),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1242),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1240),
.B(n_1045),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1240),
.A2(n_1045),
.B1(n_1151),
.B2(n_1219),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1240),
.A2(n_1045),
.B1(n_1151),
.B2(n_1219),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1231),
.A2(n_1221),
.B(n_1320),
.Y(n_1525)
);

AO31x2_ASAP7_75t_L g1526 ( 
.A1(n_1360),
.A2(n_1300),
.A3(n_1270),
.B(n_1356),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1259),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1216),
.A2(n_1211),
.B(n_1300),
.Y(n_1528)
);

AOI21xp33_ASAP7_75t_L g1529 ( 
.A1(n_1222),
.A2(n_1045),
.B(n_1151),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1231),
.A2(n_1221),
.B(n_1320),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1240),
.B(n_1045),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1240),
.B(n_1045),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1306),
.B(n_1217),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1307),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1229),
.B(n_1217),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_SL g1536 ( 
.A1(n_1228),
.A2(n_1045),
.B(n_1187),
.C(n_883),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1368),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1463),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1521),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1533),
.B(n_1520),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1484),
.B(n_1457),
.C(n_1451),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1461),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1525),
.A2(n_1436),
.B(n_1465),
.Y(n_1543)
);

O2A1O1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1535),
.A2(n_1443),
.B(n_1471),
.C(n_1477),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1447),
.B(n_1485),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1481),
.A2(n_1413),
.B(n_1529),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1439),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1419),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1389),
.A2(n_1411),
.B(n_1416),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1389),
.A2(n_1424),
.B(n_1497),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1447),
.B(n_1474),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1382),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1454),
.A2(n_1496),
.B(n_1523),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1425),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1523),
.A2(n_1524),
.B1(n_1472),
.B2(n_1531),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1439),
.B(n_1509),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1410),
.A2(n_1379),
.B(n_1383),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1426),
.A2(n_1412),
.B(n_1398),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1374),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1372),
.A2(n_1414),
.B(n_1400),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1434),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1406),
.Y(n_1562)
);

INVx4_ASAP7_75t_SL g1563 ( 
.A(n_1456),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1445),
.A2(n_1479),
.B(n_1518),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1404),
.B(n_1534),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1394),
.B(n_1511),
.Y(n_1566)
);

AOI22x1_ASAP7_75t_L g1567 ( 
.A1(n_1455),
.A2(n_1483),
.B1(n_1504),
.B2(n_1446),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1524),
.A2(n_1472),
.B1(n_1532),
.B2(n_1531),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_SL g1569 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1399),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1517),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1418),
.B(n_1394),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1390),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1437),
.A2(n_1450),
.B(n_1506),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1430),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1487),
.A2(n_1513),
.B(n_1452),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1522),
.A2(n_1478),
.B1(n_1460),
.B2(n_1468),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1433),
.Y(n_1578)
);

AND2x2_ASAP7_75t_SL g1579 ( 
.A(n_1429),
.B(n_1373),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1409),
.A2(n_1381),
.B(n_1495),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1376),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1374),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1386),
.B(n_1385),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1405),
.A2(n_1421),
.B(n_1448),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1388),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1435),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_SL g1587 ( 
.A(n_1420),
.B(n_1394),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_R g1588 ( 
.A(n_1373),
.B(n_1493),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_SL g1589 ( 
.A1(n_1469),
.A2(n_1449),
.B(n_1414),
.C(n_1422),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1388),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1387),
.B(n_1501),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1376),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1441),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1536),
.A2(n_1428),
.B(n_1407),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1483),
.A2(n_1448),
.B(n_1482),
.Y(n_1595)
);

CKINVDCx11_ASAP7_75t_R g1596 ( 
.A(n_1396),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1475),
.A2(n_1459),
.B1(n_1499),
.B2(n_1482),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1480),
.A2(n_1498),
.B(n_1503),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1442),
.Y(n_1599)
);

OAI22x1_ASAP7_75t_L g1600 ( 
.A1(n_1466),
.A2(n_1490),
.B1(n_1527),
.B2(n_1516),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1462),
.A2(n_1470),
.B1(n_1453),
.B2(n_1494),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1498),
.A2(n_1493),
.B(n_1440),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1519),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1464),
.A2(n_1427),
.B(n_1393),
.Y(n_1604)
);

BUFx8_ASAP7_75t_L g1605 ( 
.A(n_1537),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1423),
.B(n_1397),
.Y(n_1606)
);

AOI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1415),
.A2(n_1380),
.B(n_1378),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1508),
.A2(n_1492),
.B(n_1510),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1473),
.A2(n_1500),
.B(n_1488),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1510),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1438),
.A2(n_1489),
.B(n_1486),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1505),
.B(n_1417),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1456),
.Y(n_1613)
);

OAI222xp33_ASAP7_75t_L g1614 ( 
.A1(n_1401),
.A2(n_1505),
.B1(n_1486),
.B2(n_1408),
.C1(n_1392),
.C2(n_1423),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1438),
.A2(n_1489),
.B(n_1453),
.C(n_1458),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1391),
.Y(n_1616)
);

AND2x6_ASAP7_75t_L g1617 ( 
.A(n_1467),
.B(n_1395),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1395),
.B(n_1467),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1403),
.A2(n_1375),
.B(n_1526),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1512),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1431),
.A2(n_1526),
.B1(n_1507),
.B2(n_1375),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1375),
.A2(n_1526),
.B(n_1403),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1476),
.A2(n_1458),
.B(n_1507),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1476),
.A2(n_1525),
.B(n_1377),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1476),
.A2(n_1151),
.B1(n_1229),
.B2(n_1255),
.Y(n_1625)
);

OAI222xp33_ASAP7_75t_L g1626 ( 
.A1(n_1472),
.A2(n_1151),
.B1(n_1363),
.B2(n_1478),
.C1(n_1524),
.C2(n_1523),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1509),
.B(n_1439),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1454),
.A2(n_1045),
.B1(n_1229),
.B2(n_1520),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1467),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1484),
.A2(n_1151),
.B1(n_1251),
.B2(n_1248),
.Y(n_1631)
);

AOI22x1_ASAP7_75t_L g1632 ( 
.A1(n_1502),
.A2(n_1151),
.B1(n_900),
.B2(n_1326),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1454),
.A2(n_758),
.B1(n_874),
.B2(n_883),
.C(n_1229),
.Y(n_1633)
);

AO31x2_ASAP7_75t_L g1634 ( 
.A1(n_1515),
.A2(n_1528),
.A3(n_1432),
.B(n_1360),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1384),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_SL g1636 ( 
.A1(n_1460),
.A2(n_1418),
.B(n_1444),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_SL g1637 ( 
.A1(n_1460),
.A2(n_1418),
.B(n_1444),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1382),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1515),
.A2(n_1528),
.B(n_1045),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1419),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1384),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1454),
.A2(n_758),
.B1(n_874),
.B2(n_883),
.C(n_1229),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1515),
.A2(n_1528),
.B(n_1045),
.Y(n_1645)
);

OAI21xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1455),
.A2(n_1045),
.B(n_1219),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1382),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1382),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1454),
.B(n_1229),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1509),
.B(n_1439),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1384),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1419),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1533),
.B(n_1447),
.Y(n_1654)
);

AO32x2_ASAP7_75t_L g1655 ( 
.A1(n_1523),
.A2(n_1524),
.A3(n_1472),
.B1(n_1405),
.B2(n_1421),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1419),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1463),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1515),
.A2(n_1528),
.B(n_1045),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1419),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1382),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1382),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_SL g1665 ( 
.A1(n_1460),
.A2(n_1418),
.B(n_1444),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1447),
.B(n_1533),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1520),
.B(n_1535),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_SL g1669 ( 
.A1(n_1381),
.A2(n_1432),
.B(n_1477),
.C(n_1471),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1484),
.A2(n_1151),
.B1(n_1229),
.B2(n_1255),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1491),
.B(n_1400),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1419),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1520),
.B(n_1535),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_SL g1674 ( 
.A1(n_1381),
.A2(n_1432),
.B(n_1477),
.C(n_1471),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1461),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1447),
.B(n_1533),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1533),
.B(n_1447),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1521),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1454),
.B(n_1229),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1384),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1463),
.Y(n_1682)
);

CKINVDCx14_ASAP7_75t_R g1683 ( 
.A(n_1419),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1402),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1454),
.A2(n_1045),
.B(n_883),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1384),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1377),
.A2(n_1530),
.B(n_1525),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1484),
.A2(n_1151),
.B1(n_1229),
.B2(n_1255),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1384),
.Y(n_1689)
);

BUFx4f_ASAP7_75t_L g1690 ( 
.A(n_1461),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1463),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1484),
.A2(n_1151),
.B1(n_1251),
.B2(n_1248),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1586),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1586),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1599),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1633),
.A2(n_1644),
.B(n_1680),
.C(n_1649),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1629),
.B(n_1649),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1680),
.A2(n_1671),
.B(n_1565),
.Y(n_1698)
);

AOI31xp33_ASAP7_75t_L g1699 ( 
.A1(n_1631),
.A2(n_1692),
.A3(n_1541),
.B(n_1553),
.Y(n_1699)
);

CKINVDCx11_ASAP7_75t_R g1700 ( 
.A(n_1656),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1667),
.B(n_1676),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1685),
.B(n_1670),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1677),
.B(n_1591),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1605),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1646),
.A2(n_1669),
.B(n_1674),
.C(n_1544),
.Y(n_1705)
);

O2A1O1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1669),
.A2(n_1674),
.B(n_1626),
.C(n_1580),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1573),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1671),
.A2(n_1560),
.B(n_1668),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1624),
.A2(n_1622),
.B(n_1604),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1671),
.A2(n_1673),
.B(n_1668),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1569),
.A2(n_1670),
.B(n_1688),
.C(n_1555),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1583),
.B(n_1540),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1624),
.A2(n_1615),
.B(n_1602),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1673),
.A2(n_1587),
.B(n_1566),
.Y(n_1714)
);

BUFx12f_ASAP7_75t_L g1715 ( 
.A(n_1570),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1688),
.A2(n_1597),
.B1(n_1555),
.B2(n_1577),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1551),
.B(n_1606),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1597),
.A2(n_1577),
.B1(n_1568),
.B2(n_1567),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1538),
.B(n_1658),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1568),
.A2(n_1566),
.B1(n_1572),
.B2(n_1620),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1615),
.A2(n_1602),
.B(n_1576),
.Y(n_1721)
);

OA22x2_ASAP7_75t_L g1722 ( 
.A1(n_1600),
.A2(n_1594),
.B1(n_1572),
.B2(n_1665),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1605),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1572),
.A2(n_1620),
.B1(n_1579),
.B2(n_1625),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1625),
.A2(n_1690),
.B1(n_1691),
.B2(n_1682),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1563),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1562),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1589),
.A2(n_1637),
.B(n_1636),
.C(n_1614),
.Y(n_1729)
);

A2O1A1Ixp33_ASAP7_75t_SL g1730 ( 
.A1(n_1601),
.A2(n_1613),
.B(n_1684),
.C(n_1554),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1557),
.A2(n_1549),
.B(n_1623),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1539),
.Y(n_1732)
);

NOR2xp67_ASAP7_75t_L g1733 ( 
.A(n_1603),
.B(n_1559),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1679),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1690),
.A2(n_1632),
.B1(n_1592),
.B2(n_1581),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1563),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1595),
.A2(n_1542),
.B(n_1675),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1563),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1610),
.B(n_1552),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1575),
.B(n_1578),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1612),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1650),
.B(n_1552),
.Y(n_1742)
);

INVxp33_ASAP7_75t_L g1743 ( 
.A(n_1618),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1650),
.B(n_1561),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1593),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1571),
.B(n_1638),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1635),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1642),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1651),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1556),
.A2(n_1689),
.B1(n_1686),
.B2(n_1681),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1638),
.B(n_1647),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1647),
.B(n_1648),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1648),
.B(n_1663),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1595),
.B(n_1663),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1664),
.B(n_1609),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1664),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1590),
.B(n_1618),
.Y(n_1758)
);

AOI221x1_ASAP7_75t_SL g1759 ( 
.A1(n_1621),
.A2(n_1655),
.B1(n_1596),
.B2(n_1616),
.C(n_1584),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1617),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1596),
.B(n_1588),
.C(n_1546),
.Y(n_1761)
);

BUFx12f_ASAP7_75t_L g1762 ( 
.A(n_1570),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1608),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1590),
.B(n_1655),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1605),
.B(n_1617),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1588),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1630),
.B(n_1585),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1585),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1619),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1550),
.A2(n_1574),
.B(n_1564),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1582),
.A2(n_1630),
.B(n_1662),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1585),
.A2(n_1683),
.B1(n_1662),
.B2(n_1653),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1598),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1611),
.B(n_1634),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1598),
.B(n_1558),
.Y(n_1777)
);

OAI22x1_ASAP7_75t_L g1778 ( 
.A1(n_1548),
.A2(n_1641),
.B1(n_1672),
.B2(n_1656),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1558),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1640),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1548),
.B(n_1641),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1643),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1652),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1657),
.B(n_1678),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1659),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1672),
.B(n_1543),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1666),
.Y(n_1787)
);

INVx3_ASAP7_75t_SL g1788 ( 
.A(n_1627),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1660),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1687),
.B(n_1629),
.Y(n_1790)
);

CKINVDCx16_ASAP7_75t_R g1791 ( 
.A(n_1548),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1629),
.B(n_1668),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1545),
.B(n_1654),
.Y(n_1793)
);

NOR2xp67_ASAP7_75t_L g1794 ( 
.A(n_1583),
.B(n_989),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1649),
.A2(n_1680),
.B(n_1644),
.Y(n_1795)
);

AO21x2_ASAP7_75t_L g1796 ( 
.A1(n_1639),
.A2(n_1661),
.B(n_1645),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1667),
.B(n_1676),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1629),
.B(n_1668),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1649),
.A2(n_1680),
.B(n_1644),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1541),
.A2(n_1644),
.B1(n_1633),
.B2(n_1631),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1653),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1563),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1563),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1649),
.B(n_1680),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1583),
.B(n_989),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1541),
.A2(n_1644),
.B1(n_1633),
.B2(n_1631),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1639),
.A2(n_1661),
.B(n_1645),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1649),
.A2(n_1680),
.B(n_1644),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1629),
.B(n_1668),
.Y(n_1809)
);

O2A1O1Ixp5_ASAP7_75t_L g1810 ( 
.A1(n_1580),
.A2(n_1649),
.B(n_1680),
.C(n_1045),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1649),
.A2(n_1680),
.B(n_1644),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1633),
.A2(n_1644),
.B1(n_1541),
.B2(n_1631),
.Y(n_1812)
);

O2A1O1Ixp5_ASAP7_75t_L g1813 ( 
.A1(n_1580),
.A2(n_1649),
.B(n_1680),
.C(n_1045),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1545),
.B(n_1654),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1547),
.B(n_1628),
.Y(n_1815)
);

O2A1O1Ixp5_ASAP7_75t_L g1816 ( 
.A1(n_1580),
.A2(n_1649),
.B(n_1680),
.C(n_1045),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1764),
.B(n_1766),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1755),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1719),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1766),
.B(n_1771),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1708),
.B(n_1737),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1751),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1804),
.B(n_1717),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_SL g1824 ( 
.A(n_1761),
.B(n_1697),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1804),
.B(n_1712),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1696),
.B(n_1810),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1790),
.B(n_1707),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1728),
.B(n_1746),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1792),
.B(n_1798),
.Y(n_1829)
);

INVx6_ASAP7_75t_L g1830 ( 
.A(n_1760),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1740),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1809),
.B(n_1741),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1727),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1727),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_SL g1835 ( 
.A(n_1715),
.B(n_1762),
.Y(n_1835)
);

AO21x2_ASAP7_75t_L g1836 ( 
.A1(n_1730),
.A2(n_1779),
.B(n_1796),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1748),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1769),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1694),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1701),
.B(n_1797),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1749),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1736),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1738),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_R g1844 ( 
.A(n_1801),
.B(n_1791),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1763),
.B(n_1775),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1693),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1695),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1738),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1750),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1774),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1757),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1756),
.Y(n_1852)
);

BUFx12f_ASAP7_75t_L g1853 ( 
.A(n_1700),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1697),
.B(n_1703),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1786),
.B(n_1723),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1780),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1723),
.A2(n_1782),
.B(n_1787),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1787),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1786),
.B(n_1726),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1742),
.B(n_1745),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1793),
.B(n_1814),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1781),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_SL g1863 ( 
.A(n_1718),
.B(n_1725),
.Y(n_1863)
);

AO21x2_ASAP7_75t_L g1864 ( 
.A1(n_1702),
.A2(n_1777),
.B(n_1785),
.Y(n_1864)
);

OR2x4_ASAP7_75t_L g1865 ( 
.A(n_1699),
.B(n_1765),
.Y(n_1865)
);

OA21x2_ASAP7_75t_L g1866 ( 
.A1(n_1702),
.A2(n_1816),
.B(n_1813),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1758),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1795),
.B(n_1799),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1802),
.B(n_1803),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1803),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1744),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1747),
.Y(n_1872)
);

AO21x2_ASAP7_75t_L g1873 ( 
.A1(n_1711),
.A2(n_1784),
.B(n_1811),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1770),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1808),
.B(n_1739),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1732),
.B(n_1734),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1752),
.Y(n_1877)
);

AO21x2_ASAP7_75t_L g1878 ( 
.A1(n_1784),
.A2(n_1698),
.B(n_1716),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1789),
.B(n_1753),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1704),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1754),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1783),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1767),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1743),
.B(n_1722),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1743),
.B(n_1722),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1709),
.Y(n_1886)
);

BUFx2_ASAP7_75t_L g1887 ( 
.A(n_1788),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1817),
.B(n_1721),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1818),
.B(n_1759),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1849),
.Y(n_1892)
);

INVx4_ASAP7_75t_R g1893 ( 
.A(n_1880),
.Y(n_1893)
);

OR2x6_ASAP7_75t_L g1894 ( 
.A(n_1821),
.B(n_1714),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1857),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1887),
.Y(n_1896)
);

AND2x4_ASAP7_75t_SL g1897 ( 
.A(n_1821),
.B(n_1815),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1857),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1826),
.A2(n_1812),
.B1(n_1806),
.B2(n_1720),
.Y(n_1899)
);

OAI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1868),
.A2(n_1706),
.B1(n_1705),
.B2(n_1829),
.C(n_1866),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1855),
.B(n_1852),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1857),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1820),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1820),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1845),
.B(n_1713),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1882),
.B(n_1815),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1821),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1855),
.B(n_1710),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1864),
.B(n_1731),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1831),
.B(n_1788),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1839),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1839),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1842),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1845),
.B(n_1864),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1887),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_1731),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1845),
.B(n_1850),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1832),
.A2(n_1729),
.B1(n_1735),
.B2(n_1778),
.C(n_1773),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1837),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1819),
.B(n_1807),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1874),
.B(n_1807),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1874),
.Y(n_1922)
);

NOR3xp33_ASAP7_75t_SL g1923 ( 
.A(n_1900),
.B(n_1862),
.C(n_1875),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1899),
.A2(n_1873),
.B1(n_1821),
.B2(n_1878),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1899),
.A2(n_1794),
.B(n_1805),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1892),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1900),
.A2(n_1865),
.B1(n_1859),
.B2(n_1821),
.Y(n_1927)
);

AO21x2_ASAP7_75t_L g1928 ( 
.A1(n_1895),
.A2(n_1886),
.B(n_1836),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1918),
.A2(n_1865),
.B1(n_1859),
.B2(n_1822),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1918),
.A2(n_1854),
.B1(n_1825),
.B2(n_1835),
.C(n_1823),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1888),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1901),
.B(n_1840),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1892),
.Y(n_1933)
);

A2O1A1Ixp33_ASAP7_75t_L g1934 ( 
.A1(n_1908),
.A2(n_1863),
.B(n_1884),
.C(n_1885),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1896),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1891),
.B(n_1831),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1908),
.B(n_1867),
.Y(n_1937)
);

OAI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1890),
.A2(n_1866),
.B(n_1884),
.C(n_1885),
.Y(n_1938)
);

AO21x2_ASAP7_75t_L g1939 ( 
.A1(n_1895),
.A2(n_1886),
.B(n_1836),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1906),
.Y(n_1940)
);

CKINVDCx20_ASAP7_75t_R g1941 ( 
.A(n_1897),
.Y(n_1941)
);

BUFx10_ASAP7_75t_L g1942 ( 
.A(n_1906),
.Y(n_1942)
);

NAND2xp33_ASAP7_75t_R g1943 ( 
.A(n_1894),
.B(n_1844),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1890),
.B(n_1872),
.Y(n_1944)
);

OA222x2_ASAP7_75t_L g1945 ( 
.A1(n_1894),
.A2(n_1833),
.B1(n_1834),
.B2(n_1824),
.C1(n_1910),
.C2(n_1893),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1894),
.A2(n_1866),
.B1(n_1873),
.B2(n_1878),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1911),
.Y(n_1947)
);

AOI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1904),
.A2(n_1876),
.B1(n_1861),
.B2(n_1877),
.C(n_1871),
.Y(n_1948)
);

AOI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1904),
.A2(n_1861),
.B1(n_1871),
.B2(n_1881),
.C(n_1841),
.Y(n_1949)
);

AO21x1_ASAP7_75t_SL g1950 ( 
.A1(n_1910),
.A2(n_1827),
.B(n_1824),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1911),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1894),
.A2(n_1866),
.B1(n_1873),
.B2(n_1878),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1922),
.A2(n_1858),
.B(n_1856),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1903),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1903),
.B(n_1881),
.Y(n_1955)
);

AOI222xp33_ASAP7_75t_L g1956 ( 
.A1(n_1897),
.A2(n_1863),
.B1(n_1853),
.B2(n_1828),
.C1(n_1879),
.C2(n_1733),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1912),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1906),
.B(n_1917),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1894),
.A2(n_1865),
.B1(n_1830),
.B2(n_1880),
.Y(n_1959)
);

AOI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1914),
.A2(n_1841),
.B1(n_1828),
.B2(n_1879),
.C(n_1846),
.Y(n_1960)
);

INVxp67_ASAP7_75t_SL g1961 ( 
.A(n_1898),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1912),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1913),
.B(n_1883),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1896),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1894),
.A2(n_1830),
.B1(n_1880),
.B2(n_1772),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1919),
.B(n_1860),
.Y(n_1966)
);

OR2x6_ASAP7_75t_L g1967 ( 
.A(n_1907),
.B(n_1830),
.Y(n_1967)
);

OAI211xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1920),
.A2(n_1846),
.B(n_1847),
.C(n_1851),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1906),
.B(n_1869),
.Y(n_1969)
);

NOR4xp25_ASAP7_75t_SL g1970 ( 
.A(n_1896),
.B(n_1843),
.C(n_1870),
.D(n_1848),
.Y(n_1970)
);

OAI211xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1920),
.A2(n_1913),
.B(n_1909),
.C(n_1916),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1947),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1951),
.Y(n_1973)
);

NOR2x1p5_ASAP7_75t_L g1974 ( 
.A(n_1944),
.B(n_1853),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1957),
.Y(n_1975)
);

OA21x2_ASAP7_75t_L g1976 ( 
.A1(n_1961),
.A2(n_1952),
.B(n_1946),
.Y(n_1976)
);

INVx4_ASAP7_75t_SL g1977 ( 
.A(n_1967),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1923),
.B(n_1907),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_SL g1979 ( 
.A(n_1923),
.B(n_1915),
.C(n_1914),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1930),
.B(n_1776),
.Y(n_1980)
);

OA21x2_ASAP7_75t_L g1981 ( 
.A1(n_1961),
.A2(n_1916),
.B(n_1909),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1954),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1942),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1962),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1953),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1953),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1954),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1945),
.B(n_1914),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1948),
.B(n_1917),
.Y(n_1989)
);

BUFx8_ASAP7_75t_L g1990 ( 
.A(n_1938),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1926),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1935),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1933),
.Y(n_1993)
);

BUFx3_ASAP7_75t_L g1994 ( 
.A(n_1964),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1967),
.B(n_1905),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1950),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1931),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1936),
.B(n_1919),
.Y(n_1998)
);

INVx4_ASAP7_75t_SL g1999 ( 
.A(n_1967),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1931),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1937),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1955),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1932),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1946),
.A2(n_1916),
.B(n_1909),
.Y(n_2004)
);

OR2x6_ASAP7_75t_L g2005 ( 
.A(n_1965),
.B(n_1907),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1968),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1952),
.A2(n_1922),
.B(n_1921),
.Y(n_2007)
);

OA21x2_ASAP7_75t_L g2008 ( 
.A1(n_1934),
.A2(n_1902),
.B(n_1921),
.Y(n_2008)
);

NOR2xp67_ASAP7_75t_L g2009 ( 
.A(n_1924),
.B(n_1907),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1966),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1958),
.B(n_1889),
.Y(n_2011)
);

OA21x2_ASAP7_75t_L g2012 ( 
.A1(n_1934),
.A2(n_1902),
.B(n_1921),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1928),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1963),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1977),
.B(n_1940),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1994),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1996),
.B(n_1969),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_1929),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2006),
.B(n_1949),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1972),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1996),
.B(n_1940),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1996),
.B(n_1942),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1972),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1987),
.B(n_1982),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1996),
.B(n_1977),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1994),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2002),
.B(n_1960),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1996),
.B(n_1970),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1973),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1973),
.Y(n_2030)
);

AND2x4_ASAP7_75t_SL g2031 ( 
.A(n_1992),
.B(n_1941),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2002),
.B(n_2010),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1975),
.Y(n_2033)
);

HB1xp67_ASAP7_75t_L g2034 ( 
.A(n_2003),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1975),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1984),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1980),
.B(n_1925),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1984),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1977),
.B(n_1905),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1999),
.B(n_1988),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1998),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_1999),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1989),
.B(n_1927),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1981),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1997),
.B(n_1939),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1985),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1983),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1985),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1999),
.B(n_1988),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_2009),
.B(n_1956),
.Y(n_2050)
);

XNOR2x1_ASAP7_75t_L g2051 ( 
.A(n_1974),
.B(n_1959),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1991),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1991),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1986),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2025),
.B(n_1995),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2019),
.B(n_1974),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2025),
.B(n_2008),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2035),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2046),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2036),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2018),
.B(n_2011),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_L g2062 ( 
.A(n_2042),
.B(n_1978),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2024),
.B(n_1997),
.Y(n_2063)
);

AND3x2_ASAP7_75t_L g2064 ( 
.A(n_2040),
.B(n_2049),
.C(n_2028),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2040),
.B(n_2008),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2020),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2020),
.Y(n_2067)
);

NOR2x1p5_ASAP7_75t_L g2068 ( 
.A(n_2049),
.B(n_1979),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2046),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2024),
.B(n_2000),
.Y(n_2070)
);

INVxp67_ASAP7_75t_L g2071 ( 
.A(n_2034),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2017),
.B(n_2008),
.Y(n_2072)
);

O2A1O1Ixp5_ASAP7_75t_R g2073 ( 
.A1(n_2043),
.A2(n_1990),
.B(n_1976),
.C(n_2012),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2023),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2037),
.B(n_2011),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2023),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2017),
.B(n_2008),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2014),
.B(n_1993),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2079)
);

AND2x4_ASAP7_75t_SL g2080 ( 
.A(n_2015),
.B(n_2005),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2046),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2029),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2029),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2027),
.B(n_2000),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2030),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2014),
.B(n_2041),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2048),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2021),
.B(n_2012),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_2050),
.A2(n_2004),
.B(n_1971),
.C(n_2007),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2030),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2033),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2016),
.B(n_1993),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2031),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2021),
.B(n_2005),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2042),
.B(n_2005),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2033),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2090),
.A2(n_2051),
.B(n_2062),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_SL g2100 ( 
.A(n_2073),
.B(n_2028),
.C(n_2027),
.Y(n_2100)
);

AND3x1_ASAP7_75t_L g2101 ( 
.A(n_2073),
.B(n_2026),
.C(n_2016),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_2071),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2059),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_2056),
.B(n_2051),
.Y(n_2104)
);

NOR2x1_ASAP7_75t_L g2105 ( 
.A(n_2068),
.B(n_2044),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2055),
.Y(n_2106)
);

AO21x2_ASAP7_75t_L g2107 ( 
.A1(n_2065),
.A2(n_2013),
.B(n_2048),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2059),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2063),
.B(n_2032),
.Y(n_2109)
);

NOR2x1_ASAP7_75t_L g2110 ( 
.A(n_2068),
.B(n_2044),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2066),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2055),
.B(n_2047),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2080),
.B(n_2015),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2086),
.A2(n_2026),
.B(n_2031),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2095),
.B(n_2047),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2064),
.B(n_2031),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2058),
.B(n_2038),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2096),
.B(n_2015),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2066),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_2096),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2067),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2058),
.B(n_2038),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2060),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_2097),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2080),
.B(n_2015),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2080),
.B(n_2097),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_2060),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2067),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2124),
.B(n_2120),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2127),
.Y(n_2130)
);

NAND3x2_ASAP7_75t_L g2131 ( 
.A(n_2120),
.B(n_2084),
.C(n_2065),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2106),
.Y(n_2133)
);

NAND2x1p5_ASAP7_75t_L g2134 ( 
.A(n_2105),
.B(n_1704),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2124),
.B(n_2061),
.Y(n_2135)
);

NAND3xp33_ASAP7_75t_L g2136 ( 
.A(n_2099),
.B(n_1990),
.C(n_2084),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2106),
.B(n_2075),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2112),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_2105),
.B(n_2110),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2127),
.Y(n_2140)
);

AND2x2_ASAP7_75t_SL g2141 ( 
.A(n_2104),
.B(n_2057),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2112),
.B(n_2057),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2126),
.B(n_2089),
.Y(n_2143)
);

O2A1O1Ixp33_ASAP7_75t_SL g2144 ( 
.A1(n_2100),
.A2(n_2094),
.B(n_2044),
.C(n_2076),
.Y(n_2144)
);

AOI31xp33_ASAP7_75t_SL g2145 ( 
.A1(n_2116),
.A2(n_2070),
.A3(n_2063),
.B(n_2078),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2126),
.B(n_2089),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_2110),
.A2(n_2077),
.B(n_2072),
.C(n_2079),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2115),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2113),
.B(n_2074),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2123),
.Y(n_2150)
);

OAI21xp33_ASAP7_75t_L g2151 ( 
.A1(n_2115),
.A2(n_2077),
.B(n_2072),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2102),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2133),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2133),
.B(n_2113),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_2130),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2148),
.B(n_2118),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2139),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2138),
.B(n_2114),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_2149),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2143),
.B(n_2118),
.Y(n_2160)
);

INVxp67_ASAP7_75t_SL g2161 ( 
.A(n_2139),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2134),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_2141),
.A2(n_1990),
.B1(n_2125),
.B2(n_2113),
.Y(n_2163)
);

INVx2_ASAP7_75t_SL g2164 ( 
.A(n_2149),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2138),
.B(n_2113),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2152),
.B(n_2125),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2136),
.A2(n_2141),
.B1(n_2125),
.B2(n_2101),
.Y(n_2167)
);

OAI211xp5_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_2131),
.B(n_2144),
.C(n_2129),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2163),
.B(n_2125),
.Y(n_2169)
);

AOI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_2161),
.A2(n_2145),
.B(n_2144),
.C(n_2147),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2163),
.A2(n_2161),
.B1(n_2101),
.B2(n_2157),
.Y(n_2171)
);

OAI211xp5_ASAP7_75t_L g2172 ( 
.A1(n_2157),
.A2(n_2166),
.B(n_2158),
.C(n_2147),
.Y(n_2172)
);

NOR3xp33_ASAP7_75t_SL g2173 ( 
.A(n_2166),
.B(n_2137),
.C(n_2150),
.Y(n_2173)
);

AOI221xp5_ASAP7_75t_L g2174 ( 
.A1(n_2154),
.A2(n_2140),
.B1(n_2132),
.B2(n_2151),
.C(n_2143),
.Y(n_2174)
);

OAI211xp5_ASAP7_75t_SL g2175 ( 
.A1(n_2165),
.A2(n_2135),
.B(n_2162),
.C(n_2153),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2154),
.B(n_2149),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2159),
.B(n_2146),
.Y(n_2177)
);

AOI211x1_ASAP7_75t_L g2178 ( 
.A1(n_2160),
.A2(n_2156),
.B(n_2146),
.C(n_2142),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2164),
.A2(n_2134),
.B(n_2117),
.Y(n_2179)
);

O2A1O1Ixp5_ASAP7_75t_L g2180 ( 
.A1(n_2155),
.A2(n_2122),
.B(n_2142),
.C(n_2103),
.Y(n_2180)
);

NAND2x1_ASAP7_75t_L g2181 ( 
.A(n_2155),
.B(n_2103),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2181),
.Y(n_2182)
);

NOR2x1_ASAP7_75t_L g2183 ( 
.A(n_2172),
.B(n_2155),
.Y(n_2183)
);

AOI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2171),
.A2(n_2155),
.B1(n_2122),
.B2(n_2128),
.C(n_2121),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2170),
.A2(n_2128),
.B(n_2119),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2178),
.B(n_2109),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2176),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2177),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2187),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2183),
.B(n_2174),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2188),
.B(n_2173),
.Y(n_2191)
);

NOR2x1_ASAP7_75t_L g2192 ( 
.A(n_2182),
.B(n_2175),
.Y(n_2192)
);

NOR2xp67_ASAP7_75t_L g2193 ( 
.A(n_2185),
.B(n_2179),
.Y(n_2193)
);

OAI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2186),
.A2(n_2168),
.B(n_2169),
.Y(n_2194)
);

NOR3xp33_ASAP7_75t_L g2195 ( 
.A(n_2184),
.B(n_2180),
.C(n_2119),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2183),
.Y(n_2196)
);

AOI222xp33_ASAP7_75t_L g2197 ( 
.A1(n_2194),
.A2(n_2111),
.B1(n_2121),
.B2(n_2103),
.C1(n_2108),
.C2(n_2087),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_2192),
.B(n_2111),
.C(n_2108),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2196),
.Y(n_2199)
);

INVxp33_ASAP7_75t_L g2200 ( 
.A(n_2190),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_2191),
.Y(n_2201)
);

A2O1A1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2193),
.A2(n_2109),
.B(n_2108),
.C(n_2079),
.Y(n_2202)
);

OAI332xp33_ASAP7_75t_L g2203 ( 
.A1(n_2189),
.A2(n_2081),
.A3(n_2088),
.B1(n_2069),
.B2(n_2091),
.B3(n_2093),
.C1(n_2092),
.C2(n_2076),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2199),
.Y(n_2204)
);

INVx2_ASAP7_75t_SL g2205 ( 
.A(n_2198),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2201),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2197),
.B(n_2195),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_2202),
.B(n_2087),
.C(n_2081),
.Y(n_2208)
);

NOR2x1_ASAP7_75t_L g2209 ( 
.A(n_2206),
.B(n_2200),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2204),
.B(n_2070),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2205),
.Y(n_2211)
);

AOI322xp5_ASAP7_75t_L g2212 ( 
.A1(n_2209),
.A2(n_2207),
.A3(n_2208),
.B1(n_2044),
.B2(n_2203),
.C1(n_2069),
.C2(n_2088),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2210),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_2213),
.Y(n_2214)
);

NOR2xp67_ASAP7_75t_L g2215 ( 
.A(n_2212),
.B(n_2211),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2213),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2216),
.A2(n_2091),
.B1(n_2107),
.B2(n_2093),
.Y(n_2217)
);

INVxp67_ASAP7_75t_L g2218 ( 
.A(n_2214),
.Y(n_2218)
);

OAI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2215),
.A2(n_2083),
.B1(n_2098),
.B2(n_2092),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2218),
.A2(n_2082),
.B1(n_2098),
.B2(n_2085),
.Y(n_2220)
);

OAI22x1_ASAP7_75t_L g2221 ( 
.A1(n_2220),
.A2(n_2219),
.B1(n_2217),
.B2(n_2082),
.Y(n_2221)
);

AOI21x1_ASAP7_75t_L g2222 ( 
.A1(n_2221),
.A2(n_2083),
.B(n_2074),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_2222),
.B(n_2085),
.Y(n_2223)
);

AOI31xp33_ASAP7_75t_L g2224 ( 
.A1(n_2223),
.A2(n_1943),
.A3(n_1768),
.B(n_2039),
.Y(n_2224)
);

AOI221xp5_ASAP7_75t_L g2225 ( 
.A1(n_2224),
.A2(n_2107),
.B1(n_2054),
.B2(n_2053),
.C(n_2052),
.Y(n_2225)
);

AOI211xp5_ASAP7_75t_L g2226 ( 
.A1(n_2225),
.A2(n_1724),
.B(n_2054),
.C(n_2045),
.Y(n_2226)
);


endmodule