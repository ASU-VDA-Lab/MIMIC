module fake_ariane_3099_n_1924 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1924);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1924;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_42),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_23),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_123),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_37),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_127),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_95),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_20),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_52),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_0),
.Y(n_188)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_20),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_93),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_87),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_4),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_89),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_47),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_57),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_71),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_113),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_112),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_31),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_19),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_39),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_2),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_125),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_69),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_23),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_90),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_118),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_24),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_37),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_126),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_133),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_73),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_60),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_96),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_82),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_65),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_48),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_32),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_41),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_40),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_77),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_68),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_101),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_25),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_43),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_29),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_24),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_8),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_108),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_140),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_117),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_67),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_156),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_149),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_50),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_34),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_63),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_51),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_99),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_7),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_26),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_70),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_64),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_26),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_6),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_12),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_19),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_98),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_137),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_151),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_72),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_34),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_7),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_44),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_11),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_111),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_85),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_167),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_271),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_168),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_175),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_285),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_229),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_206),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_217),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_177),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_229),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_196),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_217),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_217),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_187),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_197),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_169),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_227),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_233),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_208),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_278),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_190),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_274),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_281),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_234),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_234),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_260),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_197),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_260),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_218),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_263),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_263),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_280),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_193),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_170),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_193),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_280),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_170),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_280),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_218),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_173),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_290),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_158),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_237),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_173),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_232),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_164),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_174),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_174),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_165),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_176),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_171),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_171),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_381),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_290),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_378),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_237),
.B1(n_266),
.B2(n_306),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_290),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_372),
.B(n_213),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_351),
.B(n_159),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_338),
.A2(n_266),
.B1(n_306),
.B2(n_296),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_372),
.B(n_213),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_367),
.A2(n_223),
.B1(n_264),
.B2(n_239),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_326),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_386),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_369),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_389),
.A2(n_180),
.B(n_172),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_335),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_379),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_315),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_366),
.B(n_210),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_318),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_332),
.Y(n_438)
);

AND2x2_ASAP7_75t_SL g439 ( 
.A(n_370),
.B(n_232),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_361),
.B(n_187),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_365),
.B(n_313),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_323),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_363),
.B(n_249),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_354),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_324),
.B(n_249),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_328),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_341),
.B(n_300),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_342),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_354),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_344),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_321),
.A2(n_286),
.B1(n_225),
.B2(n_309),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_350),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_439),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_403),
.B1(n_393),
.B2(n_396),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_439),
.B(n_376),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_439),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_426),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_442),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

AND3x2_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_345),
.C(n_265),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_426),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_393),
.B(n_376),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_442),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_380),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_396),
.B(n_380),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_373),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_405),
.A2(n_182),
.B(n_181),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_405),
.B(n_317),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_423),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_397),
.B(n_355),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_396),
.B(n_353),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_416),
.B(n_356),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_411),
.B(n_320),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_403),
.A2(n_339),
.B1(n_347),
.B2(n_375),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_444),
.A2(n_347),
.B1(n_385),
.B2(n_384),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_411),
.A2(n_374),
.B1(n_359),
.B2(n_358),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_442),
.B(n_320),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

CKINVDCx6p67_ASAP7_75t_R g512 ( 
.A(n_444),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_454),
.B(n_384),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_415),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_406),
.B(n_443),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_456),
.B(n_300),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_408),
.A2(n_387),
.B1(n_385),
.B2(n_261),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_444),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_398),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_416),
.B(n_454),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_SL g523 ( 
.A1(n_444),
.A2(n_186),
.B(n_185),
.Y(n_523)
);

CKINVDCx6p67_ASAP7_75t_R g524 ( 
.A(n_418),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_416),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_397),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_399),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_421),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_406),
.B(n_387),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_401),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_416),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_443),
.B(n_176),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_401),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_416),
.B(n_178),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_443),
.B(n_179),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_454),
.B(n_355),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_456),
.B(n_246),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_454),
.B(n_179),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_414),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_454),
.B(n_455),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_455),
.B(n_248),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_440),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_427),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_408),
.A2(n_269),
.B1(n_188),
.B2(n_198),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_455),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_455),
.B(n_248),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_404),
.B(n_364),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_455),
.B(n_284),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_400),
.B(n_364),
.C(n_307),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_424),
.A2(n_244),
.B1(n_183),
.B2(n_252),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_400),
.A2(n_362),
.B1(n_357),
.B2(n_343),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_440),
.B(n_262),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_437),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_424),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_424),
.A2(n_242),
.B1(n_253),
.B2(n_256),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_425),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_203),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_R g576 ( 
.A(n_438),
.B(n_322),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_430),
.B(n_207),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_451),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_391),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_425),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_391),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_425),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_391),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_451),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_448),
.B(n_284),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_391),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_448),
.B(n_287),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_391),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_390),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_434),
.B(n_287),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_448),
.B(n_294),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_418),
.B(n_294),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_390),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_446),
.A2(n_228),
.B1(n_259),
.B2(n_235),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_390),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_392),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_392),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_392),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_402),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_447),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_418),
.B(n_451),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_450),
.A2(n_209),
.B1(n_275),
.B2(n_214),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

NOR2x1p5_ASAP7_75t_L g606 ( 
.A(n_452),
.B(n_430),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_450),
.B(n_301),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_451),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_489),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_514),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_466),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_461),
.A2(n_435),
.B1(n_436),
.B2(n_441),
.Y(n_615)
);

AND2x2_ASAP7_75t_SL g616 ( 
.A(n_567),
.B(n_573),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_486),
.B(n_433),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_460),
.B(n_451),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_L g619 ( 
.A1(n_543),
.A2(n_485),
.B(n_484),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_565),
.B(n_211),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_497),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_460),
.B(n_457),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_525),
.A2(n_449),
.B1(n_445),
.B2(n_432),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_466),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_545),
.B(n_435),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_506),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_506),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_564),
.A2(n_221),
.B(n_236),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_514),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_511),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_471),
.B(n_457),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_511),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_520),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_471),
.B(n_457),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_520),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_535),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_508),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_473),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_522),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_537),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_464),
.B(n_436),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_602),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_480),
.B(n_441),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_474),
.B(n_457),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_473),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_473),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_522),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_576),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_457),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_494),
.B(n_433),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_450),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_474),
.B(n_457),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_566),
.B(n_432),
.Y(n_660)
);

AOI22x1_ASAP7_75t_L g661 ( 
.A1(n_558),
.A2(n_449),
.B1(n_445),
.B2(n_453),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_542),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_566),
.B(n_453),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_527),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_527),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_494),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_542),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_481),
.B(n_457),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_544),
.A2(n_413),
.B1(n_453),
.B2(n_458),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_481),
.B(n_446),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_547),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_602),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_534),
.B(n_446),
.Y(n_673)
);

NAND3x1_ASAP7_75t_L g674 ( 
.A(n_604),
.B(n_340),
.C(n_333),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_496),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_561),
.B(n_526),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_486),
.B(n_446),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_548),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_525),
.B(n_301),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_524),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_531),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_496),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_561),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_519),
.B(n_304),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_550),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_513),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_531),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_538),
.Y(n_691)
);

INVx3_ASAP7_75t_R g692 ( 
.A(n_568),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_486),
.B(n_446),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_523),
.A2(n_458),
.B1(n_304),
.B2(n_428),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_540),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_534),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_473),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_524),
.B(n_458),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_486),
.B(n_498),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_550),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_534),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_498),
.B(n_428),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_483),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_499),
.B(n_429),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_540),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_483),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_553),
.B(n_429),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_473),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_523),
.B(n_571),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_499),
.B(n_325),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_492),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_492),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_534),
.B(n_219),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_517),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_553),
.B(n_240),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_555),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_555),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_502),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_501),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_586),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_501),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_503),
.A2(n_276),
.B1(n_257),
.B2(n_413),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_504),
.B(n_254),
.Y(n_724)
);

BUFx4f_ASAP7_75t_L g725 ( 
.A(n_512),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_255),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_459),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_507),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_459),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_588),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_419),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_462),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_579),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_606),
.B(n_419),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_492),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_507),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_463),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_604),
.B(n_431),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_477),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_521),
.B(n_273),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_509),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_551),
.B(n_289),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_515),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_463),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_295),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_592),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_462),
.B(n_302),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_465),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_491),
.A2(n_303),
.B1(n_241),
.B2(n_195),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_509),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_516),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_516),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_465),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_468),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_512),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_462),
.B(n_467),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_518),
.B(n_431),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_468),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_467),
.B(n_262),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_467),
.B(n_262),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_2),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_528),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_572),
.B(n_232),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_475),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_544),
.A2(n_166),
.B1(n_163),
.B2(n_160),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_472),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_492),
.B(n_262),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_492),
.B(n_262),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_591),
.B(n_3),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_544),
.A2(n_517),
.B1(n_572),
.B2(n_557),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_539),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_472),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_607),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_475),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_518),
.B(n_8),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_528),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_557),
.B(n_9),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_469),
.B(n_402),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_517),
.B(n_10),
.Y(n_779)
);

AO21x2_ASAP7_75t_L g780 ( 
.A1(n_596),
.A2(n_488),
.B(n_578),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_701),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_642),
.Y(n_783)
);

AND2x6_ASAP7_75t_L g784 ( 
.A(n_678),
.B(n_470),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_609),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_696),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_610),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_613),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_724),
.A2(n_643),
.B1(n_699),
.B2(n_770),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_688),
.A2(n_595),
.B1(n_544),
.B2(n_577),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_646),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_643),
.B(n_575),
.C(n_559),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_611),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_731),
.B(n_734),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_612),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_688),
.B(n_475),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_617),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_622),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_621),
.B(n_624),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_629),
.B(n_493),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_653),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_633),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_630),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_696),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_635),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_732),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_622),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_638),
.B(n_493),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_639),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_641),
.B(n_493),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_SL g811 ( 
.A(n_685),
.B(n_593),
.C(n_536),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_645),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_654),
.B(n_500),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_648),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_699),
.B(n_529),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_756),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_732),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_756),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_685),
.B(n_541),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_724),
.A2(n_517),
.B1(n_488),
.B2(n_552),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_665),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_672),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_628),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_619),
.A2(n_479),
.B(n_470),
.C(n_476),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_616),
.A2(n_488),
.B1(n_530),
.B2(n_533),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_662),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_667),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_672),
.Y(n_828)
);

BUFx8_ASAP7_75t_SL g829 ( 
.A(n_655),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_678),
.B(n_500),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_SL g831 ( 
.A1(n_692),
.A2(n_505),
.B1(n_308),
.B2(n_283),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_677),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_698),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_770),
.A2(n_546),
.B1(n_562),
.B2(n_500),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_657),
.B(n_666),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_765),
.B(n_649),
.C(n_723),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_683),
.B(n_476),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_773),
.B(n_579),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_682),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_671),
.Y(n_840)
);

CKINVDCx16_ASAP7_75t_R g841 ( 
.A(n_617),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_759),
.A2(n_479),
.B(n_482),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_689),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_759),
.A2(n_482),
.B(n_596),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_627),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_617),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_690),
.B(n_530),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_691),
.Y(n_848)
);

OR2x2_ASAP7_75t_SL g849 ( 
.A(n_777),
.B(n_584),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_695),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_675),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_693),
.B(n_755),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_679),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_705),
.B(n_532),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_681),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_660),
.B(n_495),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_755),
.B(n_579),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_702),
.B(n_581),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_719),
.B(n_495),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_647),
.A2(n_585),
.B1(n_608),
.B2(n_605),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_616),
.A2(n_532),
.B1(n_533),
.B2(n_605),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_627),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_687),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_627),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_716),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_717),
.B(n_581),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_718),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_719),
.B(n_495),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_727),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_631),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_729),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_731),
.B(n_10),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_725),
.B(n_585),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_631),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_710),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_647),
.A2(n_585),
.B1(n_608),
.B2(n_495),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_760),
.A2(n_608),
.B(n_584),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_725),
.B(n_495),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_734),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_721),
.B(n_730),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_721),
.B(n_581),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_737),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_702),
.B(n_589),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_744),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_773),
.B(n_510),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_700),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_765),
.B(n_510),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_666),
.B(n_589),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_761),
.A2(n_589),
.B(n_587),
.C(n_563),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_714),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_730),
.B(n_510),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_703),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_660),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_746),
.B(n_587),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_714),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_746),
.B(n_510),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_669),
.A2(n_510),
.B1(n_549),
.B2(n_554),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_738),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_709),
.A2(n_569),
.B(n_560),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_631),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_669),
.A2(n_549),
.B1(n_554),
.B2(n_599),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_634),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_771),
.B(n_560),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_757),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_748),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_753),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_775),
.A2(n_549),
.B1(n_554),
.B2(n_599),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_634),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_754),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_769),
.A2(n_549),
.B1(n_554),
.B2(n_598),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_769),
.A2(n_549),
.B1(n_554),
.B2(n_598),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_714),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_634),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_739),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_733),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_706),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_743),
.B(n_563),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_570),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_SL g919 ( 
.A1(n_713),
.A2(n_569),
.B(n_582),
.C(n_570),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_658),
.A2(n_590),
.B1(n_600),
.B2(n_597),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_673),
.B(n_574),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_673),
.B(n_574),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_704),
.B(n_779),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_758),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_766),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_658),
.B(n_580),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_704),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_772),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_615),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_649),
.A2(n_580),
.B1(n_583),
.B2(n_582),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_658),
.B(n_583),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_658),
.B(n_590),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_713),
.B(n_594),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_749),
.B(n_201),
.C(n_310),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_620),
.A2(n_601),
.B1(n_600),
.B2(n_597),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_676),
.B(n_594),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_720),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_723),
.B(n_194),
.C(n_282),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_722),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_620),
.B(n_601),
.Y(n_940)
);

AND2x6_ASAP7_75t_SL g941 ( 
.A(n_761),
.B(n_715),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_660),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_686),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_764),
.B(n_262),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_686),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_764),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_SL g948 ( 
.A(n_625),
.B(n_707),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_670),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_650),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_650),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_774),
.B(n_262),
.Y(n_952)
);

BUFx4f_ASAP7_75t_L g953 ( 
.A(n_745),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_745),
.B(n_625),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_659),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_659),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_670),
.B(n_13),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_680),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_715),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_774),
.B(n_402),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_668),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_674),
.B(n_313),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_668),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_736),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_707),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_747),
.B(n_313),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_614),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_676),
.B(n_243),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_694),
.A2(n_660),
.B1(n_751),
.B2(n_776),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_741),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_750),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_781),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_833),
.B(n_747),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_740),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_833),
.B(n_636),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_781),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_959),
.B(n_740),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_856),
.Y(n_978)
);

AND3x2_ASAP7_75t_SL g979 ( 
.A(n_836),
.B(n_626),
.C(n_637),
.Y(n_979)
);

CKINVDCx8_ASAP7_75t_R g980 ( 
.A(n_788),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_949),
.B(n_726),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_781),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_929),
.B(n_684),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_789),
.A2(n_709),
.B(n_726),
.C(n_742),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_814),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_802),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_783),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_785),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_829),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_782),
.B(n_684),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_852),
.B(n_890),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_852),
.B(n_644),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_787),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_895),
.B(n_644),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_950),
.B(n_742),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_798),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_839),
.Y(n_997)
);

NOR2x2_ASAP7_75t_L g998 ( 
.A(n_962),
.B(n_752),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_823),
.B(n_632),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_807),
.Y(n_1000)
);

BUFx2_ASAP7_75t_SL g1001 ( 
.A(n_782),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_880),
.B(n_663),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_927),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_875),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_880),
.B(n_663),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_782),
.B(n_644),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_832),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_793),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_790),
.A2(n_632),
.B(n_661),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_835),
.Y(n_1010)
);

CKINVDCx8_ASAP7_75t_R g1011 ( 
.A(n_794),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_791),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_831),
.A2(n_663),
.B1(n_640),
.B2(n_623),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_951),
.B(n_663),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_795),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_845),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_898),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_790),
.A2(n_618),
.B1(n_623),
.B2(n_640),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_955),
.B(n_956),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_803),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_820),
.A2(n_618),
.B(n_760),
.C(n_768),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_801),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_826),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_904),
.B(n_762),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_805),
.Y(n_1026)
);

CKINVDCx14_ASAP7_75t_R g1027 ( 
.A(n_797),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_953),
.B(n_651),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_SL g1029 ( 
.A1(n_962),
.A2(n_763),
.B1(n_656),
.B2(n_636),
.Y(n_1029)
);

AND3x1_ASAP7_75t_SL g1030 ( 
.A(n_809),
.B(n_13),
.C(n_14),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_953),
.B(n_651),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_961),
.B(n_656),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_827),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_786),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_893),
.B(n_651),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_840),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_963),
.B(n_799),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_812),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_944),
.A2(n_763),
.B1(n_652),
.B2(n_712),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_843),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_799),
.A2(n_652),
.B1(n_697),
.B2(n_708),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_848),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_778),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_851),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_923),
.B(n_778),
.Y(n_1045)
);

INVx6_ASAP7_75t_L g1046 ( 
.A(n_841),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_849),
.B(n_780),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_797),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_821),
.B(n_652),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_821),
.B(n_697),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_845),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_828),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_879),
.B(n_815),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_893),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_850),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_853),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_858),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_893),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_838),
.B(n_697),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_908),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_865),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_846),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_855),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_815),
.B(n_780),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_867),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_869),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_893),
.B(n_708),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_819),
.B(n_708),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_914),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_938),
.B(n_768),
.C(n_767),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_796),
.B(n_735),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_796),
.B(n_735),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_871),
.Y(n_1073)
);

AND3x1_ASAP7_75t_SL g1074 ( 
.A(n_882),
.B(n_14),
.C(n_15),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_858),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_863),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_948),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_845),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_884),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_942),
.B(n_711),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_946),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_881),
.B(n_735),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_941),
.B(n_712),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_905),
.B(n_906),
.Y(n_1084)
);

CKINVDCx12_ASAP7_75t_R g1085 ( 
.A(n_962),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_942),
.B(n_711),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_870),
.Y(n_1087)
);

INVxp33_ASAP7_75t_L g1088 ( 
.A(n_967),
.Y(n_1088)
);

AOI21xp33_ASAP7_75t_L g1089 ( 
.A1(n_954),
.A2(n_767),
.B(n_712),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_870),
.Y(n_1090)
);

BUFx8_ASAP7_75t_L g1091 ( 
.A(n_870),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_909),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_940),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_924),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_925),
.B(n_711),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_883),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_811),
.B(n_763),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_886),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_928),
.B(n_763),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_894),
.B(n_800),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_912),
.B(n_16),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_313),
.Y(n_1102)
);

INVxp33_ASAP7_75t_L g1103 ( 
.A(n_883),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_SL g1104 ( 
.A(n_857),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_888),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_786),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_874),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_894),
.B(n_17),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_800),
.B(n_17),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_804),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_808),
.B(n_18),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_942),
.B(n_202),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_892),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_916),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_SL g1115 ( 
.A1(n_957),
.A2(n_232),
.B1(n_312),
.B2(n_204),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_808),
.B(n_21),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_810),
.B(n_21),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_874),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_810),
.B(n_33),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_857),
.B(n_36),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_874),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_942),
.B(n_36),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_813),
.B(n_38),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_937),
.A2(n_312),
.B1(n_247),
.B2(n_279),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_983),
.B(n_1103),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1010),
.B(n_915),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1054),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1054),
.B(n_1058),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_988),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1054),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_987),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_985),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_993),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1012),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1004),
.B(n_915),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_974),
.B(n_903),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1008),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1077),
.A2(n_919),
.B(n_813),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_1054),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1120),
.A2(n_966),
.B1(n_872),
.B2(n_792),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_997),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1077),
.A2(n_889),
.B(n_854),
.Y(n_1142)
);

NOR2x1_ASAP7_75t_SL g1143 ( 
.A(n_1058),
.B(n_966),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_975),
.B(n_900),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_974),
.B(n_903),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1023),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1015),
.Y(n_1147)
);

BUFx2_ASAP7_75t_SL g1148 ( 
.A(n_980),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1058),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1021),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_984),
.A2(n_792),
.B(n_934),
.C(n_834),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1091),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1026),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_989),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1091),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_SL g1156 ( 
.A1(n_1037),
.A2(n_837),
.B(n_854),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1024),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1058),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1041),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1046),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1016),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1046),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1038),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_978),
.B(n_816),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1016),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1096),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1040),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1042),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1037),
.B(n_918),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1055),
.Y(n_1170)
);

NAND2x1p5_ASAP7_75t_L g1171 ( 
.A(n_992),
.B(n_900),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_975),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1016),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1081),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1061),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_975),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1027),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1033),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_986),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1060),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1065),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_995),
.B(n_918),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1100),
.A2(n_847),
.B(n_887),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1007),
.B(n_864),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1066),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_973),
.B(n_902),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1018),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_973),
.B(n_902),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_973),
.B(n_864),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1036),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_999),
.A2(n_970),
.B1(n_933),
.B2(n_971),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1009),
.A2(n_897),
.B(n_907),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1009),
.A2(n_896),
.B(n_891),
.C(n_969),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1052),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1100),
.A2(n_847),
.B(n_842),
.Y(n_1195)
);

AO21x2_ASAP7_75t_L g1196 ( 
.A1(n_1022),
.A2(n_899),
.B(n_842),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1051),
.Y(n_1197)
);

BUFx12f_ASAP7_75t_L g1198 ( 
.A(n_1069),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1017),
.Y(n_1199)
);

OAI222xp33_ASAP7_75t_L g1200 ( 
.A1(n_1019),
.A2(n_911),
.B1(n_910),
.B2(n_825),
.C1(n_861),
.C2(n_837),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1122),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1051),
.Y(n_1202)
);

AND2x6_ASAP7_75t_L g1203 ( 
.A(n_1122),
.B(n_818),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_981),
.A2(n_876),
.B(n_860),
.C(n_885),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1064),
.A2(n_964),
.B1(n_939),
.B2(n_943),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1075),
.B(n_913),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1051),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1120),
.A2(n_784),
.B1(n_830),
.B2(n_958),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_992),
.B(n_784),
.Y(n_1209)
);

INVx6_ASAP7_75t_L g1210 ( 
.A(n_982),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1044),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1053),
.B(n_913),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_977),
.A2(n_901),
.B1(n_784),
.B2(n_917),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1075),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_995),
.B(n_947),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1057),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1000),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_981),
.A2(n_866),
.B1(n_947),
.B2(n_920),
.Y(n_1218)
);

BUFx8_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1104),
.A2(n_1047),
.B1(n_1063),
.B2(n_1098),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_996),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_982),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1048),
.B(n_1043),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1070),
.A2(n_824),
.B(n_899),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1073),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1101),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1003),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1078),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1090),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1041),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1105),
.B(n_913),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1056),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1076),
.A2(n_784),
.B1(n_932),
.B2(n_936),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1011),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1109),
.A2(n_868),
.B(n_859),
.C(n_968),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1049),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1101),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_1089),
.A2(n_921),
.B(n_922),
.C(n_844),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_977),
.A2(n_866),
.B1(n_935),
.B2(n_932),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1115),
.B(n_930),
.C(n_952),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1025),
.B(n_862),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1113),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1062),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1068),
.B(n_936),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1090),
.Y(n_1245)
);

BUFx4f_ASAP7_75t_L g1246 ( 
.A(n_991),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1090),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1079),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1087),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1084),
.A2(n_806),
.B1(n_817),
.B2(n_804),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1107),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1107),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1084),
.A2(n_806),
.B1(n_817),
.B2(n_818),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1045),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1001),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1093),
.A2(n_931),
.B1(n_926),
.B2(n_945),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1107),
.Y(n_1257)
);

AOI222xp33_ASAP7_75t_L g1258 ( 
.A1(n_1092),
.A2(n_926),
.B1(n_931),
.B2(n_251),
.C1(n_250),
.C2(n_216),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1082),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1121),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1114),
.A2(n_952),
.B1(n_945),
.B2(n_844),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1121),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_972),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_972),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1083),
.B(n_1088),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_991),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1002),
.B(n_878),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1020),
.A2(n_960),
.B1(n_878),
.B2(n_873),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1094),
.B(n_960),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1108),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_976),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1102),
.A2(n_312),
.B1(n_873),
.B2(n_245),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_1095),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_994),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_976),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1097),
.A2(n_877),
.B(n_231),
.C(n_230),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1162),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_L g1279 ( 
.A1(n_1151),
.A2(n_1089),
.B(n_1123),
.C(n_1119),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1140),
.A2(n_1020),
.B1(n_1102),
.B2(n_1013),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1192),
.A2(n_1099),
.B(n_1014),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1217),
.A2(n_1108),
.B1(n_1102),
.B2(n_1119),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1059),
.B(n_1099),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1195),
.A2(n_1071),
.B(n_1072),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1254),
.B(n_1118),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_R g1286 ( 
.A(n_1164),
.B(n_1085),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1129),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1164),
.B(n_1005),
.Y(n_1288)
);

BUFx8_ASAP7_75t_SL g1289 ( 
.A(n_1154),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1254),
.B(n_1049),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1201),
.B(n_1109),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1201),
.B(n_994),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1255),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1133),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1137),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1166),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1195),
.A2(n_1072),
.B(n_1071),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1138),
.A2(n_1014),
.B(n_1082),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1125),
.B(n_1028),
.Y(n_1299)
);

CKINVDCx8_ASAP7_75t_R g1300 ( 
.A(n_1148),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1140),
.A2(n_1074),
.B1(n_1030),
.B2(n_1029),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1271),
.A2(n_1123),
.B(n_1117),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_1152),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1139),
.B(n_1080),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1147),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_1177),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1192),
.A2(n_1117),
.B(n_1116),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1259),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1221),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1135),
.B(n_1095),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1142),
.A2(n_1183),
.B(n_1224),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1150),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1156),
.A2(n_1116),
.B(n_1111),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1142),
.A2(n_1224),
.B(n_1183),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1172),
.B(n_1050),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1204),
.A2(n_1111),
.B(n_1050),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1130),
.Y(n_1317)
);

NOR2x1_ASAP7_75t_R g1318 ( 
.A(n_1155),
.B(n_1031),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1234),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1259),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1132),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1212),
.B(n_1244),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1139),
.B(n_1067),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1199),
.B(n_1110),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1223),
.B(n_1110),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1216),
.B(n_38),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1131),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1126),
.B(n_990),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_SL g1329 ( 
.A1(n_1215),
.A2(n_1032),
.B(n_1039),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1134),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1146),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1269),
.A2(n_1238),
.B(n_1250),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1226),
.A2(n_979),
.B1(n_998),
.B2(n_1124),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1219),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1139),
.B(n_1086),
.Y(n_1335)
);

BUFx2_ASAP7_75t_R g1336 ( 
.A(n_1179),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1139),
.B(n_1035),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1144),
.B(n_1106),
.Y(n_1338)
);

BUFx4_ASAP7_75t_SL g1339 ( 
.A(n_1187),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1238),
.A2(n_1032),
.B(n_1106),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1223),
.B(n_1034),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1203),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1208),
.A2(n_1034),
.B1(n_979),
.B2(n_1006),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1193),
.A2(n_1112),
.B(n_258),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1250),
.A2(n_312),
.B(n_226),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1269),
.A2(n_410),
.B(n_55),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1144),
.B(n_45),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1159),
.A2(n_224),
.B1(n_277),
.B2(n_272),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1184),
.B(n_268),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1141),
.Y(n_1350)
);

OAI222xp33_ASAP7_75t_L g1351 ( 
.A1(n_1191),
.A2(n_1136),
.B1(n_1145),
.B2(n_1182),
.C1(n_1169),
.C2(n_1213),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1157),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1174),
.B(n_267),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1159),
.A2(n_1230),
.B(n_1240),
.C(n_1215),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1236),
.A2(n_220),
.B(n_215),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1153),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1258),
.A2(n_212),
.B1(n_205),
.B2(n_410),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1178),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1261),
.A2(n_410),
.B(n_66),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1190),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1230),
.A2(n_410),
.B1(n_78),
.B2(n_79),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1130),
.B(n_410),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1130),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1198),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1227),
.B(n_61),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1219),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1163),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1167),
.Y(n_1368)
);

AOI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1258),
.A2(n_410),
.B(n_88),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1274),
.B(n_410),
.C(n_92),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1194),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1253),
.A2(n_1169),
.A3(n_1218),
.B(n_1277),
.Y(n_1372)
);

OAI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1227),
.A2(n_81),
.B1(n_105),
.B2(n_106),
.C(n_120),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1236),
.A2(n_124),
.B(n_129),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1136),
.B(n_155),
.Y(n_1375)
);

INVx4_ASAP7_75t_SL g1376 ( 
.A(n_1203),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1145),
.B(n_131),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1168),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1266),
.B(n_135),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1170),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1191),
.A2(n_138),
.B(n_139),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1200),
.A2(n_1253),
.B(n_1182),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1211),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1256),
.A2(n_142),
.B(n_147),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1237),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1231),
.B(n_1274),
.Y(n_1386)
);

AOI222xp33_ASAP7_75t_L g1387 ( 
.A1(n_1175),
.A2(n_1248),
.B1(n_1185),
.B2(n_1181),
.C1(n_1225),
.C2(n_1246),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1268),
.A2(n_1128),
.B(n_1127),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1214),
.B(n_1241),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1232),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1242),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1180),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1160),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1270),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1200),
.A2(n_1196),
.B(n_1235),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1127),
.A2(n_1158),
.B(n_1256),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1239),
.A2(n_1218),
.B(n_1213),
.C(n_1273),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1214),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1275),
.B(n_1206),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1203),
.A2(n_1143),
.B1(n_1246),
.B2(n_1267),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1272),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1267),
.B(n_1275),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1267),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1228),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1251),
.B(n_1263),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1239),
.A2(n_1205),
.B(n_1220),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1262),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1247),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1176),
.B(n_1188),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1276),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1158),
.A2(n_1233),
.B(n_1245),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1273),
.A2(n_1203),
.B1(n_1209),
.B2(n_1188),
.Y(n_1414)
);

OR2x6_ASAP7_75t_SL g1415 ( 
.A(n_1203),
.B(n_1210),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1264),
.B(n_1265),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1189),
.B(n_1186),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1189),
.A2(n_1186),
.B(n_1209),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1197),
.A2(n_1260),
.B(n_1252),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1196),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1149),
.A2(n_1171),
.B(n_1252),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1197),
.A2(n_1260),
.B(n_1245),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1207),
.A2(n_1171),
.B(n_1149),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1310),
.B(n_1207),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_L g1425 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1308),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1322),
.B(n_1229),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1311),
.A2(n_1279),
.B(n_1332),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1320),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1373),
.A2(n_1210),
.B1(n_1149),
.B2(n_1222),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1289),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1296),
.B(n_1161),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1309),
.B(n_1161),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1380),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1386),
.B(n_1161),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_L g1436 ( 
.A(n_1301),
.B(n_1165),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1357),
.A2(n_1369),
.B1(n_1387),
.B2(n_1408),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1376),
.B(n_1263),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1365),
.A2(n_1222),
.B(n_1251),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1406),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1357),
.A2(n_1210),
.B1(n_1247),
.B2(n_1202),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1280),
.A2(n_1348),
.B1(n_1398),
.B2(n_1361),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1395),
.B(n_1165),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1291),
.A2(n_1165),
.B(n_1173),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_SL g1445 ( 
.A(n_1336),
.B(n_1173),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1308),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1303),
.A2(n_1247),
.B1(n_1202),
.B2(n_1229),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1381),
.A2(n_1173),
.B1(n_1202),
.B2(n_1229),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1408),
.A2(n_1257),
.B1(n_1280),
.B2(n_1333),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1390),
.B(n_1257),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1320),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1386),
.B(n_1257),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1321),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1409),
.B(n_1403),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1376),
.B(n_1411),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1327),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1279),
.A2(n_1345),
.B(n_1348),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_SL g1459 ( 
.A(n_1282),
.B(n_1393),
.C(n_1406),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1284),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1380),
.B(n_1290),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1408),
.A2(n_1382),
.B1(n_1381),
.B2(n_1355),
.Y(n_1462)
);

INVx4_ASAP7_75t_SL g1463 ( 
.A(n_1334),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1398),
.A2(n_1354),
.A3(n_1345),
.B(n_1343),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1331),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1302),
.A2(n_1354),
.B1(n_1351),
.B2(n_1316),
.C(n_1373),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1326),
.B(n_1324),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1300),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1399),
.B(n_1287),
.Y(n_1470)
);

AND2x2_ASAP7_75t_SL g1471 ( 
.A(n_1342),
.B(n_1381),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1292),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1361),
.A2(n_1365),
.B1(n_1328),
.B2(n_1350),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1328),
.A2(n_1299),
.B1(n_1303),
.B2(n_1414),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1306),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1294),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1295),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1342),
.B(n_1366),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1382),
.A2(n_1355),
.B1(n_1384),
.B2(n_1344),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1305),
.B(n_1312),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1356),
.B(n_1367),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1355),
.A2(n_1384),
.B1(n_1344),
.B2(n_1360),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1339),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1400),
.B(n_1368),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1342),
.B(n_1291),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1378),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1292),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1389),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1391),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1342),
.B(n_1347),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1400),
.B(n_1285),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1376),
.B(n_1411),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1397),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1293),
.B(n_1286),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1341),
.B(n_1416),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1351),
.A2(n_1349),
.B1(n_1375),
.B2(n_1377),
.C(n_1307),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1392),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1319),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1278),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1346),
.A2(n_1283),
.B(n_1298),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1307),
.A2(n_1353),
.B1(n_1379),
.B2(n_1394),
.C(n_1420),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1293),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1317),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1412),
.B(n_1417),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1414),
.A2(n_1415),
.B1(n_1278),
.B2(n_1384),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1338),
.B(n_1404),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1352),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1358),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1421),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1286),
.A2(n_1347),
.B1(n_1288),
.B2(n_1385),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1315),
.B(n_1383),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1359),
.A2(n_1340),
.B(n_1413),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1314),
.A2(n_1288),
.B(n_1313),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_R g1516 ( 
.A(n_1364),
.B(n_1371),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1418),
.B(n_1401),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1338),
.B(n_1401),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1405),
.A2(n_1315),
.B1(n_1410),
.B2(n_1419),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1313),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1315),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1317),
.B(n_1363),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1363),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1420),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1289),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1314),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1339),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1344),
.A2(n_1329),
.B1(n_1281),
.B2(n_1396),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1422),
.B(n_1421),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1423),
.B(n_1407),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1372),
.B(n_1318),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1336),
.A2(n_1402),
.B1(n_1370),
.B2(n_1314),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1304),
.B(n_1323),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_SL g1534 ( 
.A(n_1402),
.B(n_1304),
.C(n_1323),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_R g1535 ( 
.A(n_1374),
.B(n_1388),
.Y(n_1535)
);

AOI221xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1372),
.A2(n_1396),
.B1(n_1374),
.B2(n_1281),
.C(n_1335),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1372),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1374),
.A2(n_1335),
.B(n_1337),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_SL g1539 ( 
.A(n_1337),
.B(n_1372),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1362),
.A2(n_400),
.B1(n_408),
.B2(n_790),
.C(n_724),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1362),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1339),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1376),
.B(n_1411),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1310),
.B(n_1395),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1442),
.A2(n_1540),
.B1(n_1437),
.B2(n_1467),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1524),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1524),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1517),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1498),
.A2(n_1474),
.B1(n_1475),
.B2(n_1449),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_SL g1550 ( 
.A(n_1431),
.B(n_1527),
.C(n_1516),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_R g1551 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1500),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1457),
.A2(n_1503),
.B(n_1512),
.C(n_1532),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_SL g1554 ( 
.A(n_1469),
.B(n_1484),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1468),
.B(n_1485),
.Y(n_1555)
);

NAND2xp33_ASAP7_75t_SL g1556 ( 
.A(n_1542),
.B(n_1469),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1529),
.B(n_1489),
.Y(n_1557)
);

OAI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1537),
.A2(n_1480),
.B(n_1459),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1489),
.B(n_1433),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1429),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1453),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1469),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1451),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1462),
.A2(n_1471),
.B1(n_1507),
.B2(n_1448),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1432),
.B(n_1427),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_R g1566 ( 
.A(n_1534),
.B(n_1445),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1435),
.B(n_1452),
.Y(n_1567)
);

INVxp33_ASAP7_75t_SL g1568 ( 
.A(n_1525),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_SL g1569 ( 
.A1(n_1444),
.A2(n_1482),
.B(n_1481),
.Y(n_1569)
);

AND2x4_ASAP7_75t_SL g1570 ( 
.A(n_1501),
.B(n_1453),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1536),
.A2(n_1515),
.B(n_1502),
.Y(n_1571)
);

NAND2xp33_ASAP7_75t_SL g1572 ( 
.A(n_1447),
.B(n_1453),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1472),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_R g1574 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1472),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1454),
.B(n_1497),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1490),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1520),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1461),
.B(n_1492),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1476),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1506),
.B(n_1495),
.Y(n_1581)
);

AND2x4_ASAP7_75t_SL g1582 ( 
.A(n_1473),
.B(n_1488),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1430),
.A2(n_1440),
.B1(n_1441),
.B2(n_1531),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1530),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_SL g1585 ( 
.A(n_1522),
.B(n_1434),
.C(n_1424),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_R g1586 ( 
.A(n_1491),
.B(n_1455),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1438),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1470),
.B(n_1477),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1476),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1425),
.A2(n_1504),
.B1(n_1463),
.B2(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1478),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_R g1592 ( 
.A(n_1455),
.B(n_1493),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1487),
.B(n_1450),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1439),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1499),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1483),
.A2(n_1537),
.B1(n_1544),
.B2(n_1510),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1463),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1517),
.B(n_1538),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1530),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1426),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1426),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1504),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1473),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1438),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1505),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1486),
.B(n_1543),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1508),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1446),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1479),
.A2(n_1518),
.B1(n_1428),
.B2(n_1523),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_R g1611 ( 
.A(n_1473),
.B(n_1488),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1460),
.B(n_1465),
.C(n_1526),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_R g1613 ( 
.A(n_1488),
.B(n_1523),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1505),
.B(n_1521),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1494),
.B(n_1539),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1526),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1509),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1533),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_R g1619 ( 
.A(n_1493),
.B(n_1543),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1571),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1585),
.B(n_1594),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1616),
.B(n_1428),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1616),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1571),
.B(n_1460),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1546),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.B(n_1465),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1612),
.B(n_1514),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1612),
.B(n_1528),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1546),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1547),
.Y(n_1631)
);

INVx2_ASAP7_75t_R g1632 ( 
.A(n_1615),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1578),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1600),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1547),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1555),
.B(n_1464),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1609),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1569),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1584),
.B(n_1464),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1577),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1584),
.B(n_1464),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1595),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1560),
.B(n_1511),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1591),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1563),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1588),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1599),
.B(n_1511),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1608),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1579),
.B(n_1519),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1557),
.B(n_1513),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1598),
.B(n_1533),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1607),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1598),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1598),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1576),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1557),
.B(n_1456),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1581),
.B(n_1458),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1558),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1596),
.B(n_1466),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1548),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1621),
.A2(n_1545),
.B(n_1549),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1621),
.B(n_1553),
.C(n_1545),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1660),
.B(n_1559),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1660),
.B(n_1565),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1567),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1614),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1663),
.A2(n_1566),
.B1(n_1574),
.B2(n_1583),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1624),
.A2(n_1596),
.B(n_1564),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1561),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1663),
.A2(n_1549),
.B1(n_1564),
.B2(n_1606),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1640),
.A2(n_1606),
.B(n_1548),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1666),
.B(n_1572),
.C(n_1556),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1666),
.A2(n_1606),
.B1(n_1590),
.B2(n_1548),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1574),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1637),
.B(n_1568),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1666),
.A2(n_1605),
.B(n_1619),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1647),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1624),
.Y(n_1685)
);

AND2x2_ASAP7_75t_SL g1686 ( 
.A(n_1629),
.B(n_1570),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1624),
.A2(n_1603),
.B(n_1602),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1649),
.B(n_1587),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1649),
.B(n_1587),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1648),
.B(n_1587),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1647),
.B(n_1587),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1628),
.A2(n_1604),
.B(n_1618),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1604),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1629),
.B(n_1620),
.C(n_1640),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1653),
.B(n_1618),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1629),
.B(n_1620),
.C(n_1640),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1640),
.B(n_1575),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1654),
.A2(n_1619),
.B1(n_1592),
.B2(n_1586),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1637),
.A2(n_1573),
.B1(n_1589),
.B2(n_1580),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1628),
.A2(n_1622),
.B(n_1620),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1554),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1626),
.B(n_1552),
.C(n_1592),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1637),
.A2(n_1562),
.B1(n_1550),
.B2(n_1566),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1620),
.B(n_1550),
.C(n_1586),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1620),
.B(n_1551),
.C(n_1611),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1657),
.B(n_1582),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1684),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1687),
.Y(n_1712)
);

INVxp33_ASAP7_75t_L g1713 ( 
.A(n_1682),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1685),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1685),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1637),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1632),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1670),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1706),
.B(n_1643),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1687),
.B(n_1632),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1687),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1670),
.B(n_1631),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1697),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1674),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1674),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1686),
.B(n_1646),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1675),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1623),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1690),
.B(n_1672),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1667),
.B(n_1631),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1695),
.B(n_1643),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1680),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1708),
.B(n_1643),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1671),
.B(n_1630),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1669),
.B(n_1630),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1669),
.B(n_1626),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1672),
.B(n_1623),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1688),
.Y(n_1739)
);

AND2x4_ASAP7_75t_SL g1740 ( 
.A(n_1701),
.B(n_1655),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1692),
.B(n_1623),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1636),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_SL g1743 ( 
.A(n_1686),
.B(n_1665),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1636),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1699),
.B(n_1622),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1689),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1692),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1694),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1724),
.A2(n_1668),
.B1(n_1676),
.B2(n_1673),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1731),
.B(n_1646),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1742),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1711),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1714),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1718),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1713),
.B(n_1703),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1732),
.B(n_1709),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1730),
.B(n_1704),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1714),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1718),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1735),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1723),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1735),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1722),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1716),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1740),
.B(n_1701),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1736),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1723),
.B(n_1622),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1737),
.Y(n_1771)
);

NAND2x1_ASAP7_75t_L g1772 ( 
.A(n_1712),
.B(n_1696),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1651),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1726),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1715),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1738),
.B(n_1696),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.B(n_1633),
.Y(n_1777)
);

NAND2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1712),
.B(n_1656),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1628),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.B(n_1633),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1729),
.B(n_1705),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1729),
.B(n_1683),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1715),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1733),
.B(n_1651),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1747),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1744),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1747),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1712),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1748),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1719),
.B(n_1691),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1762),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1740),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1678),
.Y(n_1795)
);

OAI33xp33_ASAP7_75t_L g1796 ( 
.A1(n_1752),
.A2(n_1727),
.A3(n_1725),
.B1(n_1724),
.B2(n_1745),
.B3(n_1748),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_L g1797 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1797)
);

NAND4xp75_ASAP7_75t_SL g1798 ( 
.A(n_1782),
.B(n_1717),
.C(n_1720),
.D(n_1741),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1768),
.B(n_1741),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1781),
.B(n_1719),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1786),
.B(n_1725),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1753),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1750),
.A2(n_1727),
.B(n_1721),
.C(n_1732),
.Y(n_1804)
);

OAI32xp33_ASAP7_75t_L g1805 ( 
.A1(n_1752),
.A2(n_1721),
.A3(n_1720),
.B1(n_1707),
.B2(n_1654),
.Y(n_1805)
);

AO22x1_ASAP7_75t_L g1806 ( 
.A1(n_1788),
.A2(n_1721),
.B1(n_1734),
.B2(n_1719),
.Y(n_1806)
);

OAI33xp33_ASAP7_75t_L g1807 ( 
.A1(n_1752),
.A2(n_1645),
.A3(n_1679),
.B1(n_1702),
.B2(n_1625),
.B3(n_1633),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1753),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1761),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1751),
.B(n_1746),
.Y(n_1811)
);

OAI32xp33_ASAP7_75t_L g1812 ( 
.A1(n_1766),
.A2(n_1739),
.A3(n_1710),
.B1(n_1633),
.B2(n_1625),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1785),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1765),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1761),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1765),
.Y(n_1817)
);

OR2x6_ASAP7_75t_L g1818 ( 
.A(n_1778),
.B(n_1677),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1781),
.B(n_1732),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1763),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1734),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1766),
.A2(n_1732),
.B(n_1693),
.C(n_1620),
.Y(n_1823)
);

OAI32xp33_ASAP7_75t_L g1824 ( 
.A1(n_1766),
.A2(n_1778),
.A3(n_1782),
.B1(n_1758),
.B2(n_1779),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1763),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1799),
.B(n_1758),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1795),
.B(n_1769),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1822),
.B(n_1771),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1791),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1811),
.B(n_1764),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1797),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1793),
.B(n_1769),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1800),
.B(n_1771),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1804),
.A2(n_1772),
.B(n_1757),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1815),
.B(n_1764),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1817),
.B(n_1809),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1821),
.B(n_1789),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1794),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1802),
.B(n_1760),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1810),
.B(n_1789),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1816),
.B(n_1755),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1804),
.A2(n_1757),
.B(n_1772),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1794),
.B(n_1776),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1819),
.A2(n_1757),
.B1(n_1778),
.B2(n_1790),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1802),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1820),
.B(n_1760),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1801),
.B(n_1776),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1798),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1825),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1835),
.A2(n_1805),
.B(n_1824),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_L g1852 ( 
.A(n_1827),
.B(n_1796),
.C(n_1806),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1846),
.A2(n_1807),
.B1(n_1812),
.B2(n_1823),
.C(n_1808),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1849),
.A2(n_1807),
.B1(n_1814),
.B2(n_1803),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1826),
.B(n_1813),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1828),
.B(n_1792),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1832),
.B(n_1818),
.Y(n_1857)
);

AOI222xp33_ASAP7_75t_L g1858 ( 
.A1(n_1843),
.A2(n_1779),
.B1(n_1620),
.B2(n_1787),
.C1(n_1785),
.C2(n_1770),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1841),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1842),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1844),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1838),
.A2(n_1798),
.B(n_1755),
.Y(n_1862)
);

AND2x2_ASAP7_75t_SL g1863 ( 
.A(n_1832),
.B(n_1787),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1826),
.B(n_1784),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1847),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1839),
.A2(n_1818),
.B1(n_1777),
.B2(n_1780),
.Y(n_1866)
);

AOI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1831),
.A2(n_1818),
.B(n_1777),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1829),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1850),
.A2(n_1620),
.B1(n_1783),
.B2(n_1775),
.C(n_1754),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1831),
.A2(n_1783),
.B(n_1775),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1864),
.B(n_1828),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1856),
.Y(n_1872)
);

OAI32xp33_ASAP7_75t_L g1873 ( 
.A1(n_1852),
.A2(n_1845),
.A3(n_1840),
.B1(n_1830),
.B2(n_1833),
.Y(n_1873)
);

AOI21xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1851),
.A2(n_1834),
.B(n_1837),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1868),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1861),
.B(n_1848),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1848),
.Y(n_1877)
);

AOI221x1_ASAP7_75t_L g1878 ( 
.A1(n_1867),
.A2(n_1836),
.B1(n_1844),
.B2(n_1754),
.C(n_1759),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1855),
.B(n_1759),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1857),
.B(n_1780),
.Y(n_1880)
);

AOI32xp33_ASAP7_75t_L g1881 ( 
.A1(n_1853),
.A2(n_1627),
.A3(n_1641),
.B1(n_1625),
.B2(n_1658),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1874),
.A2(n_1854),
.B1(n_1862),
.B2(n_1866),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1877),
.A2(n_1854),
.B1(n_1858),
.B2(n_1857),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1871),
.A2(n_1862),
.B1(n_1859),
.B2(n_1860),
.Y(n_1884)
);

NOR3xp33_ASAP7_75t_L g1885 ( 
.A(n_1873),
.B(n_1865),
.C(n_1870),
.Y(n_1885)
);

OAI222xp33_ASAP7_75t_L g1886 ( 
.A1(n_1881),
.A2(n_1879),
.B1(n_1880),
.B2(n_1875),
.C1(n_1876),
.C2(n_1872),
.Y(n_1886)
);

AOI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1869),
.B(n_1627),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_SL g1888 ( 
.A(n_1878),
.B(n_1641),
.Y(n_1888)
);

O2A1O1Ixp5_ASAP7_75t_L g1889 ( 
.A1(n_1873),
.A2(n_1625),
.B(n_1627),
.C(n_1645),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1880),
.B(n_1641),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1884),
.Y(n_1891)
);

AO22x2_ASAP7_75t_L g1892 ( 
.A1(n_1882),
.A2(n_1659),
.B1(n_1658),
.B2(n_1665),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1886),
.A2(n_1645),
.B(n_1634),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1885),
.B(n_1639),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1891),
.B(n_1883),
.C(n_1888),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_L g1897 ( 
.A(n_1895),
.B(n_1887),
.C(n_1890),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1892),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_L g1899 ( 
.A1(n_1894),
.A2(n_1551),
.B(n_1650),
.Y(n_1899)
);

NAND4xp25_ASAP7_75t_SL g1900 ( 
.A(n_1893),
.B(n_1659),
.C(n_1658),
.D(n_1665),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1891),
.B(n_1655),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1896),
.B(n_1659),
.Y(n_1902)
);

NOR2x1_ASAP7_75t_L g1903 ( 
.A(n_1901),
.B(n_1898),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1899),
.B(n_1897),
.C(n_1900),
.Y(n_1904)
);

OAI322xp33_ASAP7_75t_L g1905 ( 
.A1(n_1896),
.A2(n_1634),
.A3(n_1635),
.B1(n_1639),
.B2(n_1664),
.C1(n_1659),
.C2(n_1658),
.Y(n_1905)
);

NAND4xp75_ASAP7_75t_L g1906 ( 
.A(n_1898),
.B(n_1650),
.C(n_1665),
.D(n_1655),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1903),
.B(n_1656),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1902),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1905),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1907),
.B(n_1904),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1910),
.Y(n_1911)
);

XOR2xp5_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1908),
.Y(n_1912)
);

XNOR2xp5_ASAP7_75t_L g1913 ( 
.A(n_1911),
.B(n_1909),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1912),
.B(n_1906),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1913),
.Y(n_1915)
);

OAI22x1_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1656),
.B1(n_1634),
.B2(n_1635),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1914),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1634),
.B1(n_1635),
.B2(n_1639),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1916),
.B1(n_1662),
.B2(n_1639),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1919),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1635),
.B1(n_1662),
.B2(n_1664),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1921),
.A2(n_1656),
.B(n_1650),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1656),
.B1(n_1642),
.B2(n_1644),
.Y(n_1923)
);

OAI31xp33_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1656),
.A3(n_1664),
.B(n_1661),
.Y(n_1924)
);


endmodule