module fake_jpeg_14633_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_182;
wire n_19;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_48),
.Y(n_78)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_22),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_23),
.B(n_38),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_58),
.Y(n_102)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_0),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_26),
.C(n_17),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_89),
.C(n_8),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_32),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_75),
.B(n_3),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_80),
.B1(n_82),
.B2(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_76),
.A2(n_96),
.B1(n_105),
.B2(n_104),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_27),
.B1(n_30),
.B2(n_37),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_16),
.B1(n_38),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_29),
.B1(n_36),
.B2(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_30),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_29),
.B(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_28),
.B1(n_36),
.B2(n_34),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_36),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_34),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_24),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_107),
.B(n_1),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_42),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_81),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_39),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_120),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_125),
.Y(n_163)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_132),
.B1(n_134),
.B2(n_83),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_7),
.Y(n_124)
);

XOR2x2_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_8),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_133),
.Y(n_155)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_70),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_79),
.Y(n_153)
);

OR2x2_ASAP7_75t_SL g131 ( 
.A(n_66),
.B(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_136),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_5),
.B1(n_13),
.B2(n_3),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_1),
.B(n_2),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_15),
.B1(n_99),
.B2(n_98),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_74),
.B(n_4),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_4),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_5),
.C(n_10),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_66),
.B(n_13),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_15),
.C(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_70),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_145),
.B(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_162),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_95),
.B1(n_81),
.B2(n_84),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_108),
.B1(n_126),
.B2(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_169),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_92),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_92),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_94),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_94),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_117),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_98),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_139),
.B(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_95),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_88),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_139),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_201),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_179),
.B1(n_117),
.B2(n_164),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_128),
.C(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_186),
.C(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_112),
.B1(n_124),
.B2(n_141),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_133),
.B(n_123),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_193),
.B(n_120),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_146),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_192),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_175),
.C(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_123),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_157),
.B(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_143),
.C(n_136),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_186),
.C(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_142),
.B1(n_131),
.B2(n_130),
.Y(n_198)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_159),
.B1(n_145),
.B2(n_166),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_215),
.B1(n_219),
.B2(n_200),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_161),
.C(n_166),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_214),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_180),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_151),
.B1(n_161),
.B2(n_152),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_199),
.B1(n_192),
.B2(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_158),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_158),
.C(n_163),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_163),
.C(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_220),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_156),
.B1(n_144),
.B2(n_173),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_186),
.C(n_191),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_165),
.C(n_147),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_176),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.C(n_235),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_232),
.B1(n_208),
.B2(n_217),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_183),
.B(n_198),
.C(n_184),
.D(n_180),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_216),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_179),
.B1(n_195),
.B2(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_189),
.C(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_210),
.C(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_235),
.C(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_204),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_209),
.B1(n_202),
.B2(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_196),
.B1(n_182),
.B2(n_154),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_202),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_222),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_233),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_241),
.A2(n_231),
.B1(n_205),
.B2(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_254),
.B(n_240),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_257),
.A3(n_251),
.B1(n_248),
.B2(n_237),
.C1(n_73),
.C2(n_88),
.Y(n_259)
);

AOI31xp33_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_253),
.A3(n_249),
.B(n_252),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_253),
.A2(n_240),
.B(n_182),
.C(n_147),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_258),
.C(n_73),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_237),
.C(n_165),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_111),
.C(n_135),
.Y(n_261)
);

XNOR2x2_ASAP7_75t_SL g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_264),
.Y(n_265)
);


endmodule