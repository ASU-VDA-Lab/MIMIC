module real_jpeg_16705_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_623, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_623;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_553;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_620;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_1),
.A2(n_84),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_1),
.A2(n_153),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_1),
.A2(n_153),
.B1(n_461),
.B2(n_464),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_1),
.A2(n_153),
.B1(n_472),
.B2(n_474),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_126),
.B1(n_196),
.B2(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_2),
.A2(n_126),
.B1(n_326),
.B2(n_335),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_2),
.A2(n_126),
.B1(n_319),
.B2(n_560),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_3),
.A2(n_129),
.B1(n_293),
.B2(n_297),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_3),
.A2(n_129),
.B1(n_438),
.B2(n_443),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_3),
.A2(n_125),
.B1(n_129),
.B2(n_494),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_4),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_4),
.Y(n_355)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_7),
.A2(n_40),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_7),
.A2(n_40),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_7),
.A2(n_40),
.B1(n_448),
.B2(n_450),
.Y(n_447)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_9),
.A2(n_72),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_9),
.A2(n_72),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_9),
.A2(n_72),
.B1(n_408),
.B2(n_413),
.Y(n_407)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_10),
.B(n_156),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g399 ( 
.A1(n_10),
.A2(n_48),
.A3(n_276),
.B1(n_400),
.B2(n_403),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_10),
.B(n_78),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_10),
.A2(n_102),
.B1(n_239),
.B2(n_493),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_10),
.A2(n_82),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_175),
.B1(n_177),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_11),
.A2(n_179),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_11),
.A2(n_179),
.B1(n_335),
.B2(n_567),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_11),
.A2(n_179),
.B1(n_597),
.B2(n_609),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_13),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_13),
.A2(n_166),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_13),
.A2(n_166),
.B1(n_551),
.B2(n_553),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_13),
.A2(n_83),
.B1(n_166),
.B2(n_597),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_14),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_14),
.A2(n_111),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_14),
.A2(n_111),
.B1(n_324),
.B2(n_327),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_14),
.A2(n_111),
.B1(n_544),
.B2(n_547),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_16),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_16),
.A2(n_234),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

OAI22x1_ASAP7_75t_SL g299 ( 
.A1(n_16),
.A2(n_234),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_16),
.A2(n_234),
.B1(n_319),
.B2(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_17),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_17),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_17),
.Y(n_237)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_17),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g131 ( 
.A(n_19),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_19),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_19),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B(n_24),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_617),
.B(n_620),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_534),
.B(n_610),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_380),
.B(n_529),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_311),
.C(n_375),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_259),
.B(n_284),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_30),
.B(n_259),
.C(n_531),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_157),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_31),
.B(n_158),
.C(n_227),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_79),
.C(n_127),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_33),
.B(n_127),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_47),
.B1(n_69),
.B2(n_77),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_35),
.A2(n_78),
.B1(n_266),
.B2(n_271),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_44),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_46),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_46),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_47),
.A2(n_69),
.B1(n_77),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_47),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_47),
.A2(n_77),
.B1(n_253),
.B2(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_47),
.A2(n_77),
.B1(n_292),
.B2(n_511),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_47),
.A2(n_77),
.B1(n_334),
.B2(n_550),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_47),
.A2(n_77),
.B1(n_550),
.B2(n_566),
.Y(n_565)
);

AO21x2_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_54),
.B(n_62),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_63),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_63),
.Y(n_233)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_67),
.Y(n_345)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_67),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_68),
.Y(n_278)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_78),
.A2(n_266),
.B1(n_271),
.B2(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_78),
.A2(n_271),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_78),
.A2(n_271),
.B(n_593),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_79),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_101),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_80),
.B(n_101),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_SL g273 ( 
.A1(n_81),
.A2(n_82),
.B(n_130),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_82),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_82),
.B(n_425),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g435 ( 
.A1(n_82),
.A2(n_424),
.B(n_436),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_82),
.B(n_306),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_82),
.B(n_183),
.Y(n_499)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_86),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_86),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_94),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_136),
.B(n_140),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_100),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_108),
.B1(n_117),
.B2(n_119),
.Y(n_101)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_102),
.A2(n_119),
.B1(n_162),
.B2(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_102),
.A2(n_174),
.B(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_102),
.A2(n_172),
.B1(n_447),
.B2(n_455),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_102),
.A2(n_471),
.B1(n_493),
.B2(n_497),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_106),
.Y(n_422)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_107),
.Y(n_301)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_107),
.Y(n_412)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22x1_ASAP7_75t_SL g298 ( 
.A1(n_109),
.A2(n_160),
.B1(n_299),
.B2(n_305),
.Y(n_298)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_114),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_115),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_122),
.Y(n_413)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_123),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_123),
.Y(n_449)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_135),
.B1(n_151),
.B2(n_156),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_128),
.A2(n_135),
.B1(n_156),
.B2(n_273),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_135),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_135),
.A2(n_156),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_135),
.A2(n_156),
.B(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g316 ( 
.A1(n_140),
.A2(n_245),
.B1(n_247),
.B2(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_140),
.A2(n_245),
.B1(n_317),
.B2(n_362),
.Y(n_361)
);

AOI22x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_146),
.B2(n_149),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_147),
.Y(n_328)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_148),
.Y(n_570)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22x1_ASAP7_75t_SL g244 ( 
.A1(n_152),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_227),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_180),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_159),
.A2(n_181),
.B(n_206),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_171),
.B2(n_173),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_160),
.A2(n_240),
.B1(n_299),
.B2(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_160),
.A2(n_470),
.B1(n_477),
.B2(n_478),
.Y(n_469)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_206),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_194),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_182),
.A2(n_207),
.B1(n_275),
.B2(n_283),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_182),
.A2(n_207),
.B1(n_339),
.B2(n_346),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_182),
.A2(n_207),
.B1(n_435),
.B2(n_437),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_182),
.A2(n_207),
.B1(n_437),
.B2(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_182),
.A2(n_207),
.B1(n_390),
.B2(n_460),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g540 ( 
.A1(n_182),
.A2(n_207),
.B(n_346),
.Y(n_540)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_220),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_183),
.A2(n_195),
.B1(n_230),
.B2(n_340),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_183),
.A2(n_230),
.B1(n_389),
.B2(n_396),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_191),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_191),
.Y(n_473)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_191),
.Y(n_490)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_193),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_219),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_216),
.B2(n_218),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_212),
.Y(n_348)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_212),
.Y(n_395)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_216),
.Y(n_423)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_222),
.Y(n_349)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_243),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_228),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

XOR2x2_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_238),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_231),
.Y(n_283)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_236),
.Y(n_465)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_239),
.Y(n_477)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_244),
.B(n_252),
.C(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_245),
.A2(n_246),
.B1(n_362),
.B2(n_543),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_245),
.A2(n_246),
.B1(n_595),
.B2(n_596),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_245),
.A2(n_246),
.B1(n_596),
.B2(n_608),
.Y(n_607)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_257),
.Y(n_554)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_258),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_264),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_261),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_264),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.C(n_274),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_274),
.Y(n_287)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_275),
.Y(n_396)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_281),
.Y(n_404)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_308),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_285),
.B(n_308),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.C(n_289),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_286),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_288),
.B(n_289),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.C(n_307),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_290),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_298),
.B(n_307),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_300),
.Y(n_494)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

A2O1A1O1Ixp25_ASAP7_75t_L g529 ( 
.A1(n_311),
.A2(n_375),
.B(n_530),
.C(n_532),
.D(n_533),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_366),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_312),
.B(n_366),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_329),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_313),
.B(n_584),
.C(n_585),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.C(n_322),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_314),
.B(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_322),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_318),
.Y(n_321)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_320),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_326),
.Y(n_512)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_326),
.Y(n_552)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_351),
.Y(n_329)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_330),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_338),
.B(n_350),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_338),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_350),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_350),
.A2(n_576),
.B1(n_578),
.B2(n_588),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_351),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_357),
.B1(n_358),
.B2(n_365),
.Y(n_351)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_352),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_353),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_353),
.A2(n_356),
.B1(n_359),
.B2(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx12f_ASAP7_75t_L g498 ( 
.A(n_355),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_359),
.A2(n_365),
.B1(n_580),
.B2(n_623),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_360),
.Y(n_581)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.C(n_372),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_368),
.B1(n_370),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_370),
.Y(n_378)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_376),
.B(n_379),
.Y(n_532)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_414),
.B(n_528),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_382),
.B(n_384),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.C(n_397),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_385),
.A2(n_386),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_388),
.A2(n_397),
.B1(n_398),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_405),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_399),
.A2(n_405),
.B1(n_406),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_521),
.B(n_527),
.Y(n_414)
);

AOI21x1_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_503),
.B(n_520),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_467),
.B(n_502),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_445),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_418),
.B(n_445),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_433),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_419),
.A2(n_433),
.B1(n_434),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

OAI32xp33_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_422),
.A3(n_423),
.B1(n_424),
.B2(n_426),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_456),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_458),
.C(n_466),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_459),
.B2(n_466),
.Y(n_456)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_481),
.B(n_501),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_479),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_479),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_495),
.B(n_500),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_492),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_491),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_499),
.Y(n_500)
);

INVx6_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_505),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_509),
.C(n_519),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_518),
.B2(n_519),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_526),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_526),
.Y(n_527)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_589),
.C(n_605),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_582),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_537),
.A2(n_613),
.B(n_614),
.Y(n_612)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_575),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_538),
.B(n_575),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_555),
.Y(n_538)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_539),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.C(n_549),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_540),
.A2(n_565),
.B1(n_571),
.B2(n_572),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_540),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_549),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_540),
.B(n_557),
.C(n_572),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_556),
.B1(n_573),
.B2(n_574),
.Y(n_555)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_543),
.Y(n_558)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_546),
.Y(n_563)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_546),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_573),
.C(n_604),
.Y(n_603)
);

XNOR2x1_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_564),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_559),
.Y(n_595)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_565),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_578),
.C(n_579),
.Y(n_575)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_586),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_583),
.B(n_586),
.Y(n_613)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

A2O1A1O1Ixp25_ASAP7_75t_L g611 ( 
.A1(n_590),
.A2(n_606),
.B(n_612),
.C(n_615),
.D(n_616),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_603),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_607),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_591),
.B(n_603),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_607),
.Y(n_616)
);

FAx1_ASAP7_75t_SL g591 ( 
.A(n_592),
.B(n_594),
.CI(n_602),
.CON(n_591),
.SN(n_591)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_598),
.Y(n_609)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_618),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_607),
.B(n_618),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_608),
.Y(n_619)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_621),
.Y(n_620)
);


endmodule