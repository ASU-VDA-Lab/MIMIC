module fake_jpeg_5695_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_29),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_63)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_16),
.Y(n_76)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_28),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_16),
.B1(n_33),
.B2(n_38),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_38),
.B1(n_22),
.B2(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_26),
.B1(n_23),
.B2(n_32),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_19),
.B1(n_42),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_80),
.B1(n_30),
.B2(n_17),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_16),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_82),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_19),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_37),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_50),
.B1(n_61),
.B2(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_87),
.C(n_12),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_42),
.C(n_33),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_67),
.C(n_80),
.Y(n_107)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_24),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_47),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_97),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_52),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_50),
.B1(n_52),
.B2(n_49),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_95),
.B(n_108),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_43),
.B(n_42),
.C(n_30),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_75),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_49),
.B1(n_42),
.B2(n_43),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_86),
.B1(n_79),
.B2(n_83),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_83),
.B1(n_86),
.B2(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_85),
.C(n_82),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_49),
.B1(n_25),
.B2(n_29),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_25),
.A3(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_95),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_63),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_120),
.C(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_85),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_66),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_130),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_91),
.B1(n_108),
.B2(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_87),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_74),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_74),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_133),
.CI(n_123),
.CON(n_137),
.SN(n_137)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_64),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_64),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_78),
.B(n_27),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_91),
.B(n_98),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_147),
.B(n_157),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_103),
.B1(n_105),
.B2(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_143),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_104),
.B1(n_98),
.B2(n_68),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_68),
.B1(n_35),
.B2(n_58),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_132),
.B(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_126),
.B1(n_130),
.B2(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_125),
.C(n_112),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_178),
.C(n_181),
.Y(n_192)
);

NAND4xp25_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_160),
.C(n_149),
.D(n_137),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_58),
.C(n_17),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_93),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_0),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_175),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_93),
.B(n_58),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_180),
.B1(n_184),
.B2(n_153),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_183),
.B1(n_162),
.B2(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_58),
.C(n_35),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_35),
.B1(n_20),
.B2(n_17),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_35),
.C(n_20),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_9),
.B(n_15),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_148),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_20),
.B1(n_17),
.B2(n_2),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_143),
.B1(n_147),
.B2(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_199),
.B1(n_201),
.B2(n_175),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_202),
.C(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_144),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_139),
.B1(n_162),
.B2(n_142),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_149),
.B1(n_139),
.B2(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_198),
.B1(n_184),
.B2(n_180),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_160),
.A3(n_140),
.B1(n_20),
.B2(n_10),
.C1(n_5),
.C2(n_6),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_140),
.B1(n_1),
.B2(n_3),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_170),
.B1(n_163),
.B2(n_176),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_198),
.B(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_1),
.C(n_4),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_173),
.B1(n_166),
.B2(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_185),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_194),
.B(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_214),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_186),
.B1(n_176),
.B2(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.C(n_192),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_203),
.B1(n_202),
.B2(n_4),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_178),
.C(n_183),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_191),
.B(n_195),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_225),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_189),
.C(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_226),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_5),
.C(n_7),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_206),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_228)
);

AOI221xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_205),
.B1(n_216),
.B2(n_206),
.C(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_232),
.C(n_221),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_204),
.B(n_214),
.C(n_212),
.D(n_208),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_13),
.B(n_14),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_213),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_13),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_223),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_242),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_8),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_237),
.B1(n_236),
.B2(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_248),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g248 ( 
.A(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_233),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_14),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_247),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_15),
.Y(n_256)
);


endmodule