module fake_jpeg_11079_n_123 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_15),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_14),
.B1(n_16),
.B2(n_25),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_48),
.B1(n_35),
.B2(n_1),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_52),
.Y(n_61)
);

OR2x4_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_25),
.B1(n_13),
.B2(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_22),
.B1(n_48),
.B2(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_21),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_19),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_68),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_42),
.B(n_55),
.C(n_53),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_22),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_86),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_66),
.B1(n_60),
.B2(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_85),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_8),
.C(n_12),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_61),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_94),
.C(n_97),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_65),
.B1(n_70),
.B2(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_91),
.B1(n_69),
.B2(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_60),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_73),
.C(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_82),
.C(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_75),
.B(n_84),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_95),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_76),
.B1(n_71),
.B2(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_98),
.B1(n_105),
.B2(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_97),
.C(n_87),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_111),
.B(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_106),
.B1(n_109),
.B2(n_58),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_57),
.B1(n_7),
.B2(n_9),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_113),
.B(n_9),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_104),
.C(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_1),
.C(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_10),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_0),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_121),
.B(n_4),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_5),
.B(n_118),
.Y(n_123)
);


endmodule