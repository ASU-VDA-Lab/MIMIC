module fake_jpeg_6311_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_61),
.B1(n_68),
.B2(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_22),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_17),
.B(n_32),
.C(n_26),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_23),
.B1(n_19),
.B2(n_31),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_28),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_64),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_29),
.CI(n_28),
.CON(n_77),
.SN(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_29),
.B(n_17),
.C(n_32),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_34),
.B1(n_16),
.B2(n_26),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_58),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_45),
.B(n_50),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_106),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_39),
.B1(n_40),
.B2(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_39),
.B(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_47),
.B1(n_56),
.B2(n_23),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_62),
.B1(n_46),
.B2(n_18),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_62),
.B1(n_46),
.B2(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_83),
.B1(n_87),
.B2(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_92),
.B1(n_90),
.B2(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_83),
.B1(n_84),
.B2(n_91),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_31),
.B(n_27),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_69),
.C(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_127),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_69),
.C(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_69),
.C(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_132),
.Y(n_165)
);

AO21x2_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_111),
.B(n_105),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_112),
.B(n_33),
.Y(n_152)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_137),
.Y(n_169)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_79),
.C(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_16),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_94),
.B(n_95),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_20),
.B(n_33),
.Y(n_161)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_99),
.B1(n_108),
.B2(n_119),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_157),
.B(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_145),
.B1(n_123),
.B2(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_98),
.B1(n_118),
.B2(n_33),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_161),
.B1(n_170),
.B2(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR4xp25_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_10),
.C(n_11),
.D(n_9),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_33),
.B(n_20),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_33),
.B1(n_20),
.B2(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_171),
.B1(n_150),
.B2(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_186),
.B1(n_171),
.B2(n_148),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_122),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_181),
.C(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_120),
.C(n_143),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_142),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_189),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_149),
.A2(n_124),
.B1(n_132),
.B2(n_139),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_191),
.C(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_130),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_114),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_214),
.B(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_220),
.B1(n_147),
.B2(n_139),
.Y(n_233)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_211),
.B(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_172),
.A2(n_152),
.B1(n_161),
.B2(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_176),
.C(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.C(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_188),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_190),
.C(n_183),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_152),
.B(n_194),
.C(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_167),
.C(n_147),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_234),
.C(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_197),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_114),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_141),
.B1(n_101),
.B2(n_2),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_238),
.B1(n_205),
.B2(n_210),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_141),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_217),
.B1(n_10),
.B2(n_11),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_1),
.C(n_3),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_249),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_252),
.B1(n_254),
.B2(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_204),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_227),
.B1(n_239),
.B2(n_224),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_201),
.C(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.C(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_256),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_200),
.B1(n_198),
.B2(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_216),
.C(n_202),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_204),
.B(n_216),
.C(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_236),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_216),
.CI(n_4),
.CON(n_256),
.SN(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_264),
.C(n_247),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_250),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_221),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_254),
.CI(n_256),
.CON(n_274),
.SN(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_226),
.C(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_229),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_254),
.B(n_241),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_234),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_248),
.C(n_254),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_275),
.B(n_277),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_280),
.B(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_272),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_245),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_240),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_9),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_238),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_284),
.B(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_289),
.C(n_4),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_1),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_8),
.B(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_7),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_271),
.B(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_292),
.B(n_295),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_294),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_7),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_8),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_15),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_296),
.A2(n_13),
.B(n_14),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_8),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_14),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_13),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_302),
.B(n_299),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_300),
.C(n_15),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_15),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_5),
.C(n_296),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_5),
.B(n_296),
.Y(n_307)
);


endmodule