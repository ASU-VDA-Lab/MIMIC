module fake_jpeg_4960_n_15 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_15);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_15;

wire n_13;
wire n_11;
wire n_14;
wire n_12;
wire n_10;
wire n_8;
wire n_9;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_1),
.Y(n_7)
);

INVxp67_ASAP7_75t_SL g8 ( 
.A(n_2),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g9 ( 
.A1(n_6),
.A2(n_5),
.B1(n_1),
.B2(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_7),
.A2(n_4),
.B(n_11),
.Y(n_12)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_13),
.B(n_14),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_7),
.B1(n_11),
.B2(n_8),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_9),
.B1(n_7),
.B2(n_11),
.Y(n_14)
);


endmodule