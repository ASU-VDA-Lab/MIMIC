module fake_ibex_241_n_837 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_158, n_132, n_157, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_837);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_158;
input n_132;
input n_157;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_837;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_801;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_782;
wire n_616;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVxp33_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_51),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_62),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_55),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_19),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_86),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_45),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_15),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_116),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_63),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_33),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_79),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_108),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_103),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_72),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_71),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_5),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_3),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_25),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g221 ( 
.A(n_120),
.B(n_73),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_68),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_43),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_23),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_89),
.Y(n_233)
);

BUFx2_ASAP7_75t_SL g234 ( 
.A(n_10),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_82),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_119),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_88),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_6),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_96),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_99),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_115),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_93),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_94),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_85),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_58),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_92),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_83),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_158),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_69),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_80),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_66),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_163),
.Y(n_263)
);

AOI22x1_ASAP7_75t_SL g264 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_160),
.B(n_1),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_2),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_3),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_166),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_4),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_159),
.B(n_7),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_165),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_186),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_169),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_182),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_180),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_196),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_201),
.A2(n_70),
.B(n_152),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_159),
.B(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_168),
.B(n_9),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_181),
.B(n_10),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_170),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_202),
.A2(n_74),
.B(n_149),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_203),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_216),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_206),
.A2(n_67),
.B(n_148),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_230),
.A2(n_65),
.B(n_146),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_11),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_230),
.A2(n_75),
.B(n_144),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_196),
.B(n_30),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_173),
.B(n_13),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_14),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_212),
.B(n_16),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_77),
.B(n_142),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_241),
.A2(n_76),
.B(n_141),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_255),
.B(n_17),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

OAI22x1_ASAP7_75t_R g314 ( 
.A1(n_219),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_212),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_176),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_252),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_216),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_215),
.B(n_18),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_216),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_255),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_184),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_218),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_185),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_307),
.B(n_187),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_188),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

OR2x6_ASAP7_75t_L g336 ( 
.A(n_273),
.B(n_234),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_273),
.B(n_191),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_264),
.A2(n_189),
.B1(n_261),
.B2(n_224),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g345 ( 
.A1(n_264),
.A2(n_267),
.B1(n_327),
.B2(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_313),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_281),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_276),
.Y(n_356)
);

NOR2x1p5_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_229),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_269),
.B(n_192),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_275),
.A2(n_235),
.B1(n_253),
.B2(n_258),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_275),
.B(n_161),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_219),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_311),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_285),
.B(n_228),
.C(n_259),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_311),
.Y(n_371)
);

OR2x6_ASAP7_75t_L g372 ( 
.A(n_272),
.B(n_221),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_280),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_277),
.B(n_172),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_319),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_279),
.B(n_177),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_270),
.A2(n_178),
.B1(n_257),
.B2(n_210),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_279),
.B(n_194),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_289),
.B(n_179),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_289),
.B(n_195),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_291),
.B(n_207),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_306),
.B(n_211),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_296),
.Y(n_385)
);

NOR2x1p5_ASAP7_75t_L g386 ( 
.A(n_286),
.B(n_217),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_220),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_265),
.B(n_223),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_292),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_326),
.B(n_225),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_293),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_292),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

AND3x2_ASAP7_75t_L g395 ( 
.A(n_314),
.B(n_244),
.C(n_256),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_283),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_334),
.A2(n_302),
.B1(n_293),
.B2(n_288),
.Y(n_398)
);

OR2x6_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_338),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_210),
.B1(n_257),
.B2(n_178),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_347),
.B(n_299),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_328),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_162),
.B1(n_183),
.B2(n_249),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_322),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_329),
.A2(n_297),
.B(n_284),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_315),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_174),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_316),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_316),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_332),
.B(n_198),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_318),
.Y(n_412)
);

OR2x6_ASAP7_75t_L g413 ( 
.A(n_336),
.B(n_314),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_190),
.Y(n_415)
);

BUFx6f_ASAP7_75t_SL g416 ( 
.A(n_336),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_366),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_365),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_369),
.Y(n_421)
);

OR2x6_ASAP7_75t_L g422 ( 
.A(n_338),
.B(n_265),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_329),
.A2(n_295),
.B(n_284),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_356),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_331),
.A2(n_295),
.B(n_297),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_345),
.A2(n_231),
.B1(n_245),
.B2(n_232),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_371),
.B(n_204),
.Y(n_431)
);

BUFx12f_ASAP7_75t_SL g432 ( 
.A(n_372),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_348),
.B(n_214),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_345),
.A2(n_250),
.B1(n_240),
.B2(n_246),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_392),
.A2(n_290),
.B1(n_300),
.B2(n_308),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_193),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_366),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_345),
.A2(n_254),
.B1(n_199),
.B2(n_200),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_342),
.A2(n_290),
.B1(n_300),
.B2(n_308),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_362),
.B(n_197),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_290),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_362),
.B(n_205),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_237),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_382),
.B(n_248),
.Y(n_449)
);

BUFx5_ASAP7_75t_L g450 ( 
.A(n_374),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_372),
.B(n_251),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_382),
.B(n_260),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_309),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_364),
.A2(n_323),
.B1(n_312),
.B2(n_310),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_337),
.B(n_237),
.Y(n_458)
);

NOR2x1p5_ASAP7_75t_L g459 ( 
.A(n_395),
.B(n_237),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_405),
.A2(n_379),
.B(n_384),
.C(n_383),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_455),
.A2(n_396),
.B(n_383),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_398),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_419),
.B(n_408),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_403),
.Y(n_464)
);

AO21x1_ASAP7_75t_L g465 ( 
.A1(n_427),
.A2(n_423),
.B(n_406),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_437),
.A2(n_396),
.B(n_391),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_437),
.A2(n_391),
.B(n_397),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_443),
.A2(n_330),
.B(n_333),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_400),
.B(n_357),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_435),
.A2(n_378),
.B1(n_344),
.B2(n_282),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_443),
.A2(n_330),
.B(n_333),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_426),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_401),
.A2(n_344),
.B1(n_282),
.B2(n_310),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

OAI21xp33_ASAP7_75t_L g477 ( 
.A1(n_415),
.A2(n_344),
.B(n_335),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_21),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_441),
.A2(n_340),
.B(n_341),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_435),
.A2(n_323),
.B1(n_310),
.B2(n_312),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_399),
.B(n_22),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_24),
.Y(n_485)
);

AO21x1_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_394),
.B(n_393),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_24),
.Y(n_487)
);

CKINVDCx10_ASAP7_75t_R g488 ( 
.A(n_416),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_418),
.B(n_312),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_430),
.Y(n_490)
);

AO21x1_ASAP7_75t_L g491 ( 
.A1(n_409),
.A2(n_393),
.B(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_25),
.Y(n_493)
);

OR2x6_ASAP7_75t_SL g494 ( 
.A(n_404),
.B(n_26),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_414),
.B(n_320),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_26),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_27),
.Y(n_497)
);

AND2x6_ASAP7_75t_SL g498 ( 
.A(n_413),
.B(n_27),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_452),
.B(n_28),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_29),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_453),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_29),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_457),
.B(n_31),
.Y(n_503)
);

AO22x1_ASAP7_75t_L g504 ( 
.A1(n_447),
.A2(n_324),
.B1(n_34),
.B2(n_35),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_399),
.B(n_360),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_420),
.B(n_32),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_36),
.Y(n_507)
);

AO21x1_ASAP7_75t_L g508 ( 
.A1(n_410),
.A2(n_360),
.B(n_359),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_412),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_447),
.B(n_37),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_431),
.B(n_39),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_153),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_422),
.B(n_47),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_413),
.B(n_140),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g516 ( 
.A(n_459),
.B(n_49),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_50),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_422),
.B(n_53),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_440),
.B(n_57),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_438),
.A2(n_87),
.B(n_91),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_456),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

INVx8_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_492),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_95),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_98),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_473),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_511),
.A2(n_450),
.B(n_102),
.C(n_105),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_480),
.Y(n_530)
);

INVx3_ASAP7_75t_SL g531 ( 
.A(n_488),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_461),
.A2(n_450),
.B(n_113),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_464),
.A2(n_110),
.B1(n_114),
.B2(n_118),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_479),
.A2(n_123),
.B(n_125),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_490),
.B(n_126),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_467),
.A2(n_131),
.B(n_137),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

AO31x2_ASAP7_75t_L g540 ( 
.A1(n_491),
.A2(n_508),
.A3(n_486),
.B(n_466),
.Y(n_540)
);

AO221x1_ASAP7_75t_L g541 ( 
.A1(n_476),
.A2(n_519),
.B1(n_494),
.B2(n_523),
.C(n_520),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_510),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_469),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_469),
.B(n_501),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_515),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

BUFx2_ASAP7_75t_R g548 ( 
.A(n_518),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_505),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_474),
.B(n_487),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_SL g551 ( 
.A(n_481),
.B(n_485),
.C(n_493),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_476),
.B(n_519),
.Y(n_552)
);

AO21x1_ASAP7_75t_L g553 ( 
.A1(n_521),
.A2(n_522),
.B(n_497),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_512),
.B(n_514),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_502),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_499),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_506),
.Y(n_557)
);

AO31x2_ASAP7_75t_L g558 ( 
.A1(n_507),
.A2(n_517),
.A3(n_489),
.B(n_500),
.Y(n_558)
);

AO31x2_ASAP7_75t_L g559 ( 
.A1(n_503),
.A2(n_504),
.A3(n_495),
.B(n_516),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_462),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

OAI21x1_ASAP7_75t_SL g562 ( 
.A1(n_490),
.A2(n_518),
.B(n_513),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_462),
.B(n_402),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_473),
.Y(n_564)
);

AOI221x1_ASAP7_75t_L g565 ( 
.A1(n_467),
.A2(n_466),
.B1(n_437),
.B2(n_477),
.C(n_471),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_462),
.B(n_402),
.Y(n_567)
);

NOR2x1_ASAP7_75t_SL g568 ( 
.A(n_476),
.B(n_399),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_461),
.A2(n_455),
.B(n_352),
.Y(n_569)
);

AO31x2_ASAP7_75t_L g570 ( 
.A1(n_465),
.A2(n_491),
.A3(n_508),
.B(n_467),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_509),
.B(n_462),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_509),
.B(n_462),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_473),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_492),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_509),
.B(n_414),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_509),
.B(n_462),
.Y(n_577)
);

INVx6_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

AO21x1_ASAP7_75t_L g579 ( 
.A1(n_467),
.A2(n_466),
.B(n_468),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_509),
.B(n_414),
.Y(n_580)
);

BUFx4_ASAP7_75t_SL g581 ( 
.A(n_498),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_473),
.B(n_414),
.Y(n_582)
);

NAND3x1_ASAP7_75t_L g583 ( 
.A(n_474),
.B(n_293),
.C(n_429),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_462),
.B(n_402),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_488),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_473),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_509),
.B(n_462),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_473),
.B(n_399),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_460),
.A2(n_509),
.B(n_467),
.C(n_477),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_414),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_492),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_463),
.A2(n_332),
.B(n_347),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_509),
.B(n_414),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_467),
.A2(n_466),
.B(n_427),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_473),
.B(n_414),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_460),
.A2(n_509),
.B(n_467),
.C(n_477),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

AO31x2_ASAP7_75t_L g602 ( 
.A1(n_465),
.A2(n_491),
.A3(n_508),
.B(n_467),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_473),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_470),
.A2(n_401),
.B1(n_404),
.B2(n_426),
.Y(n_604)
);

NOR2x1_ASAP7_75t_SL g605 ( 
.A(n_539),
.B(n_596),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_576),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_533),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_601),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_598),
.A2(n_553),
.B(n_569),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_603),
.Y(n_611)
);

NOR2x1_ASAP7_75t_R g612 ( 
.A(n_584),
.B(n_564),
.Y(n_612)
);

AO21x2_ASAP7_75t_L g613 ( 
.A1(n_591),
.A2(n_562),
.B(n_579),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_601),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

BUFx2_ASAP7_75t_SL g616 ( 
.A(n_542),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_556),
.A2(n_537),
.B(n_534),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_571),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_563),
.B(n_567),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_566),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_594),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_576),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_530),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

AO31x2_ASAP7_75t_L g625 ( 
.A1(n_536),
.A2(n_535),
.A3(n_550),
.B(n_570),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_587),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_580),
.B(n_592),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_527),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

AO31x2_ASAP7_75t_L g630 ( 
.A1(n_570),
.A2(n_602),
.A3(n_540),
.B(n_555),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_577),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_582),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_529),
.A2(n_527),
.B(n_589),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_532),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_583),
.A2(n_557),
.B1(n_546),
.B2(n_547),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_546),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_592),
.B(n_597),
.Y(n_638)
);

OA21x2_ASAP7_75t_L g639 ( 
.A1(n_602),
.A2(n_541),
.B(n_575),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_597),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_599),
.B(n_552),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_593),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_526),
.A2(n_551),
.B(n_543),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_568),
.B(n_530),
.Y(n_644)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_559),
.B(n_544),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_585),
.B(n_590),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_554),
.B(n_545),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

AO21x2_ASAP7_75t_L g649 ( 
.A1(n_558),
.A2(n_559),
.B(n_549),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_558),
.A2(n_524),
.B(n_548),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_578),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_578),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_558),
.A2(n_595),
.B(n_581),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_595),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_531),
.B(n_524),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_576),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_539),
.B(n_596),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_604),
.B(n_462),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_563),
.B(n_402),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_563),
.B(n_402),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_542),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_539),
.A2(n_401),
.B1(n_426),
.B2(n_470),
.Y(n_664)
);

AO31x2_ASAP7_75t_L g665 ( 
.A1(n_565),
.A2(n_579),
.A3(n_600),
.B(n_591),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_539),
.B(n_596),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_541),
.A2(n_470),
.B1(n_523),
.B2(n_477),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_591),
.A2(n_600),
.B(n_467),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_565),
.A2(n_579),
.A3(n_600),
.B(n_591),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_591),
.A2(n_600),
.B(n_467),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_661),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_637),
.B(n_658),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_608),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_615),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_614),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_611),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_657),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_638),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_619),
.B(n_659),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_659),
.B(n_666),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_668),
.A2(n_671),
.B(n_609),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_637),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_638),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_618),
.B(n_631),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_609),
.A2(n_671),
.B(n_668),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_623),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_618),
.B(n_631),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_628),
.B(n_650),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_633),
.A2(n_617),
.B(n_664),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_605),
.B(n_648),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_640),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_630),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_630),
.Y(n_696)
);

AOI221xp5_ASAP7_75t_L g697 ( 
.A1(n_621),
.A2(n_635),
.B1(n_634),
.B2(n_607),
.C(n_669),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_635),
.B(n_640),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_610),
.B(n_620),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_644),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_627),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_667),
.A2(n_621),
.B1(n_628),
.B2(n_647),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_641),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_665),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_665),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_662),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_633),
.A2(n_643),
.B(n_650),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_686),
.B(n_690),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_694),
.B(n_649),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_694),
.B(n_649),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_672),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_684),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_674),
.B(n_639),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_674),
.B(n_613),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_681),
.B(n_629),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_699),
.B(n_636),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_703),
.A2(n_653),
.B1(n_627),
.B2(n_632),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_675),
.B(n_670),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_675),
.B(n_677),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_689),
.B(n_641),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_695),
.Y(n_722)
);

CKINVDCx6p67_ASAP7_75t_R g723 ( 
.A(n_707),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_673),
.B(n_653),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_699),
.B(n_663),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_696),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_696),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_676),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_679),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_691),
.B(n_625),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_698),
.B(n_606),
.Y(n_732)
);

INVx3_ASAP7_75t_SL g733 ( 
.A(n_693),
.Y(n_733)
);

AOI21xp33_ASAP7_75t_L g734 ( 
.A1(n_708),
.A2(n_612),
.B(n_645),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_710),
.B(n_683),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_710),
.B(n_683),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_711),
.B(n_683),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_719),
.B(n_697),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_711),
.B(n_688),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_722),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_719),
.B(n_715),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_715),
.B(n_688),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_733),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_730),
.B(n_704),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_714),
.B(n_688),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_730),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_713),
.Y(n_747)
);

NAND2x1_ASAP7_75t_L g748 ( 
.A(n_730),
.B(n_691),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_720),
.B(n_687),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_724),
.B(n_698),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_713),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_730),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_731),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_739),
.B(n_741),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_751),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_752),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_743),
.B(n_733),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_748),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_739),
.B(n_731),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_743),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_750),
.B(n_724),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_741),
.B(n_731),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_735),
.B(n_731),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_735),
.B(n_705),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_750),
.B(n_726),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_736),
.B(n_727),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_736),
.B(n_705),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_738),
.B(n_728),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_740),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_737),
.B(n_727),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_737),
.B(n_742),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_742),
.B(n_706),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_772),
.B(n_747),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_762),
.B(n_755),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_772),
.B(n_769),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_770),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_766),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_755),
.B(n_745),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_773),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_757),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_766),
.B(n_747),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_762),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_763),
.B(n_752),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_773),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_754),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_767),
.B(n_738),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_783),
.B(n_756),
.Y(n_788)
);

NAND3x2_ASAP7_75t_L g789 ( 
.A(n_775),
.B(n_761),
.C(n_784),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_781),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_787),
.B(n_767),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_779),
.B(n_771),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_778),
.A2(n_764),
.B1(n_760),
.B2(n_763),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_779),
.B(n_771),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_776),
.A2(n_764),
.B1(n_760),
.B2(n_732),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_781),
.B(n_733),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_786),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_774),
.A2(n_732),
.B1(n_765),
.B2(n_768),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_790),
.Y(n_799)
);

AOI322xp5_ASAP7_75t_L g800 ( 
.A1(n_791),
.A2(n_782),
.A3(n_785),
.B1(n_780),
.B2(n_729),
.C1(n_712),
.C2(n_678),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_L g801 ( 
.A1(n_793),
.A2(n_785),
.B(n_780),
.Y(n_801)
);

AOI211x1_ASAP7_75t_SL g802 ( 
.A1(n_788),
.A2(n_734),
.B(n_716),
.C(n_709),
.Y(n_802)
);

OAI322xp33_ASAP7_75t_L g803 ( 
.A1(n_797),
.A2(n_777),
.A3(n_749),
.B1(n_758),
.B2(n_717),
.C1(n_725),
.C2(n_748),
.Y(n_803)
);

NOR4xp25_ASAP7_75t_L g804 ( 
.A(n_799),
.B(n_654),
.C(n_796),
.D(n_721),
.Y(n_804)
);

OAI21xp33_ASAP7_75t_SL g805 ( 
.A1(n_800),
.A2(n_789),
.B(n_794),
.Y(n_805)
);

AOI211xp5_ASAP7_75t_L g806 ( 
.A1(n_803),
.A2(n_654),
.B(n_626),
.C(n_655),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_805),
.B(n_626),
.C(n_652),
.Y(n_807)
);

OAI221xp5_ASAP7_75t_SL g808 ( 
.A1(n_806),
.A2(n_801),
.B1(n_795),
.B2(n_798),
.C(n_691),
.Y(n_808)
);

NAND4xp25_ASAP7_75t_L g809 ( 
.A(n_807),
.B(n_802),
.C(n_718),
.D(n_759),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_808),
.B(n_723),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_810),
.B(n_651),
.C(n_646),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_809),
.B(n_723),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_811),
.B(n_812),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_812),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_814),
.Y(n_815)
);

BUFx8_ASAP7_75t_L g816 ( 
.A(n_813),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_813),
.B(n_662),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_816),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_817),
.A2(n_815),
.B(n_804),
.Y(n_819)
);

XNOR2x1_ASAP7_75t_L g820 ( 
.A(n_815),
.B(n_616),
.Y(n_820)
);

AO21x1_ASAP7_75t_L g821 ( 
.A1(n_817),
.A2(n_792),
.B(n_744),
.Y(n_821)
);

XOR2xp5_ASAP7_75t_L g822 ( 
.A(n_815),
.B(n_701),
.Y(n_822)
);

OAI222xp33_ASAP7_75t_L g823 ( 
.A1(n_818),
.A2(n_691),
.B1(n_759),
.B2(n_704),
.C1(n_744),
.C2(n_685),
.Y(n_823)
);

AOI21xp33_ASAP7_75t_SL g824 ( 
.A1(n_820),
.A2(n_759),
.B(n_685),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_819),
.B(n_777),
.Y(n_825)
);

XNOR2xp5_ASAP7_75t_L g826 ( 
.A(n_822),
.B(n_606),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_821),
.A2(n_622),
.B(n_624),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_818),
.A2(n_704),
.B1(n_744),
.B2(n_746),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_818),
.A2(n_622),
.B(n_624),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_824),
.B(n_704),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_825),
.B(n_753),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_828),
.A2(n_656),
.B1(n_680),
.B2(n_692),
.C(n_682),
.Y(n_832)
);

INVxp33_ASAP7_75t_SL g833 ( 
.A(n_829),
.Y(n_833)
);

AOI221xp5_ASAP7_75t_L g834 ( 
.A1(n_833),
.A2(n_826),
.B1(n_827),
.B2(n_823),
.C(n_656),
.Y(n_834)
);

OA22x2_ASAP7_75t_L g835 ( 
.A1(n_830),
.A2(n_746),
.B1(n_702),
.B2(n_700),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_834),
.B(n_831),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_836),
.A2(n_835),
.B1(n_832),
.B2(n_746),
.Y(n_837)
);


endmodule