module fake_jpeg_27007_n_240 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_28),
.B1(n_23),
.B2(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_14),
.B1(n_23),
.B2(n_15),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_56),
.Y(n_68)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_53),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_52),
.B1(n_27),
.B2(n_29),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_28),
.B1(n_29),
.B2(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_26),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_31),
.B1(n_27),
.B2(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_11),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_17),
.Y(n_69)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_76),
.B1(n_62),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_84),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_27),
.B1(n_44),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_23),
.B1(n_44),
.B2(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_35),
.B1(n_23),
.B2(n_37),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_43),
.Y(n_91)
);

NOR2x1p5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_37),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_24),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_37),
.B1(n_16),
.B2(n_17),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_93),
.B1(n_95),
.B2(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_91),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_103),
.B(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_55),
.B1(n_51),
.B2(n_56),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_52),
.B1(n_62),
.B2(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_12),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_77),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_0),
.C(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_22),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_22),
.A3(n_20),
.B1(n_63),
.B2(n_21),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_16),
.B1(n_19),
.B2(n_17),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_66),
.B1(n_64),
.B2(n_17),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_72),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_20),
.B(n_22),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_81),
.B(n_70),
.C(n_66),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_118),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_115),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_66),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_125),
.B1(n_118),
.B2(n_126),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_133),
.B1(n_86),
.B2(n_107),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_123),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_49),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_134),
.C(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_21),
.B(n_19),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_65),
.B(n_1),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_20),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_64),
.B1(n_16),
.B2(n_67),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_49),
.C(n_24),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_18),
.B(n_11),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_49),
.C(n_65),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_148),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_95),
.C(n_86),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_112),
.C(n_132),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_160),
.B1(n_137),
.B2(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_119),
.B1(n_85),
.B2(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_112),
.B1(n_117),
.B2(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_97),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_106),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_88),
.B(n_135),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_173),
.B1(n_171),
.B2(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_154),
.B1(n_151),
.B2(n_152),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_117),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_179),
.B(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_65),
.B1(n_16),
.B2(n_67),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_177),
.B1(n_181),
.B2(n_158),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_157),
.B1(n_148),
.B2(n_149),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_49),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_138),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_0),
.B(n_2),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_19),
.B1(n_18),
.B2(n_11),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_142),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_141),
.A3(n_146),
.B1(n_145),
.B2(n_143),
.C1(n_138),
.C2(n_144),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_188),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_192),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_144),
.B(n_163),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_176),
.B1(n_175),
.B2(n_165),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_193),
.B1(n_183),
.B2(n_194),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_196),
.B1(n_181),
.B2(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_12),
.C(n_19),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_168),
.C(n_167),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_18),
.B1(n_12),
.B2(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_182),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_187),
.C(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_179),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_191),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_2),
.C(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_191),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_4),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_214),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_187),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_5),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_197),
.B1(n_199),
.B2(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_5),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_202),
.B(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_198),
.B(n_6),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_5),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_215),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_231),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_210),
.B(n_6),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_222),
.B(n_6),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_234),
.B1(n_227),
.B2(n_228),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_225),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_5),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_7),
.B(n_8),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_237),
.B(n_232),
.Y(n_238)
);

NOR4xp25_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_8),
.C(n_9),
.D(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_8),
.Y(n_240)
);


endmodule