module real_jpeg_26830_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_38;
wire n_35;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_76;
wire n_58;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_75;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_71;
wire n_47;
wire n_45;
wire n_25;
wire n_51;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_70;
wire n_74;
wire n_26;
wire n_32;
wire n_56;
wire n_48;
wire n_19;
wire n_20;
wire n_27;
wire n_41;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_5),
.B(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_1),
.A2(n_15),
.B1(n_18),
.B2(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_16),
.B1(n_17),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_4),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_71)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_16),
.B1(n_17),
.B2(n_40),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_7),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_56),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_44),
.B(n_55),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_26),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_13),
.B(n_26),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_20),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_15),
.A2(n_24),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_18),
.Y(n_15)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_16),
.A2(n_17),
.B1(n_34),
.B2(n_35),
.Y(n_36)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_38),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_42),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_29),
.A2(n_36),
.B1(n_39),
.B2(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_35),
.B(n_38),
.C(n_43),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_54),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_76),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);


endmodule