module fake_jpeg_12359_n_24 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

INVx1_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_11),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_16),
.B(n_10),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_13),
.B1(n_5),
.B2(n_9),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_18),
.A2(n_19),
.B1(n_13),
.B2(n_6),
.Y(n_20)
);

OAI211xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.C(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_20),
.C(n_7),
.Y(n_24)
);


endmodule