module fake_jpeg_19148_n_258 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_47),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_20),
.A3(n_18),
.B1(n_22),
.B2(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_31),
.B1(n_34),
.B2(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_57),
.B1(n_44),
.B2(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_35),
.B1(n_44),
.B2(n_39),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_33),
.B2(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_65),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_41),
.B1(n_26),
.B2(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_20),
.B(n_18),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_18),
.B(n_12),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_90),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_53),
.B1(n_52),
.B2(n_54),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_59),
.C(n_48),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_14),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_60),
.B1(n_43),
.B2(n_54),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_97),
.B1(n_65),
.B2(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_71),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_62),
.B(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_43),
.B1(n_26),
.B2(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_100),
.B(n_103),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_97),
.B1(n_87),
.B2(n_91),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_70),
.B(n_79),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_77),
.B(n_80),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_63),
.B1(n_74),
.B2(n_73),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_109),
.B1(n_87),
.B2(n_67),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_68),
.B1(n_67),
.B2(n_78),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_68),
.B(n_71),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_29),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_114),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_71),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_110),
.Y(n_125)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_126),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_127),
.B1(n_104),
.B2(n_135),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_103),
.B(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_95),
.B1(n_61),
.B2(n_37),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_109),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_20),
.C(n_7),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_37),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_139),
.B(n_132),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_102),
.B1(n_104),
.B2(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_158),
.B1(n_139),
.B2(n_66),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_107),
.C(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_153),
.C(n_157),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_105),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_22),
.B(n_29),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_138),
.B1(n_137),
.B2(n_126),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_71),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_156),
.B1(n_162),
.B2(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_58),
.C(n_24),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_58),
.B1(n_66),
.B2(n_21),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_24),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_161),
.C(n_129),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_19),
.C(n_13),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_176),
.B1(n_178),
.B2(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_172),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_182),
.B(n_12),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_181),
.B1(n_0),
.B2(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_159),
.B1(n_143),
.B2(n_153),
.Y(n_176)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_9),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_161),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_150),
.C(n_25),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.C(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_25),
.C(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_22),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_25),
.C(n_19),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_25),
.C(n_19),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_19),
.C(n_13),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_168),
.B1(n_173),
.B2(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_1),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_10),
.B(n_11),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_6),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_165),
.B1(n_167),
.B2(n_176),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_185),
.B1(n_189),
.B2(n_204),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_190),
.B1(n_188),
.B2(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_177),
.C(n_19),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_6),
.B1(n_7),
.B2(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_194),
.B(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_199),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_206),
.B(n_208),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_195),
.B1(n_192),
.B2(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_17),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_211),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_13),
.C(n_19),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_17),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_13),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_232),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_17),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_239),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_222),
.A3(n_231),
.B1(n_234),
.B2(n_226),
.C(n_22),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_241),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_222),
.C(n_13),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_13),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_242),
.B(n_13),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_247),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_22),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_236),
.C(n_23),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_12),
.Y(n_247)
);

AOI21x1_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_244),
.B(n_3),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_236),
.B(n_3),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_246),
.B(n_23),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_252),
.B(n_250),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_2),
.B(n_3),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_2),
.B1(n_5),
.B2(n_207),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_2),
.Y(n_258)
);


endmodule