module fake_jpeg_14290_n_611 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g192 ( 
.A(n_72),
.Y(n_192)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_75),
.B(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_80),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_84),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_88),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_100),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g180 ( 
.A(n_97),
.B(n_47),
.Y(n_180)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_11),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_29),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_120),
.Y(n_133)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_26),
.Y(n_166)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_9),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_75),
.Y(n_140)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_127),
.Y(n_205)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_57),
.B1(n_38),
.B2(n_36),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_130),
.A2(n_149),
.B(n_47),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_29),
.Y(n_139)
);

NAND2x1_ASAP7_75t_SL g263 ( 
.A(n_139),
.B(n_0),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_34),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_60),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_144),
.B(n_145),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_60),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_86),
.A2(n_57),
.B1(n_36),
.B2(n_28),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_39),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_150),
.B(n_166),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_SL g153 ( 
.A(n_64),
.Y(n_153)
);

INVx11_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_47),
.B1(n_57),
.B2(n_59),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_154),
.A2(n_47),
.B1(n_46),
.B2(n_41),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_66),
.B(n_26),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_171),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_68),
.B(n_56),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_70),
.B(n_24),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_172),
.B(n_176),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_43),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_43),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_177),
.A2(n_194),
.B(n_14),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_180),
.Y(n_225)
);

INVx6_ASAP7_75t_SL g187 ( 
.A(n_72),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g273 ( 
.A(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_91),
.B(n_56),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_40),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_198),
.B(n_208),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_93),
.B(n_55),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_223),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_141),
.A2(n_58),
.B1(n_44),
.B2(n_55),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_213),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_214),
.B(n_237),
.Y(n_327)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_215),
.Y(n_312)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_81),
.B1(n_80),
.B2(n_84),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_217),
.A2(n_231),
.B1(n_195),
.B2(n_189),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_52),
.B1(n_41),
.B2(n_28),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_218),
.A2(n_269),
.B1(n_272),
.B2(n_178),
.Y(n_323)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_219),
.Y(n_342)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_222),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_224),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_129),
.B(n_59),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_260),
.Y(n_288)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_228),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_112),
.B1(n_111),
.B2(n_89),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_229),
.A2(n_253),
.B1(n_203),
.B2(n_189),
.Y(n_287)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_230),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_154),
.A2(n_115),
.B1(n_88),
.B2(n_85),
.Y(n_231)
);

AO21x1_ASAP7_75t_SL g294 ( 
.A1(n_232),
.A2(n_178),
.B(n_192),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_233),
.Y(n_331)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_234),
.Y(n_334)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_47),
.B(n_40),
.C(n_33),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_238),
.Y(n_341)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_175),
.A2(n_46),
.B1(n_41),
.B2(n_36),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_242),
.A2(n_254),
.B(n_278),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_261),
.B1(n_280),
.B2(n_199),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

BUFx24_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_197),
.A2(n_46),
.B1(n_33),
.B2(n_23),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_149),
.A2(n_205),
.B(n_199),
.Y(n_254)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_255),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_135),
.B(n_23),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_259),
.C(n_16),
.Y(n_336)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_267),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_185),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_262),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_142),
.B(n_23),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_0),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_202),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_170),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_263),
.B(n_152),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_266),
.B(n_178),
.C(n_201),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.C(n_5),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_275),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_175),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_190),
.B(n_1),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_221),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_162),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_274),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_131),
.A2(n_15),
.B1(n_6),
.B2(n_12),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_200),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_277),
.B(n_284),
.Y(n_315)
);

NAND2x1p5_ASAP7_75t_L g278 ( 
.A(n_158),
.B(n_1),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_167),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_146),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_282),
.Y(n_321)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_165),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_283),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_297),
.B1(n_302),
.B2(n_316),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_291),
.B(n_273),
.Y(n_378)
);

OR2x2_ASAP7_75t_SL g292 ( 
.A(n_263),
.B(n_147),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_319),
.C(n_293),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_278),
.B(n_237),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_238),
.A2(n_174),
.B1(n_169),
.B2(n_148),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_336),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_248),
.A2(n_173),
.B1(n_191),
.B2(n_207),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_307),
.A2(n_310),
.B1(n_314),
.B2(n_338),
.Y(n_381)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_173),
.B(n_203),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_225),
.A2(n_260),
.B1(n_270),
.B2(n_261),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_232),
.A2(n_207),
.B1(n_191),
.B2(n_206),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_162),
.B1(n_211),
.B2(n_163),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_322),
.B1(n_325),
.B2(n_329),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_225),
.A2(n_158),
.B1(n_165),
.B2(n_152),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_151),
.B1(n_16),
.B2(n_17),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_226),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_264),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_284),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_256),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_229),
.A2(n_18),
.B1(n_242),
.B2(n_253),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_266),
.B(n_265),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_256),
.A2(n_18),
.B1(n_259),
.B2(n_214),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_224),
.B(n_246),
.C(n_236),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_240),
.C(n_259),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_214),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_345),
.C(n_356),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_303),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_243),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_289),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_348),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_285),
.B(n_227),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_250),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_314),
.A2(n_304),
.B1(n_310),
.B2(n_306),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_352),
.A2(n_355),
.B1(n_359),
.B2(n_366),
.Y(n_421)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_353),
.A2(n_286),
.B(n_330),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_362),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_304),
.A2(n_252),
.B1(n_257),
.B2(n_219),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_340),
.B(n_251),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_296),
.C(n_293),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_358),
.B(n_361),
.C(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_216),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_220),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_367),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_327),
.B(n_275),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_310),
.A2(n_234),
.B1(n_228),
.B2(n_239),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_277),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_295),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_368),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_222),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_374),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_294),
.A2(n_222),
.B(n_215),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_378),
.B(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_271),
.B(n_273),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_373),
.A2(n_322),
.B(n_286),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_281),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_301),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_376),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_336),
.C(n_342),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_244),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_379),
.Y(n_407)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_295),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_307),
.A2(n_230),
.B1(n_282),
.B2(n_267),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_385),
.A2(n_311),
.B1(n_321),
.B2(n_324),
.Y(n_424)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_299),
.Y(n_387)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

A2O1A1Ixp33_ASAP7_75t_SL g441 ( 
.A1(n_390),
.A2(n_396),
.B(n_400),
.C(n_385),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_376),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_338),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_410),
.C(n_416),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g396 ( 
.A1(n_362),
.A2(n_291),
.B1(n_316),
.B2(n_337),
.Y(n_396)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_292),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_382),
.A2(n_298),
.B1(n_321),
.B2(n_311),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_342),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_352),
.A2(n_298),
.B1(n_291),
.B2(n_287),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_412),
.A2(n_351),
.B1(n_375),
.B2(n_382),
.Y(n_435)
);

BUFx8_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_413),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_419),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_303),
.C(n_300),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_417),
.A2(n_305),
.B(n_335),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_343),
.B(n_300),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_295),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_375),
.C(n_344),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_424),
.A2(n_366),
.B1(n_381),
.B2(n_367),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_399),
.B(n_363),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g486 ( 
.A(n_427),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_428),
.A2(n_443),
.B1(n_396),
.B2(n_398),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_431),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_378),
.B(n_370),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_432),
.A2(n_441),
.B(n_445),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_354),
.A3(n_355),
.B1(n_353),
.B2(n_381),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_437),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_440),
.B1(n_444),
.B2(n_446),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_415),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_442),
.C(n_458),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_399),
.B(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_421),
.A2(n_351),
.B1(n_384),
.B2(n_368),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_389),
.C(n_420),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_395),
.A2(n_365),
.B1(n_359),
.B2(n_350),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_421),
.A2(n_384),
.B1(n_365),
.B2(n_359),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_407),
.A2(n_365),
.B1(n_369),
.B2(n_346),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_390),
.A2(n_372),
.B1(n_371),
.B2(n_387),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_380),
.Y(n_447)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_449),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_397),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_459),
.C(n_439),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_400),
.A2(n_374),
.B1(n_324),
.B2(n_331),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_451),
.A2(n_456),
.B1(n_424),
.B2(n_388),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_400),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_406),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_453),
.B(n_413),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_305),
.Y(n_454)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_454),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_400),
.A2(n_331),
.B1(n_233),
.B2(n_249),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_320),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_334),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_430),
.B(n_411),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_469),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_447),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_463),
.B(n_459),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_465),
.A2(n_476),
.B(n_489),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_468),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_428),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_429),
.B(n_394),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_482),
.Y(n_496)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_416),
.C(n_401),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_431),
.Y(n_505)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_396),
.B1(n_413),
.B2(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_403),
.Y(n_477)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_477),
.Y(n_511)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_419),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_440),
.B1(n_444),
.B2(n_451),
.Y(n_493)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_410),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_445),
.C(n_458),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_455),
.B(n_404),
.Y(n_487)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_435),
.A2(n_396),
.B1(n_422),
.B2(n_405),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_454),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_446),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_491),
.B(n_505),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_493),
.A2(n_513),
.B1(n_514),
.B2(n_475),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_427),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_497),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_448),
.C(n_433),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_515),
.C(n_517),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_499),
.Y(n_529)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_477),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_504),
.B(n_510),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_489),
.A2(n_443),
.B1(n_432),
.B2(n_434),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_426),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_516),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_486),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_460),
.A2(n_456),
.B1(n_441),
.B2(n_448),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_460),
.A2(n_441),
.B1(n_453),
.B2(n_436),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_473),
.B(n_441),
.C(n_436),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_441),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_405),
.C(n_392),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_423),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_334),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_492),
.A2(n_467),
.B(n_476),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_521),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_492),
.A2(n_467),
.B(n_502),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_503),
.A2(n_461),
.B1(n_478),
.B2(n_490),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_466),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_528),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_496),
.B(n_485),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_531),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_482),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_481),
.C(n_462),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_536),
.C(n_491),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_512),
.B(n_466),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_534),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_498),
.B(n_461),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_471),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_535),
.B(n_540),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_471),
.C(n_488),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_493),
.A2(n_472),
.B1(n_488),
.B2(n_479),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_501),
.C(n_513),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_518),
.Y(n_542)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_542),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_505),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_543),
.B(n_546),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_531),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_536),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_516),
.C(n_501),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_548),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_520),
.C(n_526),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_550),
.B(n_556),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_514),
.C(n_500),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_553),
.C(n_557),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_506),
.C(n_511),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_526),
.B(n_495),
.C(n_509),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_495),
.C(n_508),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_525),
.B(n_508),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_555),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_562),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_554),
.A2(n_519),
.B(n_524),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_564),
.B(n_573),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_537),
.C(n_539),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_568),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_544),
.A2(n_521),
.B(n_522),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_566),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_539),
.C(n_540),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_551),
.A2(n_524),
.B1(n_522),
.B2(n_507),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_571),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_541),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_507),
.B1(n_423),
.B2(n_331),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_559),
.B(n_328),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_574),
.B(n_549),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_557),
.A2(n_328),
.B1(n_247),
.B2(n_241),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_575),
.B(n_332),
.Y(n_578)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_577),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_579),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_545),
.C(n_328),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_572),
.B(n_317),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_583),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_317),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_563),
.A2(n_328),
.B(n_255),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_584),
.B(n_587),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_313),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_564),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_588),
.B(n_589),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_585),
.B(n_560),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_580),
.B(n_571),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_591),
.B(n_592),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_586),
.B(n_565),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_SL g595 ( 
.A1(n_581),
.A2(n_562),
.B(n_566),
.C(n_567),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_595),
.A2(n_593),
.B(n_596),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_594),
.A2(n_581),
.B(n_576),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_598),
.B(n_599),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_590),
.A2(n_568),
.B(n_574),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_602),
.C(n_326),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_595),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_235),
.C(n_312),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_603),
.Y(n_606)
);

NAND4xp25_ASAP7_75t_SL g607 ( 
.A(n_604),
.B(n_597),
.C(n_332),
.D(n_312),
.Y(n_607)
);

AO21x2_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_605),
.B(n_235),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_606),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_313),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_610),
.B(n_283),
.Y(n_611)
);


endmodule