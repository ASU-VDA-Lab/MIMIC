module fake_jpeg_21918_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_13),
.B1(n_29),
.B2(n_31),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_26),
.B(n_13),
.C(n_29),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_14),
.B1(n_22),
.B2(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_70),
.Y(n_79)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_78),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_76),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_54),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_26),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_54),
.C(n_42),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_47),
.B(n_50),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_43),
.B1(n_48),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_61),
.B1(n_70),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_94),
.B1(n_95),
.B2(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_42),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_24),
.B1(n_16),
.B2(n_48),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_46),
.Y(n_114)
);

NOR2x1_ASAP7_75t_R g94 ( 
.A(n_77),
.B(n_43),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_48),
.B1(n_29),
.B2(n_13),
.Y(n_95)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_60),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_72),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_100),
.B(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_121),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_113),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_119),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_52),
.B1(n_51),
.B2(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_64),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_52),
.B1(n_51),
.B2(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_46),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_33),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_33),
.Y(n_137)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_64),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_91),
.B1(n_97),
.B2(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_97),
.B1(n_91),
.B2(n_84),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_80),
.B(n_94),
.C(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_101),
.B(n_86),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_145),
.B(n_150),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_85),
.C(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_85),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_97),
.B1(n_85),
.B2(n_88),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_144),
.B1(n_60),
.B2(n_65),
.Y(n_165)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_85),
.B1(n_62),
.B2(n_69),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_13),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_69),
.B1(n_60),
.B2(n_65),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_52),
.B1(n_67),
.B2(n_58),
.Y(n_148)
);

XOR2x2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_62),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_153),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_102),
.B1(n_124),
.B2(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_133),
.B1(n_130),
.B2(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_170),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_105),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_131),
.B(n_125),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_117),
.B1(n_111),
.B2(n_112),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_167),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_62),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_116),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_116),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_32),
.C(n_36),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_174),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_121),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_136),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_176),
.B1(n_150),
.B2(n_131),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_183),
.B1(n_187),
.B2(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_195),
.B(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_185),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_190),
.B1(n_192),
.B2(n_173),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_133),
.B1(n_144),
.B2(n_132),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_165),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_137),
.B1(n_145),
.B2(n_67),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_58),
.B1(n_78),
.B2(n_51),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_49),
.C(n_34),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_197),
.C(n_155),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_0),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_49),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_66),
.B1(n_55),
.B2(n_14),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_24),
.B1(n_14),
.B2(n_66),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_215),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_208),
.B(n_226),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_152),
.B(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_153),
.B(n_167),
.C(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_220),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_218),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_159),
.C(n_167),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_208),
.C(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_179),
.B1(n_199),
.B2(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_188),
.B1(n_186),
.B2(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_233),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_182),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_205),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_184),
.B(n_181),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_209),
.B(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_213),
.B1(n_23),
.B2(n_20),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_246),
.C(n_213),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_225),
.B1(n_212),
.B2(n_220),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_242),
.B1(n_244),
.B2(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_199),
.B1(n_189),
.B2(n_201),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_159),
.B1(n_195),
.B2(n_66),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_17),
.B1(n_26),
.B2(n_20),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_195),
.B1(n_55),
.B2(n_23),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_21),
.C(n_26),
.Y(n_246)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_205),
.B1(n_219),
.B2(n_215),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_261),
.B1(n_264),
.B2(n_0),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_237),
.B(n_211),
.CI(n_222),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_265),
.C(n_229),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_12),
.B(n_1),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_37),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_37),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_27),
.B1(n_20),
.B2(n_19),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_36),
.B1(n_32),
.B2(n_27),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_235),
.B1(n_246),
.B2(n_236),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_19),
.B(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_4),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_279),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_3),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_0),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_253),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_285),
.B(n_293),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_250),
.B1(n_254),
.B2(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_263),
.C(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_271),
.C(n_269),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_257),
.B1(n_261),
.B2(n_3),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_6),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_4),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_304),
.C(n_6),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_273),
.B(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_281),
.B(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_281),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_287),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_26),
.B(n_7),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_6),
.B(n_8),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_312),
.C(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_303),
.B(n_300),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_307),
.B(n_10),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.C(n_9),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_305),
.B(n_26),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.C(n_10),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_11),
.C(n_9),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_11),
.B(n_9),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_11),
.B(n_9),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_10),
.C(n_321),
.Y(n_325)
);


endmodule