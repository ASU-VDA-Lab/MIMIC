module fake_jpeg_15341_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_25),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_54),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_31),
.Y(n_104)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_43),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_25),
.A3(n_33),
.B1(n_29),
.B2(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_20),
.B1(n_33),
.B2(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_45),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_36),
.B1(n_39),
.B2(n_45),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_93),
.B1(n_56),
.B2(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_92),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_36),
.B1(n_69),
.B2(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_2),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_2),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_4),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_53),
.A2(n_31),
.A3(n_18),
.B1(n_16),
.B2(n_7),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_99),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_115),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_57),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_127),
.B(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_4),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_129),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_5),
.B(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_76),
.A2(n_92),
.B1(n_102),
.B2(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_75),
.B1(n_49),
.B2(n_62),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_97),
.C(n_95),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_105),
.C(n_81),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_149),
.B(n_125),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.C(n_144),
.Y(n_167)
);

NOR2x1_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_85),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_112),
.B(n_111),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_7),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_84),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_155),
.B1(n_132),
.B2(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_87),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_91),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_107),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_75),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_114),
.B1(n_121),
.B2(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_8),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_8),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_15),
.C(n_12),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_118),
.C(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_9),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_9),
.Y(n_170)
);

XNOR2x2_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_127),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_14),
.B(n_15),
.C(n_168),
.D(n_181),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_112),
.B(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_182),
.B1(n_9),
.B2(n_13),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_155),
.B1(n_153),
.B2(n_152),
.C(n_136),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_135),
.B(n_156),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_170),
.B(n_161),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_183),
.B1(n_137),
.B2(n_158),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_14),
.B1(n_164),
.B2(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_109),
.B1(n_124),
.B2(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_131),
.B(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_131),
.C(n_13),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_140),
.C(n_159),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_199),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_205),
.B(n_206),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_142),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_138),
.C(n_148),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_162),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_137),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_136),
.C(n_141),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_183),
.B1(n_177),
.B2(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_171),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_178),
.B(n_174),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_185),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_198),
.B1(n_175),
.B2(n_204),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_200),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_205),
.C(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_191),
.B1(n_200),
.B2(n_203),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_218),
.B1(n_214),
.B2(n_207),
.Y(n_240)
);

OAI31xp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_220),
.A3(n_217),
.B(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_192),
.C(n_186),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_176),
.C(n_180),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_209),
.C(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_238),
.C(n_243),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_225),
.B(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_212),
.C(n_208),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_208),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_232),
.C(n_226),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_235),
.C(n_242),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_251),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_247),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_201),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_227),
.B1(n_162),
.B2(n_182),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_245),
.B1(n_251),
.B2(n_163),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_260),
.B(n_163),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_259),
.C(n_256),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.C(n_170),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_253),
.Y(n_264)
);


endmodule