module fake_netlist_6_398_n_4819 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_1061, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_1072, n_677, n_969, n_988, n_805, n_396, n_495, n_1065, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_1071, n_628, n_1067, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1074, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_1057, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_1058, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_1070, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1073, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_1062, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_1048, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_1068, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_1075, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_1064, n_403, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_1066, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_1060, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_1055, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_1069, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_1052, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_1063, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_1059, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_4819);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_1061;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1072;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_1065;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_1071;
input n_628;
input n_1067;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1074;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_1057;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_1058;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_1070;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1073;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_1062;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_1068;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_1075;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_1064;
input n_403;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_1066;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_1060;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_1069;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_1052;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_1063;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_1059;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_4819;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_4730;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_4598;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4649;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_4670;
wire n_3266;
wire n_1351;
wire n_3574;
wire n_4620;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_4738;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_3178;
wire n_1307;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1581;
wire n_4504;
wire n_3844;
wire n_4395;
wire n_1237;
wire n_2534;
wire n_2353;
wire n_3301;
wire n_3089;
wire n_4388;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_2324;
wire n_1575;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_4815;
wire n_3257;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_2260;
wire n_1387;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_4699;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_4686;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_4645;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_4755;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_4777;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4591;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_4702;
wire n_2291;
wire n_4754;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1371;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_3626;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3757;
wire n_3904;
wire n_1590;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_2247;
wire n_3106;
wire n_1711;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_4666;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_4617;
wire n_4733;
wire n_2129;
wire n_2340;
wire n_4764;
wire n_1261;
wire n_4724;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_4743;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_4696;
wire n_4692;
wire n_1572;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_4814;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_2510;
wire n_2739;
wire n_3890;
wire n_2480;
wire n_1300;
wire n_3023;
wire n_1541;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3750;
wire n_3607;
wire n_4325;
wire n_3251;
wire n_3877;
wire n_3316;
wire n_4602;
wire n_2212;
wire n_3929;
wire n_3048;
wire n_3063;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1455;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_4767;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_4722;
wire n_4606;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1971;
wire n_1781;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_2873;
wire n_1345;
wire n_3452;
wire n_3655;
wire n_1820;
wire n_4563;
wire n_3107;
wire n_4556;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_4687;
wire n_3948;
wire n_2836;
wire n_3664;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_4619;
wire n_2378;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_4600;
wire n_4125;
wire n_2625;
wire n_3296;
wire n_1400;
wire n_4646;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_4262;
wire n_1088;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_4729;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_3999;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_4751;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_4605;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_4691;
wire n_1558;
wire n_3943;
wire n_2300;
wire n_1986;
wire n_1732;
wire n_4320;
wire n_4305;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_3871;
wire n_2190;
wire n_1918;
wire n_3603;
wire n_1641;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_4662;
wire n_1843;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_4314;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_3728;
wire n_2669;
wire n_2925;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_4677;
wire n_3272;
wire n_4765;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_1302;
wire n_1599;
wire n_1543;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_1762;
wire n_4641;
wire n_1910;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_4795;
wire n_3630;
wire n_4698;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_4792;
wire n_4810;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_3914;
wire n_3514;
wire n_2228;
wire n_1605;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_2714;
wire n_1289;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_4742;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1865;
wire n_1111;
wire n_2971;
wire n_1713;
wire n_4375;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_4613;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_2818;
wire n_1359;
wire n_2428;
wire n_3581;
wire n_4717;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_4585;
wire n_4731;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_4773;
wire n_3933;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3346;
wire n_2254;
wire n_2345;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_1747;
wire n_3691;
wire n_4427;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_4681;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_4072;
wire n_3940;
wire n_1655;
wire n_4220;
wire n_4523;
wire n_4752;
wire n_2347;
wire n_1214;
wire n_3917;
wire n_2092;
wire n_1886;
wire n_1654;
wire n_4371;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_2994;
wire n_1750;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4673;
wire n_4313;
wire n_2916;
wire n_3415;
wire n_4292;
wire n_4607;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_3873;
wire n_1624;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_4510;
wire n_1515;
wire n_4473;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_3009;
wire n_1709;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_3578;
wire n_1369;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_4737;
wire n_4685;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_4675;
wire n_2794;
wire n_3352;
wire n_2663;
wire n_1990;
wire n_1296;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_3696;
wire n_3780;
wire n_1420;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_3337;
wire n_3253;
wire n_1767;
wire n_1779;
wire n_3431;
wire n_1465;
wire n_3450;
wire n_4002;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_3021;
wire n_1712;
wire n_4603;
wire n_1391;
wire n_4663;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_1523;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_4697;
wire n_1735;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2712;
wire n_2684;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1100;
wire n_4588;
wire n_4653;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_2230;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_2535;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_4636;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_2693;
wire n_1293;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_4701;
wire n_4651;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_4576;
wire n_3727;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_4615;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_3293;
wire n_1646;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_4661;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4621;
wire n_4216;
wire n_3608;
wire n_4540;
wire n_4664;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_4284;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3353;
wire n_3150;
wire n_3018;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_4785;
wire n_3470;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4713;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_4688;
wire n_3166;
wire n_4753;
wire n_2316;
wire n_1771;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1707;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_4775;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_4674;
wire n_2191;
wire n_2717;
wire n_1723;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_3580;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3775;
wire n_3537;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_4634;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2667;
wire n_2698;
wire n_2539;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_3119;
wire n_1809;
wire n_4280;
wire n_2958;
wire n_2948;
wire n_1577;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_4718;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4627;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_2403;
wire n_3342;
wire n_4624;
wire n_2837;
wire n_4175;
wire n_4700;
wire n_4818;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_4659;
wire n_4771;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_2127;
wire n_2338;
wire n_1178;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3867;
wire n_3341;
wire n_4455;
wire n_4453;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_3191;
wire n_1626;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_4798;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_3987;
wire n_1857;
wire n_4806;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_2296;
wire n_1284;
wire n_3201;
wire n_3633;
wire n_1604;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_1201;
wire n_3103;
wire n_3638;
wire n_1398;
wire n_4573;
wire n_4592;
wire n_4816;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_3480;
wire n_3451;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_4695;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_4796;
wire n_3606;
wire n_3142;
wire n_1310;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3641;
wire n_3591;
wire n_3777;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_1314;
wire n_4533;
wire n_4756;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_1410;
wire n_4746;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_4658;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3944;
wire n_3909;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1785;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_4665;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_4654;
wire n_4633;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_4362;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_1773;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_4597;
wire n_1783;
wire n_1533;
wire n_2929;
wire n_3226;
wire n_2780;
wire n_3364;
wire n_3323;
wire n_1597;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_4404;
wire n_1153;
wire n_3407;
wire n_1618;
wire n_1531;
wire n_4618;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_4679;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_4805;
wire n_4063;
wire n_1679;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_1374;
wire n_2556;
wire n_4706;
wire n_2648;
wire n_4747;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_3188;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_1459;
wire n_4410;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1933;
wire n_3683;
wire n_4034;
wire n_4056;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_4622;
wire n_4721;
wire n_4807;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_4693;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_3284;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_1881;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_2720;
wire n_1520;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1733;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_3051;
wire n_1636;
wire n_1437;
wire n_4614;
wire n_4609;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_4707;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_2627;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_2777;
wire n_1134;
wire n_1668;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_4647;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_4126;
wire n_1129;
wire n_3870;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_4655;
wire n_1429;
wire n_4632;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_4470;
wire n_3466;
wire n_4801;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_4813;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_2942;
wire n_1635;
wire n_4014;
wire n_1079;
wire n_4714;
wire n_4704;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_4374;
wire n_2201;
wire n_3919;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_4668;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4635;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_3886;
wire n_2924;
wire n_4761;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_4710;
wire n_1510;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_1270;
wire n_2549;
wire n_4690;
wire n_1187;
wire n_4405;
wire n_4304;
wire n_4234;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_4759;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4667;
wire n_4182;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_3592;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_4656;
wire n_1841;
wire n_4660;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4637;
wire n_4274;
wire n_2423;
wire n_3277;
wire n_4797;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4270;
wire n_4189;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_3730;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_3011;
wire n_1601;
wire n_1960;
wire n_4808;
wire n_2694;
wire n_2061;
wire n_4611;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_4610;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_2716;
wire n_3249;
wire n_1320;
wire n_3657;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_3672;
wire n_2854;
wire n_1452;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4725;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_3137;
wire n_3382;
wire n_1535;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_3177;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_2472;
wire n_1262;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_1891;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_3424;
wire n_2894;
wire n_1272;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_4554;
wire n_3594;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_4778;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_2373;
wire n_1472;
wire n_4626;
wire n_4595;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_2964;
wire n_1870;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_4734;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_4680;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_4689;
wire n_4616;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_2699;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1828;
wire n_4258;
wire n_4547;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_4643;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_4601;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_3681;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_4623;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3988;
wire n_1974;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_3307;
wire n_1637;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_4135;
wire n_2768;
wire n_1795;
wire n_4279;
wire n_2871;
wire n_4209;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_3858;
wire n_1845;
wire n_4183;
wire n_4321;
wire n_1489;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_4644;
wire n_4790;
wire n_2258;
wire n_1485;
wire n_1544;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_2310;
wire n_4608;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_4716;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_4757;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_2195;
wire n_3208;
wire n_1633;
wire n_2809;
wire n_3007;
wire n_3528;
wire n_2172;
wire n_4682;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4715;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_3102;
wire n_1948;
wire n_4694;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_4672;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_4604;
wire n_2939;
wire n_4782;
wire n_3305;
wire n_1484;
wire n_2992;
wire n_1906;
wire n_1321;
wire n_1241;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1672;
wire n_4185;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4407;
wire n_4378;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_4774;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_2668;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_4776;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_4726;
wire n_1794;
wire n_1650;
wire n_1962;
wire n_1236;
wire n_3506;
wire n_2398;
wire n_3855;
wire n_1928;
wire n_1559;
wire n_3743;
wire n_1725;
wire n_1872;
wire n_3091;
wire n_4736;
wire n_4317;
wire n_4493;
wire n_4723;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_4315;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2923;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_1804;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_4650;
wire n_4788;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_4421;
wire n_1477;
wire n_4719;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_4793;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_4799;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_4789;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_3621;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_4505;
wire n_4657;
wire n_4708;
wire n_1562;
wire n_1690;
wire n_4365;
wire n_1191;
wire n_1826;
wire n_2951;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1929;
wire n_1807;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4741;
wire n_4543;
wire n_3343;
wire n_3303;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4630;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_4652;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_2358;
wire n_1401;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_4748;
wire n_4439;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_4783;
wire n_3874;
wire n_2814;
wire n_2528;
wire n_1379;
wire n_4639;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_3027;
wire n_3231;
wire n_1554;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4786;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_4579;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4811;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_4112;
wire n_4009;
wire n_1114;
wire n_3268;
wire n_1147;
wire n_1848;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_1754;
wire n_2584;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_4557;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_4593;
wire n_2906;
wire n_2769;
wire n_1303;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1721;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_2180;
wire n_1689;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_3604;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_4711;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_4740;
wire n_2117;
wire n_2234;
wire n_4631;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_4720;
wire n_1656;
wire n_3494;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_2430;
wire n_3584;
wire n_1464;
wire n_3486;
wire n_1414;
wire n_4678;
wire n_4086;
wire n_2649;
wire n_2721;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_4625;
wire n_4812;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_4766;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_3362;
wire n_2242;
wire n_1253;
wire n_1266;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4744;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_4817;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_4115;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_4265;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4105;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_4612;
wire n_3038;
wire n_2033;
wire n_3086;
wire n_4104;
wire n_4353;
wire n_2531;
wire n_1789;
wire n_1770;
wire n_4787;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_2071;
wire n_1144;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_4779;
wire n_4640;
wire n_3521;
wire n_3233;
wire n_4599;
wire n_2800;
wire n_1710;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_2805;
wire n_1301;
wire n_4769;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_4628;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_4784;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_4594;
wire n_1998;
wire n_3066;
wire n_4727;
wire n_3101;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_1574;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_3374;
wire n_1194;
wire n_4429;
wire n_4538;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4506;
wire n_2640;
wire n_3695;
wire n_4642;
wire n_4051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_4684;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_4768;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_4758;
wire n_4781;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4522;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_1170;
wire n_2221;
wire n_1629;
wire n_4263;
wire n_2055;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_3017;
wire n_1632;
wire n_1890;
wire n_3955;
wire n_2477;
wire n_1805;
wire n_2280;
wire n_1888;
wire n_1557;
wire n_3903;
wire n_3945;
wire n_1833;
wire n_1311;
wire n_4780;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_4803;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_4750;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_4648;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_3274;
wire n_2899;
wire n_3333;
wire n_4129;
wire n_3186;
wire n_1322;
wire n_4457;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_4804;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_4794;
wire n_4500;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1423;
wire n_1935;
wire n_4039;
wire n_4745;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_1801;
wire n_4426;
wire n_2912;
wire n_4703;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_4762;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_4030;
wire n_1612;
wire n_1240;
wire n_4809;

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_426),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1011),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1045),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_284),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_1031),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_87),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_424),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_997),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1021),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_358),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_426),
.Y(n_1086)
);

CKINVDCx16_ASAP7_75t_R g1087 ( 
.A(n_658),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_289),
.Y(n_1088)
);

CKINVDCx16_ASAP7_75t_R g1089 ( 
.A(n_998),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_526),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_513),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_314),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_510),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_409),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_88),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_360),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_169),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_858),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_859),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_628),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_374),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1050),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_124),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_749),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_913),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_203),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_874),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_257),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_857),
.Y(n_1110)
);

BUFx10_ASAP7_75t_L g1111 ( 
.A(n_292),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_182),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_886),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_909),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_742),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_935),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_685),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_886),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_338),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_34),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_745),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_277),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_500),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_718),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_683),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_949),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_905),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_299),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_835),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_176),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_911),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_56),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_892),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_958),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_896),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_539),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_199),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_646),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_39),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_277),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_606),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_563),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1012),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_217),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_49),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_482),
.Y(n_1146)
);

CKINVDCx14_ASAP7_75t_R g1147 ( 
.A(n_484),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_451),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_970),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_37),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_861),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_934),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_923),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_729),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_314),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_396),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_21),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_397),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_646),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_599),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1039),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_480),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_415),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_670),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_895),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_712),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_821),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_20),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_817),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_265),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_178),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_172),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_435),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_917),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_815),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_140),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_381),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_831),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_60),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_164),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_76),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_719),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_947),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_921),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_478),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_513),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_965),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_768),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_863),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_405),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_665),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_639),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_379),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_178),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_323),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_824),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_834),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_508),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_406),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_32),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_233),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_99),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_463),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_211),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_425),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_712),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_606),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_512),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_902),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_833),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_675),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_809),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_729),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_936),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_547),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_910),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_500),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_772),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_924),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1032),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_859),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_939),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_80),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_365),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_168),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_905),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_954),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_865),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1006),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_832),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_924),
.Y(n_1231)
);

BUFx5_ASAP7_75t_L g1232 ( 
.A(n_80),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_652),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_599),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_691),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_811),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_267),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1022),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_935),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_273),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_878),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_560),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_284),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_983),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_390),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_747),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_830),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_579),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_901),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_947),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_454),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_129),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_190),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1028),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_860),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_49),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_985),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_839),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1052),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_237),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_615),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_382),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_536),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_285),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_862),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_768),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_845),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_785),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_538),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_395),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_991),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_953),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_456),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_458),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_43),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1040),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_442),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_175),
.Y(n_1278)
);

BUFx8_ASAP7_75t_SL g1279 ( 
.A(n_780),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_697),
.Y(n_1280)
);

CKINVDCx14_ASAP7_75t_R g1281 ( 
.A(n_960),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_476),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_308),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_717),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_53),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_601),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_584),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_622),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_872),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_763),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_816),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_2),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_294),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_219),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_475),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_818),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_899),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_230),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_644),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_307),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_2),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1068),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_519),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_20),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_765),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_628),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_645),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_669),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_691),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_746),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_183),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_440),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_922),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_419),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_108),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_586),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_798),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_589),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_805),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_420),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_373),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_32),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_94),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_454),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_660),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_91),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_194),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_772),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_849),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1014),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_911),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_981),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_488),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1024),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_683),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_614),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_142),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1043),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_364),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_828),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_773),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_908),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_518),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_863),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_121),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_842),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_381),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_528),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_932),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_390),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_906),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_81),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_316),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1057),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_840),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_556),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_218),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_491),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_673),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_915),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_77),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_898),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_36),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_190),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_512),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1019),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_687),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_527),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_798),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1038),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_506),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_995),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_938),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_367),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_661),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_118),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_928),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_182),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_346),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_896),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_801),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_554),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_703),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_898),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_376),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_550),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_276),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_856),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_509),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_51),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_251),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_658),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_585),
.Y(n_1393)
);

BUFx10_ASAP7_75t_L g1394 ( 
.A(n_582),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_814),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_684),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_161),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_822),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_942),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_806),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_595),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_523),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_992),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_31),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_31),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_239),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_35),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_463),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_403),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_959),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_67),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_697),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_289),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_45),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_341),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_290),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_65),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1062),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_328),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_707),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_78),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_808),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_550),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_495),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_301),
.Y(n_1425)
);

BUFx10_ASAP7_75t_L g1426 ( 
.A(n_351),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1025),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_903),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_633),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_220),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_504),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_932),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_138),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_889),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_506),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_583),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_25),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_746),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_829),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_605),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_846),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_199),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_74),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_645),
.Y(n_1444)
);

BUFx5_ASAP7_75t_L g1445 ( 
.A(n_319),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_292),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_107),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_741),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_713),
.Y(n_1449)
);

BUFx8_ASAP7_75t_SL g1450 ( 
.A(n_810),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1074),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_893),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_881),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_833),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_61),
.Y(n_1455)
);

CKINVDCx14_ASAP7_75t_R g1456 ( 
.A(n_625),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_384),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1023),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_945),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_65),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_14),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_858),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_955),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_78),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_831),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_100),
.Y(n_1466)
);

CKINVDCx14_ASAP7_75t_R g1467 ( 
.A(n_780),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_731),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_389),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_48),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_724),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_586),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_579),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_107),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_276),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_505),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_995),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_518),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_251),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_722),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_322),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_871),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_867),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_623),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_922),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_102),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_418),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_680),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_392),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_198),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_722),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_648),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_718),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_944),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_417),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_654),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_231),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_425),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_555),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_536),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_715),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_919),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_975),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_70),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_428),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_44),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_4),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1066),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_54),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_891),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_657),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_10),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_943),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1009),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_408),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_213),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_914),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_926),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_112),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_567),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_323),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_904),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_899),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_322),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_241),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_158),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_167),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_814),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_527),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_113),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_782),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_274),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_358),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_420),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_83),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_829),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_805),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_907),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_836),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_551),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_502),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_626),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_524),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_221),
.Y(n_1544)
);

INVx4_ASAP7_75t_R g1545 ( 
.A(n_795),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_126),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_79),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_751),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1001),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_619),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_775),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_159),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_694),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_892),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_929),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_762),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_933),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_950),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_312),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_996),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_501),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_843),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_91),
.Y(n_1563)
);

INVxp33_ASAP7_75t_SL g1564 ( 
.A(n_801),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_603),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_187),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_344),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_273),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_443),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_629),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_197),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_979),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_137),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_912),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_631),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_53),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_720),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1059),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1004),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1060),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_799),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_738),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_397),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_779),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_350),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_528),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_160),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_883),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_641),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_409),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_480),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_979),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1073),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1056),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_897),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_531),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_813),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_644),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_437),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_941),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_442),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_298),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_350),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_103),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_548),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_796),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_622),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_209),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_68),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_839),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_515),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_825),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_170),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_10),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_473),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_526),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_71),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_192),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_260),
.Y(n_1619)
);

CKINVDCx12_ASAP7_75t_R g1620 ( 
.A(n_462),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_256),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_562),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_181),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_493),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_465),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_461),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_867),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_607),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_879),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_168),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_854),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_161),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_786),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1055),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_651),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_838),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_127),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_271),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_890),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_866),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_467),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_525),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_666),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_445),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_663),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_462),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_855),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_517),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_197),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_882),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_538),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_850),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_278),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_885),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_248),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_537),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_419),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_546),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_601),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_930),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_657),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_460),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_771),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_54),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_594),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_353),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_852),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_417),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_823),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_386),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_7),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_248),
.Y(n_1672)
);

CKINVDCx20_ASAP7_75t_R g1673 ( 
.A(n_451),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_488),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_321),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_220),
.Y(n_1676)
);

CKINVDCx14_ASAP7_75t_R g1677 ( 
.A(n_73),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_799),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_844),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_187),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_853),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_715),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_202),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_970),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_551),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_468),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_802),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_837),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_423),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_384),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_709),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_469),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_5),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_669),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_47),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_972),
.Y(n_1696)
);

BUFx2_ASAP7_75t_SL g1697 ( 
.A(n_940),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_807),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_840),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1015),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_755),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_482),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_760),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_57),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_471),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_304),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_448),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_478),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_948),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_894),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_395),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_826),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_705),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_936),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_687),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_954),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_240),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_664),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_50),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_195),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_969),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_880),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_163),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_389),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_808),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_937),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_887),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_183),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_430),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_957),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_75),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_423),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_504),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_252),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_468),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_714),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_589),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_137),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_888),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_786),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_703),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_705),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_521),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_14),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_15),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_418),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_812),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_414),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_673),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_118),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1070),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_887),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_169),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_796),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_819),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_355),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_92),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_827),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_965),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_272),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_714),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1046),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_453),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_869),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_310),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_166),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_215),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_690),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_902),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_916),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_906),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_720),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_201),
.Y(n_1773)
);

CKINVDCx14_ASAP7_75t_R g1774 ( 
.A(n_213),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_209),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_207),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_771),
.Y(n_1777)
);

BUFx2_ASAP7_75t_SL g1778 ( 
.A(n_115),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_285),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_516),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_634),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_918),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_643),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_764),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_448),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_219),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_138),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_486),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_67),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1017),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_956),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_354),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_619),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_820),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_87),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_553),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_926),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_827),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_268),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_263),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_415),
.Y(n_1801)
);

BUFx5_ASAP7_75t_L g1802 ( 
.A(n_618),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_850),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_424),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_242),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_745),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_416),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_841),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_73),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_822),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_223),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_372),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_626),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_664),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_510),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_834),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_640),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_367),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_736),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_868),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_39),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_921),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_647),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_335),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_127),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_150),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_951),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_875),
.Y(n_1828)
);

BUFx10_ASAP7_75t_L g1829 ( 
.A(n_976),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_443),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_894),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_176),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_191),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_126),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_946),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_931),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_309),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_877),
.Y(n_1838)
);

BUFx10_ASAP7_75t_L g1839 ( 
.A(n_469),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_223),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1051),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_761),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_348),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_851),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1036),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_660),
.Y(n_1846)
);

BUFx5_ASAP7_75t_L g1847 ( 
.A(n_791),
.Y(n_1847)
);

CKINVDCx20_ASAP7_75t_R g1848 ( 
.A(n_884),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_904),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_699),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_930),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_143),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_609),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_802),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_254),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_218),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_432),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_252),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_108),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_943),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_962),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_145),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_938),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_100),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_109),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_370),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1030),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_784),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_460),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_346),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_848),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_555),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_681),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_925),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_686),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_572),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_641),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_422),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_361),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_876),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_436),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_927),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_869),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_591),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_19),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_193),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_583),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_517),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_620),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_881),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_484),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_900),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_133),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_883),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_485),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_865),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_920),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_45),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_345),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_882),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_269),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_682),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_885),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_678),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_256),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_809),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_923),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_778),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_873),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_334),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_847),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_952),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_870),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_994),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_243),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_490),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_987),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_577),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_109),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_744),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_946),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_400),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_949),
.Y(n_1923)
);

CKINVDCx20_ASAP7_75t_R g1924 ( 
.A(n_637),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_184),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_505),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_375),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_111),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_486),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_873),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_271),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_864),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_591),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_139),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_570),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_211),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1232),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1232),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1620),
.Y(n_1939)
);

INVxp33_ASAP7_75t_SL g1940 ( 
.A(n_1106),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1232),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1279),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1084),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1232),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1279),
.Y(n_1945)
);

CKINVDCx20_ASAP7_75t_R g1946 ( 
.A(n_1083),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1083),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1450),
.Y(n_1948)
);

CKINVDCx20_ASAP7_75t_R g1949 ( 
.A(n_1508),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1232),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1077),
.Y(n_1951)
);

CKINVDCx20_ASAP7_75t_R g1952 ( 
.A(n_1508),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1232),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1450),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1129),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1265),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1232),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1445),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1445),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1080),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1445),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1445),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1169),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1287),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1549),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1169),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1445),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1445),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1445),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1802),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1102),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1802),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1349),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1802),
.Y(n_1974)
);

CKINVDCx14_ASAP7_75t_R g1975 ( 
.A(n_1147),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1549),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1802),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1354),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1089),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1169),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1802),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1802),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1143),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1802),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1439),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1847),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1847),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1847),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1328),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1077),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1281),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1328),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1847),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1259),
.Y(n_1994)
);

CKINVDCx16_ASAP7_75t_R g1995 ( 
.A(n_1087),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1847),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1847),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1847),
.Y(n_1998)
);

CKINVDCx20_ASAP7_75t_R g1999 ( 
.A(n_1456),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1467),
.Y(n_2000)
);

CKINVDCx16_ASAP7_75t_R g2001 ( 
.A(n_1138),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1462),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1328),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1349),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1363),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1471),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1302),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1338),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1408),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1408),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1677),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1408),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1880),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1748),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1514),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1880),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1578),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1579),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1880),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1774),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1181),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_1580),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1181),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1224),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1224),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1257),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1593),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1257),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1332),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1428),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1349),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1349),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1298),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1354),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1298),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1470),
.Y(n_2036)
);

INVxp33_ASAP7_75t_SL g2037 ( 
.A(n_1433),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1339),
.Y(n_2038)
);

CKINVDCx20_ASAP7_75t_R g2039 ( 
.A(n_1594),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1339),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1388),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1388),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1393),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1393),
.Y(n_2044)
);

CKINVDCx20_ASAP7_75t_R g2045 ( 
.A(n_1634),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1473),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1473),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1483),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1483),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1489),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1489),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1534),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1470),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1526),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1790),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1470),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1534),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1566),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_1841),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1566),
.Y(n_2060)
);

INVxp33_ASAP7_75t_L g2061 ( 
.A(n_1540),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1161),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1470),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1427),
.B(n_1404),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1607),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1486),
.Y(n_2066)
);

CKINVDCx16_ASAP7_75t_R g2067 ( 
.A(n_1111),
.Y(n_2067)
);

INVxp67_ASAP7_75t_SL g2068 ( 
.A(n_1613),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1607),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1081),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1649),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_1649),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1763),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1662),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1763),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1883),
.Y(n_2076)
);

INVxp33_ASAP7_75t_L g2077 ( 
.A(n_1835),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1883),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1486),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1486),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1486),
.Y(n_2081)
);

INVxp33_ASAP7_75t_SL g2082 ( 
.A(n_1899),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1511),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1511),
.Y(n_2084)
);

INVxp67_ASAP7_75t_SL g2085 ( 
.A(n_1936),
.Y(n_2085)
);

CKINVDCx20_ASAP7_75t_R g2086 ( 
.A(n_1161),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1511),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1925),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1511),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1517),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1517),
.Y(n_2091)
);

CKINVDCx14_ASAP7_75t_R g2092 ( 
.A(n_1849),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1517),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_1092),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1085),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1517),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1090),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1572),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_1897),
.B(n_0),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1572),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1572),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1572),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1585),
.Y(n_2103)
);

INVxp33_ASAP7_75t_SL g2104 ( 
.A(n_1931),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1585),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1585),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1585),
.Y(n_2107)
);

CKINVDCx16_ASAP7_75t_R g2108 ( 
.A(n_1111),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1091),
.Y(n_2109)
);

CKINVDCx20_ASAP7_75t_R g2110 ( 
.A(n_1092),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1654),
.Y(n_2111)
);

INVxp33_ASAP7_75t_SL g2112 ( 
.A(n_1934),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1654),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1654),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1111),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1654),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1681),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1681),
.Y(n_2118)
);

CKINVDCx14_ASAP7_75t_R g2119 ( 
.A(n_1174),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1681),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1681),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1682),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1682),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_1076),
.Y(n_2124)
);

CKINVDCx20_ASAP7_75t_R g2125 ( 
.A(n_1096),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1682),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1682),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1683),
.Y(n_2128)
);

CKINVDCx14_ASAP7_75t_R g2129 ( 
.A(n_1174),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1683),
.Y(n_2130)
);

INVxp67_ASAP7_75t_SL g2131 ( 
.A(n_1683),
.Y(n_2131)
);

INVxp33_ASAP7_75t_L g2132 ( 
.A(n_1079),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1683),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1076),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1978),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2131),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2004),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_L g2138 ( 
.A(n_1978),
.Y(n_2138)
);

BUFx8_ASAP7_75t_L g2139 ( 
.A(n_2115),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_2072),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2031),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2032),
.Y(n_2142)
);

CKINVDCx16_ASAP7_75t_R g2143 ( 
.A(n_1991),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2036),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2053),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2029),
.B(n_1078),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2056),
.Y(n_2147)
);

AND2x2_ASAP7_75t_SL g2148 ( 
.A(n_1995),
.B(n_1276),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2063),
.Y(n_2149)
);

OA21x2_ASAP7_75t_L g2150 ( 
.A1(n_2003),
.A2(n_1229),
.B(n_1220),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1960),
.B(n_1427),
.Y(n_2151)
);

AND2x6_ASAP7_75t_L g2152 ( 
.A(n_2021),
.B(n_1105),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1978),
.Y(n_2153)
);

AND2x2_ASAP7_75t_SL g2154 ( 
.A(n_2001),
.B(n_2099),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_1973),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1971),
.B(n_1276),
.Y(n_2156)
);

AND2x6_ASAP7_75t_L g2157 ( 
.A(n_2023),
.B(n_1159),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_2034),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_L g2159 ( 
.A1(n_1956),
.A2(n_1149),
.B1(n_1152),
.B2(n_1148),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1983),
.B(n_1366),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2030),
.B(n_1238),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_2070),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2066),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_2034),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2084),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2100),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_2034),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1973),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_2103),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_1951),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2088),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2107),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2121),
.Y(n_2173)
);

NAND2xp33_ASAP7_75t_L g2174 ( 
.A(n_2095),
.B(n_1740),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_2068),
.B(n_1254),
.Y(n_2175)
);

OA21x2_ASAP7_75t_L g2176 ( 
.A1(n_2009),
.A2(n_1334),
.B(n_1330),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_2133),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2079),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1994),
.B(n_1366),
.Y(n_2179)
);

INVx6_ASAP7_75t_L g2180 ( 
.A(n_2067),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1958),
.A2(n_1867),
.B(n_1418),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2080),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1990),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_2081),
.Y(n_2184)
);

AND2x6_ASAP7_75t_L g2185 ( 
.A(n_2024),
.B(n_1184),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2007),
.B(n_1867),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_SL g2187 ( 
.A1(n_2094),
.A2(n_1119),
.B1(n_1122),
.B2(n_1096),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2108),
.B(n_1740),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2083),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_2074),
.B(n_1370),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2087),
.Y(n_2191)
);

INVx3_ASAP7_75t_L g2192 ( 
.A(n_2089),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2022),
.B(n_1451),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_2097),
.B(n_1564),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2090),
.Y(n_2195)
);

OA21x2_ASAP7_75t_L g2196 ( 
.A1(n_2010),
.A2(n_1700),
.B(n_1458),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1975),
.B(n_1174),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2109),
.B(n_1292),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2005),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1940),
.A2(n_1406),
.B1(n_1531),
.B2(n_1135),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_2091),
.Y(n_2201)
);

INVx5_ASAP7_75t_L g2202 ( 
.A(n_1967),
.Y(n_2202)
);

CKINVDCx16_ASAP7_75t_R g2203 ( 
.A(n_1999),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2093),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2096),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2098),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2101),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2102),
.Y(n_2208)
);

BUFx12f_ASAP7_75t_L g2209 ( 
.A(n_1942),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2105),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_2039),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2106),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2085),
.B(n_1751),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2111),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2113),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_2114),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1943),
.B(n_1292),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2116),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2124),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_2117),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_2118),
.Y(n_2221)
);

INVx5_ASAP7_75t_L g2222 ( 
.A(n_1984),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2008),
.B(n_1762),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_2045),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2120),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1963),
.B(n_1292),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2122),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2123),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2126),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2127),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_2128),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2130),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1986),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1966),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_2059),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_2062),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1980),
.Y(n_2237)
);

BUFx8_ASAP7_75t_L g2238 ( 
.A(n_2025),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1989),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2026),
.Y(n_2240)
);

CKINVDCx6p67_ASAP7_75t_R g2241 ( 
.A(n_2000),
.Y(n_2241)
);

INVx4_ASAP7_75t_L g2242 ( 
.A(n_2015),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_2028),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_1997),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_2033),
.Y(n_2245)
);

AND2x6_ASAP7_75t_L g2246 ( 
.A(n_2035),
.B(n_1225),
.Y(n_2246)
);

BUFx3_ASAP7_75t_L g2247 ( 
.A(n_2038),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2092),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1937),
.Y(n_2249)
);

NAND2x1p5_ASAP7_75t_L g2250 ( 
.A(n_1956),
.B(n_1354),
.Y(n_2250)
);

BUFx3_ASAP7_75t_L g2251 ( 
.A(n_2040),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1992),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_1938),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1941),
.Y(n_2254)
);

BUFx12f_ASAP7_75t_L g2255 ( 
.A(n_1945),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2012),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1944),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2013),
.Y(n_2258)
);

CKINVDCx8_ASAP7_75t_R g2259 ( 
.A(n_1948),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_2119),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1955),
.B(n_1845),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2016),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1950),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2037),
.A2(n_1564),
.B1(n_1323),
.B2(n_1407),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1953),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_1957),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2017),
.B(n_1354),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2019),
.Y(n_2268)
);

OA21x2_ASAP7_75t_L g2269 ( 
.A1(n_2064),
.A2(n_1113),
.B(n_1088),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2082),
.A2(n_1560),
.B1(n_1547),
.B2(n_1149),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2041),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_2129),
.Y(n_2272)
);

BUFx8_ASAP7_75t_L g2273 ( 
.A(n_2042),
.Y(n_2273)
);

BUFx6f_ASAP7_75t_L g2274 ( 
.A(n_1959),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2043),
.Y(n_2275)
);

AOI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_1979),
.A2(n_1665),
.B1(n_1926),
.B2(n_1115),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1961),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1962),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2044),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1985),
.B(n_2002),
.Y(n_2280)
);

OA21x2_ASAP7_75t_L g2281 ( 
.A1(n_2064),
.A2(n_1113),
.B(n_1088),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2046),
.Y(n_2282)
);

OA21x2_ASAP7_75t_L g2283 ( 
.A1(n_1968),
.A2(n_1140),
.B(n_1139),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2047),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_2134),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2048),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1969),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1970),
.Y(n_2288)
);

BUFx8_ASAP7_75t_L g2289 ( 
.A(n_2049),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2006),
.B(n_1404),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2050),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2051),
.Y(n_2292)
);

CKINVDCx16_ASAP7_75t_R g2293 ( 
.A(n_2011),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2018),
.B(n_1740),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2052),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2057),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2027),
.B(n_1740),
.Y(n_2297)
);

BUFx3_ASAP7_75t_L g2298 ( 
.A(n_2058),
.Y(n_2298)
);

INVx4_ASAP7_75t_L g2299 ( 
.A(n_2055),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1972),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2060),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2065),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2069),
.B(n_1490),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_1974),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_2086),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2071),
.B(n_1490),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_L g2307 ( 
.A(n_1964),
.B(n_1148),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1977),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2061),
.B(n_1313),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2073),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2014),
.B(n_1612),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_1939),
.Y(n_2312)
);

AND2x6_ASAP7_75t_L g2313 ( 
.A(n_2075),
.B(n_1251),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_1954),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2020),
.A2(n_1095),
.B1(n_1099),
.B2(n_1094),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2076),
.B(n_2078),
.Y(n_2316)
);

OA21x2_ASAP7_75t_L g2317 ( 
.A1(n_1981),
.A2(n_1140),
.B(n_1139),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1982),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1987),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1988),
.Y(n_2320)
);

OAI21x1_ASAP7_75t_L g2321 ( 
.A1(n_1993),
.A2(n_1177),
.B(n_1163),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1996),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1998),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_2132),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2054),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2077),
.B(n_1313),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2104),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_1964),
.B(n_1612),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2112),
.B(n_1701),
.Y(n_2329)
);

AND2x4_ASAP7_75t_L g2330 ( 
.A(n_1946),
.B(n_1701),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_1947),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1949),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1952),
.Y(n_2333)
);

INVx2_ASAP7_75t_SL g2334 ( 
.A(n_2110),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1965),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_SL g2336 ( 
.A1(n_2125),
.A2(n_1122),
.B1(n_1126),
.B2(n_1119),
.Y(n_2336)
);

INVx6_ASAP7_75t_L g2337 ( 
.A(n_1976),
.Y(n_2337)
);

OAI21x1_ASAP7_75t_L g2338 ( 
.A1(n_1958),
.A2(n_1177),
.B(n_1163),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1960),
.B(n_1727),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2131),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2131),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1960),
.B(n_1727),
.Y(n_2342)
);

BUFx8_ASAP7_75t_SL g2343 ( 
.A(n_2094),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2004),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_2070),
.Y(n_2345)
);

OA21x2_ASAP7_75t_L g2346 ( 
.A1(n_2003),
.A2(n_1240),
.B(n_1190),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2131),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_2029),
.B(n_1768),
.Y(n_2348)
);

CKINVDCx11_ASAP7_75t_R g2349 ( 
.A(n_2094),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_1978),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2131),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_1978),
.Y(n_2352)
);

BUFx2_ASAP7_75t_L g2353 ( 
.A(n_2062),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_1940),
.A2(n_1154),
.B1(n_1155),
.B2(n_1152),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_1960),
.B(n_1768),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_2070),
.Y(n_2356)
);

OAI21x1_ASAP7_75t_L g2357 ( 
.A1(n_1958),
.A2(n_1240),
.B(n_1190),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_1975),
.B(n_1313),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_1975),
.B(n_1321),
.Y(n_2359)
);

BUFx3_ASAP7_75t_L g2360 ( 
.A(n_2072),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1978),
.Y(n_2361)
);

BUFx8_ASAP7_75t_L g2362 ( 
.A(n_2115),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1960),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2004),
.Y(n_2364)
);

INVx5_ASAP7_75t_L g2365 ( 
.A(n_1978),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2072),
.Y(n_2366)
);

AND2x2_ASAP7_75t_SL g2367 ( 
.A(n_1995),
.B(n_1252),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2004),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2004),
.Y(n_2369)
);

BUFx8_ASAP7_75t_L g2370 ( 
.A(n_2115),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2131),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2004),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_2072),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_1978),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2004),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_2062),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_1975),
.B(n_1321),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2131),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2131),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_1975),
.B(n_1321),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1960),
.B(n_1910),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_1975),
.B(n_1350),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2131),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2072),
.Y(n_2384)
);

XNOR2xp5_ASAP7_75t_L g2385 ( 
.A(n_1946),
.B(n_1126),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2131),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2029),
.B(n_1910),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2004),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_2029),
.B(n_1082),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2131),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2131),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2131),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2131),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2131),
.Y(n_2394)
);

BUFx6f_ASAP7_75t_L g2395 ( 
.A(n_1978),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_1940),
.A2(n_1155),
.B1(n_1157),
.B2(n_1154),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2072),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2131),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2072),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_1978),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2029),
.B(n_1086),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2072),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2131),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2131),
.Y(n_2404)
);

INVxp67_ASAP7_75t_L g2405 ( 
.A(n_2005),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1960),
.B(n_1100),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1960),
.B(n_1101),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_1975),
.B(n_1350),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2004),
.Y(n_2409)
);

BUFx8_ASAP7_75t_L g2410 ( 
.A(n_2115),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2131),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2131),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2131),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2070),
.B(n_1107),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1960),
.B(n_1108),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2131),
.Y(n_2416)
);

OA21x2_ASAP7_75t_L g2417 ( 
.A1(n_2003),
.A2(n_1260),
.B(n_1252),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2004),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2131),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2131),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2072),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2062),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1960),
.B(n_1109),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2004),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2131),
.Y(n_2425)
);

OA21x2_ASAP7_75t_L g2426 ( 
.A1(n_2003),
.A2(n_1271),
.B(n_1260),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2004),
.Y(n_2427)
);

BUFx8_ASAP7_75t_L g2428 ( 
.A(n_2115),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2062),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_1978),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2029),
.B(n_1093),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_1978),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2131),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2004),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1978),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_1995),
.B(n_1350),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_1978),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2131),
.Y(n_2438)
);

BUFx6f_ASAP7_75t_L g2439 ( 
.A(n_1978),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_2029),
.B(n_1097),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2131),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_1978),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2004),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2131),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_1978),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_1946),
.Y(n_2446)
);

NOR2x1_ASAP7_75t_L g2447 ( 
.A(n_2022),
.B(n_1098),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2070),
.B(n_1112),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2004),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_1995),
.B(n_1394),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2131),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_1978),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2070),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2131),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1960),
.B(n_1114),
.Y(n_2455)
);

AND2x6_ASAP7_75t_L g2456 ( 
.A(n_2021),
.B(n_1290),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2131),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_1960),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2004),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_1978),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2131),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2131),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2131),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2070),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_1960),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2004),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2131),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2004),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2004),
.Y(n_2469)
);

OAI21x1_ASAP7_75t_L g2470 ( 
.A1(n_1958),
.A2(n_1285),
.B(n_1271),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_1960),
.B(n_1116),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2072),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_1960),
.B(n_1120),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_1995),
.B(n_1394),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2004),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2004),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2267),
.B(n_1285),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2324),
.B(n_1394),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2271),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2363),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_2458),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2465),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2169),
.Y(n_2483)
);

BUFx2_ASAP7_75t_L g2484 ( 
.A(n_2324),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2343),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_R g2486 ( 
.A(n_2314),
.B(n_1121),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2169),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2349),
.Y(n_2488)
);

CKINVDCx5p33_ASAP7_75t_R g2489 ( 
.A(n_2241),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2135),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_2211),
.Y(n_2491)
);

INVx2_ASAP7_75t_SL g2492 ( 
.A(n_2198),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2224),
.Y(n_2493)
);

INVxp33_ASAP7_75t_L g2494 ( 
.A(n_2385),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2235),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2177),
.Y(n_2496)
);

AOI21x1_ASAP7_75t_L g2497 ( 
.A1(n_2319),
.A2(n_2277),
.B(n_2254),
.Y(n_2497)
);

CKINVDCx20_ASAP7_75t_R g2498 ( 
.A(n_2143),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2203),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2293),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2244),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2209),
.Y(n_2502)
);

INVxp33_ASAP7_75t_L g2503 ( 
.A(n_2309),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2255),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2170),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2242),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2326),
.B(n_1426),
.Y(n_2507)
);

AND3x1_ASAP7_75t_L g2508 ( 
.A(n_2264),
.B(n_1104),
.C(n_1103),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2275),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_R g2510 ( 
.A(n_2259),
.B(n_2174),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2177),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_2299),
.Y(n_2512)
);

CKINVDCx20_ASAP7_75t_R g2513 ( 
.A(n_2337),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2171),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2279),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2282),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2328),
.B(n_1426),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2453),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2367),
.A2(n_1352),
.B1(n_1364),
.B2(n_1322),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2464),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2248),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2244),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2284),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2331),
.Y(n_2524)
);

INVxp67_ASAP7_75t_L g2525 ( 
.A(n_2217),
.Y(n_2525)
);

CKINVDCx20_ASAP7_75t_R g2526 ( 
.A(n_2236),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2135),
.Y(n_2527)
);

CKINVDCx20_ASAP7_75t_R g2528 ( 
.A(n_2305),
.Y(n_2528)
);

CKINVDCx20_ASAP7_75t_R g2529 ( 
.A(n_2353),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_2331),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2162),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2345),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2356),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2376),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2151),
.B(n_1123),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2138),
.Y(n_2536)
);

CKINVDCx16_ASAP7_75t_R g2537 ( 
.A(n_2260),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2184),
.Y(n_2538)
);

NOR2xp67_ASAP7_75t_L g2539 ( 
.A(n_2272),
.B(n_999),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2422),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2184),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2292),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2295),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_2414),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2296),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2301),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2302),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2429),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2140),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2446),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2366),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2139),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_2362),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2370),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2384),
.Y(n_2555)
);

NAND2xp33_ASAP7_75t_SL g2556 ( 
.A(n_2219),
.B(n_1136),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2360),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2201),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2410),
.Y(n_2559)
);

INVxp67_ASAP7_75t_L g2560 ( 
.A(n_2448),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2428),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2294),
.B(n_1358),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2180),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2373),
.Y(n_2564)
);

CKINVDCx20_ASAP7_75t_R g2565 ( 
.A(n_2334),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2201),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2297),
.B(n_1358),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2310),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2212),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_2406),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2407),
.Y(n_2571)
);

HB1xp67_ASAP7_75t_L g2572 ( 
.A(n_2397),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2415),
.Y(n_2573)
);

AOI21x1_ASAP7_75t_L g2574 ( 
.A1(n_2288),
.A2(n_1117),
.B(n_1110),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2423),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2455),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2471),
.Y(n_2577)
);

CKINVDCx20_ASAP7_75t_R g2578 ( 
.A(n_2332),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2473),
.Y(n_2579)
);

XOR2xp5_ASAP7_75t_L g2580 ( 
.A(n_2333),
.B(n_1136),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2249),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2194),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2212),
.Y(n_2583)
);

CKINVDCx20_ASAP7_75t_R g2584 ( 
.A(n_2335),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2183),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2249),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_2148),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2327),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2156),
.Y(n_2589)
);

INVxp67_ASAP7_75t_SL g2590 ( 
.A(n_2399),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2253),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2253),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2160),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2257),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2179),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2216),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2186),
.Y(n_2597)
);

CKINVDCx20_ASAP7_75t_R g2598 ( 
.A(n_2315),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2402),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2421),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_2472),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2216),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2257),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2223),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2263),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_2154),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2339),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2342),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2355),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2381),
.Y(n_2610)
);

NOR2xp67_ASAP7_75t_L g2611 ( 
.A(n_2285),
.B(n_1000),
.Y(n_2611)
);

BUFx10_ASAP7_75t_L g2612 ( 
.A(n_2280),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2263),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2265),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2187),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2336),
.Y(n_2616)
);

CKINVDCx16_ASAP7_75t_R g2617 ( 
.A(n_2197),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2234),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2237),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_R g2620 ( 
.A(n_2136),
.B(n_1124),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2239),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2221),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2265),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2252),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2243),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2138),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2221),
.Y(n_2627)
);

INVxp67_ASAP7_75t_L g2628 ( 
.A(n_2307),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2245),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2266),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_R g2631 ( 
.A(n_2340),
.B(n_1125),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2341),
.B(n_1376),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2247),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2251),
.Y(n_2634)
);

CKINVDCx20_ASAP7_75t_R g2635 ( 
.A(n_2276),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_2286),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2266),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2298),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2358),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2347),
.B(n_1127),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_2359),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2377),
.Y(n_2642)
);

OAI21x1_ASAP7_75t_L g2643 ( 
.A1(n_2338),
.A2(n_1434),
.B(n_1376),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_2380),
.Y(n_2644)
);

HB1xp67_ASAP7_75t_L g2645 ( 
.A(n_2250),
.Y(n_2645)
);

CKINVDCx20_ASAP7_75t_R g2646 ( 
.A(n_2199),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2274),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2274),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2226),
.B(n_2382),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2278),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_R g2651 ( 
.A(n_2351),
.B(n_1128),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2408),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2278),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2287),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2287),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2405),
.Y(n_2656)
);

CKINVDCx20_ASAP7_75t_R g2657 ( 
.A(n_2436),
.Y(n_2657)
);

CKINVDCx20_ASAP7_75t_R g2658 ( 
.A(n_2450),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2312),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2231),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2330),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2231),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_2354),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2329),
.B(n_1426),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2348),
.B(n_1565),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_2396),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2188),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2371),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2300),
.Y(n_2669)
);

BUFx2_ASAP7_75t_L g2670 ( 
.A(n_2152),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_R g2671 ( 
.A(n_2378),
.B(n_1130),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2325),
.B(n_2379),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2137),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2300),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2383),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_2386),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2153),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2304),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2390),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2141),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2391),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_R g2682 ( 
.A(n_2392),
.B(n_1131),
.Y(n_2682)
);

BUFx10_ASAP7_75t_L g2683 ( 
.A(n_2290),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_2393),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2394),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2398),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2403),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2304),
.Y(n_2688)
);

AOI21x1_ASAP7_75t_L g2689 ( 
.A1(n_2308),
.A2(n_1145),
.B(n_1118),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2404),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2318),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2318),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2142),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2411),
.Y(n_2694)
);

OAI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2200),
.A2(n_1443),
.B1(n_1510),
.B2(n_1403),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2320),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2320),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2144),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_2412),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2283),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_R g2701 ( 
.A(n_2413),
.B(n_1132),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2416),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_R g2703 ( 
.A(n_2419),
.B(n_1133),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_R g2704 ( 
.A(n_2420),
.B(n_1134),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2317),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2425),
.B(n_1434),
.Y(n_2706)
);

CKINVDCx20_ASAP7_75t_R g2707 ( 
.A(n_2474),
.Y(n_2707)
);

HB1xp67_ASAP7_75t_L g2708 ( 
.A(n_2155),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_2433),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2438),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2441),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2444),
.Y(n_2712)
);

HB1xp67_ASAP7_75t_L g2713 ( 
.A(n_2168),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_R g2714 ( 
.A(n_2451),
.B(n_1137),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_2454),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2457),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2322),
.Y(n_2717)
);

CKINVDCx20_ASAP7_75t_R g2718 ( 
.A(n_2238),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2461),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2462),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2323),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2463),
.B(n_1522),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2467),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2256),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2147),
.Y(n_2725)
);

CKINVDCx16_ASAP7_75t_R g2726 ( 
.A(n_2447),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2163),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_2146),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2161),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2269),
.Y(n_2730)
);

NOR2xp67_ASAP7_75t_L g2731 ( 
.A(n_2202),
.B(n_1002),
.Y(n_2731)
);

CKINVDCx16_ASAP7_75t_R g2732 ( 
.A(n_2193),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2175),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2258),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2262),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2166),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2172),
.Y(n_2737)
);

CKINVDCx20_ASAP7_75t_R g2738 ( 
.A(n_2273),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2190),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2213),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2289),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2387),
.Y(n_2742)
);

CKINVDCx20_ASAP7_75t_R g2743 ( 
.A(n_2270),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2152),
.Y(n_2744)
);

NAND2xp33_ASAP7_75t_R g2745 ( 
.A(n_2389),
.B(n_1157),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2157),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2233),
.B(n_1522),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2344),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2268),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2281),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2182),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2157),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2185),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_SL g2754 ( 
.A1(n_2159),
.A2(n_1178),
.B1(n_1182),
.B2(n_1151),
.Y(n_2754)
);

CKINVDCx20_ASAP7_75t_R g2755 ( 
.A(n_2316),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2189),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2185),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2364),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2246),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2246),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2313),
.Y(n_2761)
);

INVxp67_ASAP7_75t_L g2762 ( 
.A(n_2313),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2456),
.Y(n_2763)
);

BUFx10_ASAP7_75t_L g2764 ( 
.A(n_2311),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2401),
.B(n_1141),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_R g2766 ( 
.A(n_2240),
.B(n_1142),
.Y(n_2766)
);

HB1xp67_ASAP7_75t_L g2767 ( 
.A(n_2291),
.Y(n_2767)
);

CKINVDCx20_ASAP7_75t_R g2768 ( 
.A(n_2303),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2456),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2431),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2440),
.Y(n_2771)
);

CKINVDCx20_ASAP7_75t_R g2772 ( 
.A(n_2306),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2261),
.B(n_1565),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2195),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2206),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2368),
.B(n_1527),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2153),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2158),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2158),
.Y(n_2779)
);

HB1xp67_ASAP7_75t_L g2780 ( 
.A(n_2192),
.Y(n_2780)
);

NOR2xp33_ASAP7_75t_L g2781 ( 
.A(n_2218),
.B(n_1144),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2164),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2369),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_2164),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2497),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2777),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2673),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2484),
.B(n_2505),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2480),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2604),
.B(n_2150),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2544),
.B(n_1548),
.Y(n_2791)
);

BUFx6f_ASAP7_75t_L g2792 ( 
.A(n_2490),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2589),
.B(n_2176),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2507),
.B(n_1565),
.Y(n_2794)
);

BUFx6f_ASAP7_75t_L g2795 ( 
.A(n_2490),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2593),
.B(n_2196),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2724),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2734),
.Y(n_2798)
);

AND2x6_ASAP7_75t_L g2799 ( 
.A(n_2730),
.B(n_1527),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2680),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2560),
.B(n_1551),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2595),
.B(n_2346),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2735),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2597),
.B(n_1592),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2481),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2749),
.Y(n_2806)
);

AND2x4_ASAP7_75t_L g2807 ( 
.A(n_2601),
.B(n_2228),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2570),
.B(n_2417),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2693),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2698),
.Y(n_2810)
);

NAND2x1_ASAP7_75t_L g2811 ( 
.A(n_2700),
.B(n_2426),
.Y(n_2811)
);

AND2x6_ASAP7_75t_L g2812 ( 
.A(n_2750),
.B(n_1532),
.Y(n_2812)
);

CKINVDCx16_ASAP7_75t_R g2813 ( 
.A(n_2537),
.Y(n_2813)
);

BUFx4f_ASAP7_75t_L g2814 ( 
.A(n_2670),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2725),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2607),
.B(n_2608),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2550),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2571),
.B(n_2202),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2609),
.B(n_2167),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2610),
.B(n_1630),
.Y(n_2820)
);

NAND2x1p5_ASAP7_75t_L g2821 ( 
.A(n_2557),
.B(n_2321),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2503),
.B(n_1829),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2490),
.Y(n_2823)
);

INVxp67_ASAP7_75t_SL g2824 ( 
.A(n_2501),
.Y(n_2824)
);

OR2x6_ASAP7_75t_L g2825 ( 
.A(n_2521),
.B(n_1294),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2527),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2573),
.B(n_1657),
.Y(n_2827)
);

XNOR2xp5_ASAP7_75t_L g2828 ( 
.A(n_2498),
.B(n_2499),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2527),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2727),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2575),
.B(n_1666),
.Y(n_2831)
);

AO22x2_ASAP7_75t_L g2832 ( 
.A1(n_2580),
.A2(n_1697),
.B1(n_1778),
.B2(n_1387),
.Y(n_2832)
);

BUFx10_ASAP7_75t_L g2833 ( 
.A(n_2485),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2576),
.B(n_1729),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2577),
.B(n_2222),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2479),
.Y(n_2836)
);

OR2x2_ASAP7_75t_L g2837 ( 
.A(n_2525),
.B(n_1742),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2579),
.B(n_2222),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2509),
.Y(n_2839)
);

AND2x6_ASAP7_75t_L g2840 ( 
.A(n_2705),
.B(n_1532),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2535),
.B(n_2372),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2649),
.B(n_2167),
.Y(n_2842)
);

INVx1_ASAP7_75t_SL g2843 ( 
.A(n_2478),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2517),
.B(n_1829),
.Y(n_2844)
);

AND2x6_ASAP7_75t_L g2845 ( 
.A(n_2773),
.B(n_1546),
.Y(n_2845)
);

INVx3_ASAP7_75t_L g2846 ( 
.A(n_2527),
.Y(n_2846)
);

AND2x6_ASAP7_75t_L g2847 ( 
.A(n_2562),
.B(n_1546),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2582),
.B(n_1743),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2515),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2513),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2516),
.Y(n_2851)
);

BUFx6f_ASAP7_75t_L g2852 ( 
.A(n_2778),
.Y(n_2852)
);

OR2x2_ASAP7_75t_L g2853 ( 
.A(n_2525),
.B(n_1753),
.Y(n_2853)
);

INVx5_ASAP7_75t_L g2854 ( 
.A(n_2612),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2477),
.B(n_2375),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2618),
.B(n_2350),
.Y(n_2856)
);

BUFx6f_ASAP7_75t_L g2857 ( 
.A(n_2779),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2523),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2482),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2736),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2619),
.B(n_2350),
.Y(n_2861)
);

INVx3_ASAP7_75t_L g2862 ( 
.A(n_2483),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2646),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2590),
.B(n_2538),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2628),
.A2(n_2229),
.B1(n_2191),
.B2(n_2204),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2782),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2621),
.B(n_2352),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2542),
.Y(n_2868)
);

INVx3_ASAP7_75t_L g2869 ( 
.A(n_2487),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2543),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2784),
.Y(n_2871)
);

AOI21x1_ASAP7_75t_L g2872 ( 
.A1(n_2567),
.A2(n_2470),
.B(n_2357),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2545),
.Y(n_2873)
);

BUFx4f_ASAP7_75t_L g2874 ( 
.A(n_2492),
.Y(n_2874)
);

INVx4_ASAP7_75t_L g2875 ( 
.A(n_2563),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2737),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2624),
.B(n_2742),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2683),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2546),
.Y(n_2879)
);

AND2x2_ASAP7_75t_SL g2880 ( 
.A(n_2726),
.B(n_1550),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2547),
.Y(n_2881)
);

BUFx3_ASAP7_75t_L g2882 ( 
.A(n_2524),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2568),
.Y(n_2883)
);

INVx1_ASAP7_75t_SL g2884 ( 
.A(n_2755),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2667),
.A2(n_1901),
.B1(n_1922),
.B2(n_1887),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2748),
.Y(n_2886)
);

INVx3_ASAP7_75t_L g2887 ( 
.A(n_2496),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2758),
.Y(n_2888)
);

INVx4_ASAP7_75t_L g2889 ( 
.A(n_2530),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2668),
.B(n_2352),
.Y(n_2890)
);

INVx6_ASAP7_75t_L g2891 ( 
.A(n_2612),
.Y(n_2891)
);

BUFx6f_ASAP7_75t_L g2892 ( 
.A(n_2536),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2783),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2751),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2717),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2541),
.B(n_2145),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2675),
.B(n_1146),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2756),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2676),
.B(n_2679),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2774),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2721),
.Y(n_2901)
);

INVx3_ASAP7_75t_L g2902 ( 
.A(n_2511),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2775),
.B(n_2388),
.Y(n_2903)
);

AND2x6_ASAP7_75t_L g2904 ( 
.A(n_2765),
.B(n_2519),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2681),
.B(n_2409),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2672),
.B(n_1158),
.Y(n_2906)
);

BUFx6f_ASAP7_75t_L g2907 ( 
.A(n_2536),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2712),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2640),
.A2(n_2706),
.B1(n_2722),
.B2(n_2632),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2708),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2684),
.B(n_2361),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2685),
.B(n_1829),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2713),
.Y(n_2913)
);

NAND2x1p5_ASAP7_75t_L g2914 ( 
.A(n_2501),
.B(n_2361),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2780),
.Y(n_2915)
);

INVxp67_ASAP7_75t_L g2916 ( 
.A(n_2745),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2587),
.A2(n_2205),
.B1(n_2207),
.B2(n_2178),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2776),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2564),
.Y(n_2919)
);

INVx3_ASAP7_75t_L g2920 ( 
.A(n_2626),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2767),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2522),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2686),
.B(n_2418),
.Y(n_2923)
);

OR2x2_ASAP7_75t_L g2924 ( 
.A(n_2732),
.B(n_2656),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2747),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2643),
.Y(n_2926)
);

BUFx2_ASAP7_75t_L g2927 ( 
.A(n_2526),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2574),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2558),
.B(n_2149),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2687),
.B(n_2424),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2689),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2626),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2690),
.B(n_2694),
.Y(n_2933)
);

AND2x2_ASAP7_75t_SL g2934 ( 
.A(n_2508),
.B(n_1550),
.Y(n_2934)
);

AO22x2_ASAP7_75t_L g2935 ( 
.A1(n_2754),
.A2(n_1656),
.B1(n_1661),
.B2(n_1556),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2528),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2695),
.A2(n_1656),
.B1(n_1661),
.B2(n_1556),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2677),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2683),
.Y(n_2939)
);

INVx4_ASAP7_75t_SL g2940 ( 
.A(n_2581),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2677),
.Y(n_2941)
);

INVx4_ASAP7_75t_L g2942 ( 
.A(n_2585),
.Y(n_2942)
);

NOR2xp33_ASAP7_75t_L g2943 ( 
.A(n_2699),
.B(n_1170),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_2506),
.Y(n_2944)
);

INVx3_ASAP7_75t_R g2945 ( 
.A(n_2566),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2702),
.B(n_2374),
.Y(n_2946)
);

INVx1_ASAP7_75t_SL g2947 ( 
.A(n_2529),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2569),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2583),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2709),
.A2(n_1680),
.B1(n_1714),
.B2(n_1663),
.Y(n_2950)
);

INVx1_ASAP7_75t_SL g2951 ( 
.A(n_2534),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2710),
.B(n_1839),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2711),
.B(n_2374),
.Y(n_2953)
);

BUFx10_ASAP7_75t_L g2954 ( 
.A(n_2488),
.Y(n_2954)
);

INVx3_ASAP7_75t_L g2955 ( 
.A(n_2596),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2602),
.Y(n_2956)
);

INVxp67_ASAP7_75t_L g2957 ( 
.A(n_2556),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2622),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_SL g2959 ( 
.A(n_2531),
.B(n_2532),
.Y(n_2959)
);

INVxp33_ASAP7_75t_L g2960 ( 
.A(n_2486),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2627),
.Y(n_2961)
);

INVx5_ASAP7_75t_L g2962 ( 
.A(n_2764),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2660),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_SL g2964 ( 
.A(n_2764),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2715),
.B(n_1171),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2662),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2549),
.B(n_2165),
.Y(n_2967)
);

BUFx6f_ASAP7_75t_L g2968 ( 
.A(n_2599),
.Y(n_2968)
);

BUFx4f_ASAP7_75t_L g2969 ( 
.A(n_2586),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2591),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2716),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2592),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2719),
.Y(n_2973)
);

INVx8_ASAP7_75t_L g2974 ( 
.A(n_2500),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2720),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2723),
.Y(n_2976)
);

OR2x6_ASAP7_75t_L g2977 ( 
.A(n_2645),
.B(n_1663),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2551),
.Y(n_2978)
);

INVx4_ASAP7_75t_L g2979 ( 
.A(n_2600),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2661),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2594),
.B(n_2427),
.Y(n_2981)
);

NAND3xp33_ASAP7_75t_L g2982 ( 
.A(n_2781),
.B(n_2762),
.C(n_2588),
.Y(n_2982)
);

INVx4_ASAP7_75t_L g2983 ( 
.A(n_2491),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_2512),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2603),
.Y(n_2985)
);

AND2x6_ASAP7_75t_L g2986 ( 
.A(n_2605),
.B(n_1680),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2613),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2555),
.Y(n_2988)
);

INVx3_ASAP7_75t_L g2989 ( 
.A(n_2625),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2572),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2629),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2614),
.B(n_2434),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2623),
.Y(n_2993)
);

BUFx6f_ASAP7_75t_L g2994 ( 
.A(n_2493),
.Y(n_2994)
);

INVx4_ASAP7_75t_L g2995 ( 
.A(n_2495),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2630),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2728),
.A2(n_1173),
.B1(n_1175),
.B2(n_1172),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2637),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2664),
.A2(n_1786),
.B1(n_1787),
.B2(n_1714),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2647),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2648),
.B(n_2443),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2650),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2659),
.B(n_1176),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2653),
.B(n_2449),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2633),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2665),
.B(n_1179),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2654),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2634),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2584),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2533),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2655),
.B(n_2459),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2565),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2617),
.B(n_2395),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2669),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2636),
.B(n_1180),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2639),
.B(n_1839),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2638),
.B(n_1183),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2674),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2678),
.Y(n_3019)
);

CKINVDCx16_ASAP7_75t_R g3020 ( 
.A(n_2510),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2641),
.B(n_1839),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2688),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2642),
.B(n_2173),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2691),
.B(n_2466),
.Y(n_3024)
);

NAND2xp33_ASAP7_75t_SL g3025 ( 
.A(n_2744),
.B(n_1151),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2768),
.Y(n_3026)
);

BUFx4f_ASAP7_75t_L g3027 ( 
.A(n_2692),
.Y(n_3027)
);

NAND2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2539),
.B(n_2696),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_2697),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2611),
.B(n_2468),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_2489),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2620),
.B(n_2469),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_SL g3033 ( 
.A1(n_2884),
.A2(n_2616),
.B1(n_2615),
.B2(n_2635),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2785),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2918),
.B(n_2644),
.Y(n_3035)
);

AOI22xp33_ASAP7_75t_L g3036 ( 
.A1(n_2904),
.A2(n_2666),
.B1(n_2663),
.B2(n_2598),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2925),
.B(n_2652),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2797),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2804),
.B(n_2827),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2904),
.A2(n_2606),
.B1(n_2772),
.B2(n_2658),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2909),
.B(n_2729),
.Y(n_3041)
);

BUFx6f_ASAP7_75t_L g3042 ( 
.A(n_2792),
.Y(n_3042)
);

AO22x1_ASAP7_75t_L g3043 ( 
.A1(n_2848),
.A2(n_2752),
.B1(n_2753),
.B2(n_2746),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2808),
.A2(n_2739),
.B1(n_2740),
.B2(n_2733),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2787),
.Y(n_3045)
);

AOI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2904),
.A2(n_2707),
.B1(n_2657),
.B2(n_2514),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_2802),
.A2(n_2743),
.B1(n_2759),
.B2(n_2757),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2791),
.B(n_2770),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2831),
.B(n_2518),
.Y(n_3049)
);

BUFx6f_ASAP7_75t_L g3050 ( 
.A(n_2792),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2933),
.B(n_2520),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2899),
.B(n_2760),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2800),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2809),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2801),
.B(n_2771),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2810),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2815),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2798),
.Y(n_3058)
);

NOR3xp33_ASAP7_75t_L g3059 ( 
.A(n_2816),
.B(n_2763),
.C(n_2761),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_SL g3060 ( 
.A(n_2971),
.B(n_2769),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2834),
.B(n_2631),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2973),
.B(n_2651),
.Y(n_3062)
);

OR2x2_ASAP7_75t_L g3063 ( 
.A(n_2817),
.B(n_2494),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2830),
.Y(n_3064)
);

NAND2x1p5_ASAP7_75t_L g3065 ( 
.A(n_2852),
.B(n_2395),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2795),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2841),
.B(n_2671),
.Y(n_3067)
);

OAI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_2959),
.A2(n_2548),
.B1(n_2540),
.B2(n_2578),
.Y(n_3068)
);

INVx3_ASAP7_75t_L g3069 ( 
.A(n_2788),
.Y(n_3069)
);

INVx2_ASAP7_75t_SL g3070 ( 
.A(n_3023),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2820),
.B(n_2682),
.Y(n_3071)
);

INVx8_ASAP7_75t_L g3072 ( 
.A(n_2974),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2852),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_2882),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2860),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2916),
.B(n_2975),
.Y(n_3076)
);

INVx8_ASAP7_75t_L g3077 ( 
.A(n_2974),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2790),
.B(n_2701),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2793),
.B(n_2703),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2843),
.B(n_2704),
.Y(n_3080)
);

O2A1O1Ixp5_ASAP7_75t_L g3081 ( 
.A1(n_2796),
.A2(n_2476),
.B(n_2475),
.C(n_2210),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2880),
.B(n_2714),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2855),
.B(n_2766),
.Y(n_3083)
);

OR2x2_ASAP7_75t_L g3084 ( 
.A(n_2837),
.B(n_2502),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2960),
.B(n_2552),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2876),
.Y(n_3086)
);

NOR3xp33_ASAP7_75t_L g3087 ( 
.A(n_2877),
.B(n_2554),
.C(n_2553),
.Y(n_3087)
);

INVx2_ASAP7_75t_SL g3088 ( 
.A(n_2977),
.Y(n_3088)
);

INVx1_ASAP7_75t_SL g3089 ( 
.A(n_2863),
.Y(n_3089)
);

INVx4_ASAP7_75t_L g3090 ( 
.A(n_2857),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2811),
.A2(n_1182),
.B1(n_1192),
.B2(n_1178),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_L g3092 ( 
.A(n_3009),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2803),
.B(n_2208),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2806),
.B(n_2214),
.Y(n_3094)
);

INVxp67_ASAP7_75t_L g3095 ( 
.A(n_2822),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2836),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2839),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2799),
.A2(n_2812),
.B1(n_2851),
.B2(n_2849),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2858),
.B(n_2215),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2868),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2840),
.A2(n_2181),
.B1(n_1219),
.B2(n_1222),
.Y(n_3101)
);

OR2x2_ASAP7_75t_L g3102 ( 
.A(n_2853),
.B(n_2504),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2870),
.B(n_2225),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2873),
.B(n_2879),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2881),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2883),
.B(n_2230),
.Y(n_3106)
);

NAND2xp33_ASAP7_75t_L g3107 ( 
.A(n_2799),
.B(n_2559),
.Y(n_3107)
);

NAND2xp33_ASAP7_75t_L g3108 ( 
.A(n_2799),
.B(n_2561),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2894),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_SL g3110 ( 
.A(n_2944),
.B(n_2400),
.Y(n_3110)
);

NOR2x1p5_ASAP7_75t_L g3111 ( 
.A(n_2889),
.B(n_1158),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2886),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2898),
.B(n_2232),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2888),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2984),
.B(n_2400),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_3005),
.B(n_2430),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2872),
.A2(n_2227),
.B(n_2220),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2900),
.B(n_2731),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_3005),
.B(n_2430),
.Y(n_3119)
);

INVx4_ASAP7_75t_L g3120 ( 
.A(n_2857),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2926),
.A2(n_2365),
.B(n_2432),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2794),
.B(n_2432),
.Y(n_3122)
);

INVx1_ASAP7_75t_SL g3123 ( 
.A(n_2947),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2897),
.B(n_2435),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2893),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2943),
.B(n_2435),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2989),
.B(n_2437),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2965),
.B(n_2437),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2976),
.B(n_1192),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_2789),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2903),
.Y(n_3131)
);

A2O1A1Ixp33_ASAP7_75t_L g3132 ( 
.A1(n_3006),
.A2(n_2957),
.B(n_2982),
.C(n_2931),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_SL g3133 ( 
.A(n_2991),
.B(n_2439),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2871),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2895),
.Y(n_3135)
);

NAND2xp33_ASAP7_75t_L g3136 ( 
.A(n_2812),
.B(n_1185),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_3003),
.B(n_3015),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_3008),
.B(n_2439),
.Y(n_3138)
);

BUFx3_ASAP7_75t_L g3139 ( 
.A(n_2871),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2901),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2981),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_L g3142 ( 
.A(n_2812),
.B(n_1186),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_3017),
.B(n_1219),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_2968),
.B(n_2442),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2905),
.B(n_2442),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2923),
.B(n_2445),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2928),
.Y(n_3147)
);

CKINVDCx5p33_ASAP7_75t_R g3148 ( 
.A(n_2805),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2930),
.B(n_2445),
.Y(n_3149)
);

INVx2_ASAP7_75t_SL g3150 ( 
.A(n_2967),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2968),
.B(n_2452),
.Y(n_3151)
);

AND2x4_ASAP7_75t_L g3152 ( 
.A(n_2850),
.B(n_2718),
.Y(n_3152)
);

INVxp67_ASAP7_75t_L g3153 ( 
.A(n_2912),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2864),
.B(n_2452),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_3020),
.B(n_2874),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_3032),
.B(n_2460),
.Y(n_3156)
);

HB1xp67_ASAP7_75t_L g3157 ( 
.A(n_2927),
.Y(n_3157)
);

NAND2xp33_ASAP7_75t_SL g3158 ( 
.A(n_2945),
.B(n_1222),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2818),
.B(n_2460),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2835),
.B(n_1188),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2838),
.B(n_1191),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2908),
.B(n_2365),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2952),
.B(n_1249),
.Y(n_3163)
);

OR2x2_ASAP7_75t_L g3164 ( 
.A(n_2951),
.B(n_1160),
.Y(n_3164)
);

AND2x2_ASAP7_75t_SL g3165 ( 
.A(n_2813),
.B(n_1786),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2840),
.B(n_1193),
.Y(n_3166)
);

NOR2xp67_ASAP7_75t_L g3167 ( 
.A(n_2875),
.B(n_1003),
.Y(n_3167)
);

OR2x2_ASAP7_75t_L g3168 ( 
.A(n_2906),
.B(n_1160),
.Y(n_3168)
);

INVxp67_ASAP7_75t_L g3169 ( 
.A(n_2844),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_3010),
.B(n_1249),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2896),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_3028),
.A2(n_1273),
.B1(n_1274),
.B2(n_1261),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_2983),
.B(n_2995),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2840),
.A2(n_1273),
.B1(n_1274),
.B2(n_1261),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2992),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2824),
.B(n_1194),
.Y(n_3176)
);

BUFx4f_ASAP7_75t_L g3177 ( 
.A(n_2994),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2847),
.B(n_1195),
.Y(n_3178)
);

AOI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2845),
.A2(n_1317),
.B1(n_1329),
.B2(n_1299),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2929),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_SL g3181 ( 
.A(n_2994),
.B(n_1299),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3001),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2922),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_SL g3184 ( 
.A(n_2859),
.B(n_3031),
.Y(n_3184)
);

OR2x6_ASAP7_75t_L g3185 ( 
.A(n_2891),
.B(n_1787),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2847),
.B(n_1197),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2847),
.B(n_1198),
.Y(n_3187)
);

BUFx6f_ASAP7_75t_L g3188 ( 
.A(n_2795),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_2865),
.A2(n_1153),
.B(n_1156),
.C(n_1150),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2958),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3004),
.Y(n_3191)
);

NOR3xp33_ASAP7_75t_L g3192 ( 
.A(n_3025),
.B(n_1200),
.C(n_1199),
.Y(n_3192)
);

BUFx3_ASAP7_75t_L g3193 ( 
.A(n_2980),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2970),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2942),
.B(n_2979),
.Y(n_3195)
);

OAI22xp33_ASAP7_75t_L g3196 ( 
.A1(n_2924),
.A2(n_1329),
.B1(n_1335),
.B2(n_1317),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3011),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2972),
.Y(n_3198)
);

OR2x2_ASAP7_75t_L g3199 ( 
.A(n_3026),
.B(n_1164),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2915),
.B(n_1335),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2845),
.B(n_1201),
.Y(n_3201)
);

HB1xp67_ASAP7_75t_L g3202 ( 
.A(n_2936),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_SL g3203 ( 
.A(n_2962),
.B(n_1340),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2985),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_2921),
.A2(n_1345),
.B1(n_1357),
.B2(n_1340),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3024),
.Y(n_3206)
);

AOI22xp33_ASAP7_75t_L g3207 ( 
.A1(n_2934),
.A2(n_1357),
.B1(n_1371),
.B2(n_1345),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2845),
.B(n_1202),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2986),
.A2(n_1382),
.B1(n_1410),
.B2(n_1371),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2993),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2987),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_3016),
.B(n_1382),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_3021),
.B(n_1410),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_2919),
.B(n_1457),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_2910),
.B(n_1457),
.Y(n_3215)
);

INVxp67_ASAP7_75t_L g3216 ( 
.A(n_2913),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2996),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3030),
.B(n_1203),
.Y(n_3218)
);

NAND2x1_ASAP7_75t_L g3219 ( 
.A(n_2823),
.B(n_1545),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2998),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2978),
.B(n_1463),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3002),
.Y(n_3222)
);

AO22x1_ASAP7_75t_L g3223 ( 
.A1(n_2885),
.A2(n_1164),
.B1(n_1166),
.B2(n_1165),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_2962),
.B(n_1463),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2821),
.B(n_2917),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2842),
.B(n_1206),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3000),
.Y(n_3227)
);

NAND2xp33_ASAP7_75t_SL g3228 ( 
.A(n_2786),
.B(n_2866),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_2986),
.A2(n_1481),
.B1(n_1523),
.B2(n_1466),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2988),
.B(n_1466),
.Y(n_3230)
);

INVxp67_ASAP7_75t_L g3231 ( 
.A(n_2990),
.Y(n_3231)
);

O2A1O1Ixp33_ASAP7_75t_L g3232 ( 
.A1(n_2819),
.A2(n_1803),
.B(n_1840),
.C(n_1791),
.Y(n_3232)
);

AND2x6_ASAP7_75t_SL g3233 ( 
.A(n_2825),
.B(n_1162),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2986),
.B(n_1207),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2833),
.Y(n_3235)
);

OAI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_3132),
.A2(n_3019),
.B(n_3007),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_3225),
.A2(n_2861),
.B(n_2856),
.Y(n_3237)
);

AOI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_3039),
.A2(n_2935),
.B1(n_3018),
.B2(n_3014),
.Y(n_3238)
);

O2A1O1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_3137),
.A2(n_2890),
.B(n_2911),
.C(n_2867),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3067),
.B(n_2950),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3078),
.A2(n_2953),
.B(n_2946),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3079),
.A2(n_3027),
.B(n_2969),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_3049),
.B(n_2828),
.Y(n_3243)
);

BUFx6f_ASAP7_75t_L g3244 ( 
.A(n_3042),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3038),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3083),
.A2(n_3013),
.B(n_3022),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_3061),
.B(n_3012),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3070),
.B(n_2814),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3147),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3058),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3096),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3118),
.A2(n_2807),
.B(n_2878),
.Y(n_3252)
);

OAI21x1_ASAP7_75t_L g3253 ( 
.A1(n_3117),
.A2(n_3081),
.B(n_3121),
.Y(n_3253)
);

BUFx4f_ASAP7_75t_L g3254 ( 
.A(n_3072),
.Y(n_3254)
);

OAI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3071),
.A2(n_2939),
.B1(n_2854),
.B2(n_2938),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3097),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3131),
.B(n_2920),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3100),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3141),
.B(n_3029),
.Y(n_3259)
);

OAI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3098),
.A2(n_2949),
.B(n_2948),
.Y(n_3260)
);

NOR2xp33_ASAP7_75t_L g3261 ( 
.A(n_3143),
.B(n_2980),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3035),
.B(n_2854),
.Y(n_3262)
);

INVxp67_ASAP7_75t_L g3263 ( 
.A(n_3199),
.Y(n_3263)
);

CKINVDCx20_ASAP7_75t_R g3264 ( 
.A(n_3130),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3034),
.A2(n_2961),
.B(n_2956),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_3104),
.A2(n_3122),
.B(n_3156),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3175),
.B(n_3029),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3182),
.B(n_2963),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3191),
.B(n_2999),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3197),
.B(n_2932),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_3145),
.A2(n_2826),
.B(n_2823),
.Y(n_3271)
);

AO21x1_ASAP7_75t_L g3272 ( 
.A1(n_3041),
.A2(n_3082),
.B(n_3076),
.Y(n_3272)
);

NOR2xp67_ASAP7_75t_L g3273 ( 
.A(n_3090),
.B(n_2955),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3206),
.B(n_2941),
.Y(n_3274)
);

OR2x6_ASAP7_75t_L g3275 ( 
.A(n_3120),
.B(n_3134),
.Y(n_3275)
);

NOR2xp33_ASAP7_75t_L g3276 ( 
.A(n_3048),
.B(n_2997),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_3055),
.B(n_2966),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3045),
.Y(n_3278)
);

INVx2_ASAP7_75t_SL g3279 ( 
.A(n_3177),
.Y(n_3279)
);

A2O1A1Ixp33_ASAP7_75t_L g3280 ( 
.A1(n_3095),
.A2(n_2862),
.B(n_2887),
.C(n_2869),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3105),
.B(n_2902),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3109),
.B(n_2846),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3163),
.B(n_2826),
.Y(n_3283)
);

NOR3xp33_ASAP7_75t_L g3284 ( 
.A(n_3212),
.B(n_1210),
.C(n_1209),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3042),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3037),
.B(n_2892),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3218),
.B(n_2892),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3169),
.B(n_2907),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_3213),
.B(n_2829),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_3146),
.A2(n_2829),
.B(n_2907),
.Y(n_3290)
);

O2A1O1Ixp33_ASAP7_75t_L g3291 ( 
.A1(n_3153),
.A2(n_2937),
.B(n_1187),
.C(n_1189),
.Y(n_3291)
);

OAI321xp33_ASAP7_75t_L g3292 ( 
.A1(n_3196),
.A2(n_1168),
.A3(n_1204),
.B1(n_1208),
.B2(n_1205),
.C(n_1196),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_3149),
.A2(n_2914),
.B(n_1212),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3140),
.B(n_2940),
.Y(n_3294)
);

INVx2_ASAP7_75t_SL g3295 ( 
.A(n_3073),
.Y(n_3295)
);

AND2x4_ASAP7_75t_L g3296 ( 
.A(n_3139),
.B(n_2738),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3210),
.Y(n_3297)
);

OAI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_3166),
.A2(n_1221),
.B(n_1211),
.Y(n_3298)
);

OAI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3093),
.A2(n_1234),
.B(n_1227),
.Y(n_3299)
);

OAI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_3094),
.A2(n_3103),
.B(n_3099),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3053),
.Y(n_3301)
);

AOI21x1_ASAP7_75t_L g3302 ( 
.A1(n_3106),
.A2(n_1243),
.B(n_1237),
.Y(n_3302)
);

INVx4_ASAP7_75t_L g3303 ( 
.A(n_3193),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3154),
.A2(n_1258),
.B(n_1246),
.Y(n_3304)
);

OAI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3113),
.A2(n_1275),
.B(n_1263),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3124),
.A2(n_1289),
.B(n_1282),
.Y(n_3306)
);

HB1xp67_ASAP7_75t_L g3307 ( 
.A(n_3157),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3135),
.B(n_3176),
.Y(n_3308)
);

O2A1O1Ixp33_ASAP7_75t_L g3309 ( 
.A1(n_3189),
.A2(n_1304),
.B(n_1306),
.C(n_1301),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3054),
.B(n_2832),
.Y(n_3310)
);

AO21x1_ASAP7_75t_L g3311 ( 
.A1(n_3178),
.A2(n_1311),
.B(n_1308),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3217),
.A2(n_1327),
.B(n_1318),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3126),
.A2(n_3128),
.B(n_3159),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3056),
.B(n_1213),
.Y(n_3314)
);

AO21x1_ASAP7_75t_L g3315 ( 
.A1(n_3186),
.A2(n_1356),
.B(n_1355),
.Y(n_3315)
);

AND2x4_ASAP7_75t_L g3316 ( 
.A(n_3074),
.B(n_1359),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_3080),
.A2(n_1373),
.B(n_1365),
.Y(n_3317)
);

AO21x1_ASAP7_75t_L g3318 ( 
.A1(n_3187),
.A2(n_1378),
.B(n_1374),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3129),
.B(n_2954),
.Y(n_3319)
);

NAND2x1_ASAP7_75t_L g3320 ( 
.A(n_3050),
.B(n_1791),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3220),
.Y(n_3321)
);

INVx3_ASAP7_75t_L g3322 ( 
.A(n_3050),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3160),
.A2(n_1383),
.B(n_1381),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3161),
.A2(n_3142),
.B(n_3136),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3057),
.B(n_1214),
.Y(n_3325)
);

NAND2x1p5_ASAP7_75t_L g3326 ( 
.A(n_3069),
.B(n_2964),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3064),
.A2(n_1389),
.B(n_1385),
.Y(n_3327)
);

OAI21xp33_ASAP7_75t_L g3328 ( 
.A1(n_3207),
.A2(n_1523),
.B(n_1481),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3075),
.B(n_1215),
.Y(n_3329)
);

BUFx6f_ASAP7_75t_L g3330 ( 
.A(n_3188),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3086),
.A2(n_1396),
.B(n_1391),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3112),
.B(n_3114),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3125),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3222),
.B(n_1216),
.Y(n_3334)
);

A2O1A1Ixp33_ASAP7_75t_L g3335 ( 
.A1(n_3201),
.A2(n_1409),
.B(n_1411),
.C(n_1405),
.Y(n_3335)
);

INVxp67_ASAP7_75t_SL g3336 ( 
.A(n_3050),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3173),
.B(n_1217),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3047),
.B(n_1218),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3188),
.Y(n_3339)
);

AOI21xp33_ASAP7_75t_L g3340 ( 
.A1(n_3044),
.A2(n_1561),
.B(n_1525),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3194),
.B(n_1223),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_3216),
.A2(n_1416),
.B(n_1414),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3214),
.B(n_1525),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3063),
.B(n_1165),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3198),
.B(n_1226),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3226),
.A2(n_3062),
.B(n_3171),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3204),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3180),
.A2(n_1423),
.B(n_1419),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3051),
.A2(n_1577),
.B1(n_1583),
.B2(n_1561),
.Y(n_3349)
);

NOR2x1p5_ASAP7_75t_SL g3350 ( 
.A(n_3183),
.B(n_1803),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3211),
.B(n_1228),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3190),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3227),
.B(n_1230),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_3127),
.A2(n_1431),
.B(n_1424),
.Y(n_3354)
);

BUFx6f_ASAP7_75t_L g3355 ( 
.A(n_3066),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3133),
.A2(n_1438),
.B(n_1432),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_L g3357 ( 
.A(n_3091),
.B(n_1577),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3043),
.B(n_1231),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3231),
.A2(n_1444),
.B(n_1440),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3138),
.A2(n_1454),
.B(n_1448),
.Y(n_3360)
);

AOI21x1_ASAP7_75t_L g3361 ( 
.A1(n_3208),
.A2(n_1474),
.B(n_1455),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3101),
.B(n_1233),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3234),
.A2(n_1477),
.B(n_1475),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3232),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3066),
.Y(n_3365)
);

AOI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3059),
.A2(n_1591),
.B1(n_1614),
.B2(n_1583),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3168),
.B(n_1235),
.Y(n_3367)
);

O2A1O1Ixp5_ASAP7_75t_L g3368 ( 
.A1(n_3060),
.A2(n_1858),
.B(n_1840),
.C(n_1480),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3150),
.A2(n_1482),
.B(n_1479),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3200),
.B(n_1236),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3195),
.A2(n_1492),
.B(n_1484),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3215),
.B(n_1239),
.Y(n_3372)
);

BUFx3_ASAP7_75t_L g3373 ( 
.A(n_3072),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_3202),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3165),
.B(n_1591),
.Y(n_3375)
);

NAND3xp33_ASAP7_75t_L g3376 ( 
.A(n_3170),
.B(n_1242),
.C(n_1241),
.Y(n_3376)
);

NOR3xp33_ASAP7_75t_L g3377 ( 
.A(n_3033),
.B(n_1245),
.C(n_1244),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3221),
.B(n_1247),
.Y(n_3378)
);

AOI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_3219),
.A2(n_1494),
.B(n_1493),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3066),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_L g3381 ( 
.A(n_3089),
.B(n_1614),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_3123),
.B(n_1631),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3167),
.A2(n_1497),
.B(n_1496),
.Y(n_3383)
);

A2O1A1Ixp33_ASAP7_75t_L g3384 ( 
.A1(n_3230),
.A2(n_1505),
.B(n_1518),
.C(n_1498),
.Y(n_3384)
);

INVx4_ASAP7_75t_L g3385 ( 
.A(n_3148),
.Y(n_3385)
);

INVx4_ASAP7_75t_L g3386 ( 
.A(n_3077),
.Y(n_3386)
);

OAI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_3192),
.A2(n_1520),
.B(n_1519),
.Y(n_3387)
);

INVx3_ASAP7_75t_L g3388 ( 
.A(n_3303),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_3275),
.Y(n_3389)
);

O2A1O1Ixp33_ASAP7_75t_SL g3390 ( 
.A1(n_3240),
.A2(n_3052),
.B(n_3151),
.C(n_3144),
.Y(n_3390)
);

AOI22x1_ASAP7_75t_L g3391 ( 
.A1(n_3313),
.A2(n_3111),
.B1(n_3065),
.B2(n_3102),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3324),
.A2(n_3228),
.B(n_3108),
.Y(n_3392)
);

BUFx2_ASAP7_75t_L g3393 ( 
.A(n_3307),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3276),
.B(n_3036),
.Y(n_3394)
);

O2A1O1Ixp33_ASAP7_75t_L g3395 ( 
.A1(n_3298),
.A2(n_3181),
.B(n_3172),
.C(n_3203),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3277),
.B(n_3174),
.Y(n_3396)
);

OR2x6_ASAP7_75t_L g3397 ( 
.A(n_3279),
.B(n_3077),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3245),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3266),
.A2(n_3107),
.B(n_3155),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3250),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_R g3401 ( 
.A(n_3264),
.B(n_3235),
.Y(n_3401)
);

BUFx6f_ASAP7_75t_L g3402 ( 
.A(n_3244),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_L g3403 ( 
.A(n_3243),
.B(n_3068),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3300),
.A2(n_3115),
.B(n_3110),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3343),
.B(n_3040),
.Y(n_3405)
);

HB1xp67_ASAP7_75t_L g3406 ( 
.A(n_3374),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_R g3407 ( 
.A(n_3254),
.B(n_3184),
.Y(n_3407)
);

OAI22xp5_ASAP7_75t_SL g3408 ( 
.A1(n_3357),
.A2(n_3229),
.B1(n_3209),
.B2(n_3179),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3259),
.A2(n_3046),
.B1(n_3084),
.B2(n_3092),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3251),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3256),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3258),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_3247),
.B(n_3224),
.Y(n_3413)
);

AND2x4_ASAP7_75t_L g3414 ( 
.A(n_3373),
.B(n_3088),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3261),
.B(n_3205),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3267),
.B(n_3164),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_3269),
.A2(n_3085),
.B1(n_3119),
.B2(n_3116),
.Y(n_3417)
);

BUFx8_ASAP7_75t_L g3418 ( 
.A(n_3296),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3297),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3283),
.B(n_3223),
.Y(n_3420)
);

CKINVDCx10_ASAP7_75t_R g3421 ( 
.A(n_3275),
.Y(n_3421)
);

INVxp67_ASAP7_75t_L g3422 ( 
.A(n_3381),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3375),
.B(n_3185),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_3244),
.Y(n_3424)
);

INVx5_ASAP7_75t_L g3425 ( 
.A(n_3355),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3239),
.A2(n_3158),
.B(n_3087),
.C(n_3162),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_3285),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3321),
.Y(n_3428)
);

OAI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_3257),
.A2(n_3238),
.B1(n_3308),
.B2(n_3268),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_3340),
.B(n_3152),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3382),
.B(n_3185),
.Y(n_3431)
);

OAI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3349),
.A2(n_1640),
.B1(n_1673),
.B2(n_1631),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_3385),
.Y(n_3433)
);

INVx1_ASAP7_75t_SL g3434 ( 
.A(n_3295),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3249),
.Y(n_3435)
);

INVx2_ASAP7_75t_SL g3436 ( 
.A(n_3285),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3278),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_3330),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_3330),
.Y(n_3439)
);

OR2x2_ASAP7_75t_L g3440 ( 
.A(n_3344),
.B(n_1166),
.Y(n_3440)
);

AOI21x1_ASAP7_75t_L g3441 ( 
.A1(n_3237),
.A2(n_1524),
.B(n_1521),
.Y(n_3441)
);

INVx4_ASAP7_75t_L g3442 ( 
.A(n_3339),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_3286),
.A2(n_1640),
.B1(n_1673),
.B2(n_1668),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3328),
.B(n_3233),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3289),
.B(n_2741),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_3263),
.B(n_1167),
.Y(n_3446)
);

HB1xp67_ASAP7_75t_L g3447 ( 
.A(n_3339),
.Y(n_3447)
);

OAI21xp33_ASAP7_75t_SL g3448 ( 
.A1(n_3312),
.A2(n_1533),
.B(n_1530),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3337),
.B(n_1536),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3316),
.B(n_1248),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_SL g3451 ( 
.A1(n_3319),
.A2(n_1668),
.B1(n_1706),
.B2(n_1674),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3241),
.A2(n_3346),
.B(n_3236),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3287),
.B(n_3272),
.Y(n_3453)
);

O2A1O1Ixp33_ASAP7_75t_L g3454 ( 
.A1(n_3370),
.A2(n_1552),
.B(n_1553),
.C(n_1542),
.Y(n_3454)
);

OR2x6_ASAP7_75t_L g3455 ( 
.A(n_3386),
.B(n_1858),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3316),
.B(n_1250),
.Y(n_3456)
);

NAND2xp33_ASAP7_75t_L g3457 ( 
.A(n_3284),
.B(n_3355),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3372),
.B(n_1674),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3366),
.A2(n_1928),
.B1(n_1924),
.B2(n_1723),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3332),
.Y(n_3460)
);

NOR2x1_ASAP7_75t_L g3461 ( 
.A(n_3242),
.B(n_1924),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3301),
.Y(n_3462)
);

INVx3_ASAP7_75t_L g3463 ( 
.A(n_3322),
.Y(n_3463)
);

OAI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3270),
.A2(n_1706),
.B1(n_1737),
.B2(n_1723),
.Y(n_3464)
);

O2A1O1Ixp33_ASAP7_75t_L g3465 ( 
.A1(n_3378),
.A2(n_1558),
.B(n_1563),
.C(n_1554),
.Y(n_3465)
);

NOR2xp67_ASAP7_75t_L g3466 ( 
.A(n_3252),
.B(n_1005),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3274),
.A2(n_1737),
.B1(n_1806),
.B2(n_1794),
.Y(n_3467)
);

AOI21x1_ASAP7_75t_L g3468 ( 
.A1(n_3253),
.A2(n_1571),
.B(n_1570),
.Y(n_3468)
);

OAI22x1_ASAP7_75t_L g3469 ( 
.A1(n_3262),
.A2(n_3376),
.B1(n_3310),
.B2(n_3338),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3384),
.A2(n_1582),
.B(n_1589),
.C(n_1575),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3367),
.B(n_1794),
.Y(n_3471)
);

BUFx2_ASAP7_75t_L g3472 ( 
.A(n_3380),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3333),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3246),
.A2(n_1599),
.B(n_1595),
.Y(n_3474)
);

O2A1O1Ixp33_ASAP7_75t_L g3475 ( 
.A1(n_3292),
.A2(n_1621),
.B(n_1622),
.C(n_1602),
.Y(n_3475)
);

O2A1O1Ixp5_ASAP7_75t_L g3476 ( 
.A1(n_3311),
.A2(n_1629),
.B(n_1632),
.C(n_1626),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3288),
.B(n_1806),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3342),
.B(n_1642),
.Y(n_3478)
);

NOR2x1_ASAP7_75t_L g3479 ( 
.A(n_3248),
.B(n_1826),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3377),
.A2(n_1831),
.B1(n_1848),
.B2(n_1826),
.Y(n_3480)
);

BUFx2_ASAP7_75t_L g3481 ( 
.A(n_3365),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_SL g3482 ( 
.A(n_3359),
.B(n_1831),
.Y(n_3482)
);

AOI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3362),
.A2(n_3358),
.B1(n_3255),
.B2(n_3334),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3273),
.B(n_1848),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_3260),
.A2(n_1644),
.B(n_1643),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3282),
.A2(n_3347),
.B1(n_3281),
.B2(n_3352),
.Y(n_3486)
);

AOI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_3315),
.A2(n_1928),
.B1(n_1918),
.B2(n_1852),
.Y(n_3487)
);

O2A1O1Ixp33_ASAP7_75t_SL g3488 ( 
.A1(n_3335),
.A2(n_1676),
.B(n_1686),
.C(n_1650),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3299),
.B(n_1850),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3280),
.A2(n_1850),
.B1(n_1866),
.B2(n_1852),
.Y(n_3490)
);

OR2x2_ASAP7_75t_L g3491 ( 
.A(n_3341),
.B(n_1167),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3305),
.B(n_1691),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3364),
.A2(n_1693),
.B(n_1692),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3302),
.Y(n_3494)
);

HB1xp67_ASAP7_75t_L g3495 ( 
.A(n_3336),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_3294),
.Y(n_3496)
);

BUFx3_ASAP7_75t_L g3497 ( 
.A(n_3326),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3265),
.A2(n_1696),
.B(n_1695),
.Y(n_3498)
);

A2O1A1Ixp33_ASAP7_75t_L g3499 ( 
.A1(n_3387),
.A2(n_1703),
.B(n_1704),
.C(n_1698),
.Y(n_3499)
);

A2O1A1Ixp33_ASAP7_75t_L g3500 ( 
.A1(n_3368),
.A2(n_1710),
.B(n_1711),
.C(n_1705),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3320),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3345),
.B(n_1918),
.Y(n_3502)
);

HB1xp67_ASAP7_75t_L g3503 ( 
.A(n_3314),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3350),
.Y(n_3504)
);

NOR2xp33_ASAP7_75t_L g3505 ( 
.A(n_3351),
.B(n_1866),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3325),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3353),
.B(n_1716),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3329),
.A2(n_3290),
.B1(n_3271),
.B2(n_3293),
.Y(n_3508)
);

NOR2xp33_ASAP7_75t_L g3509 ( 
.A(n_3369),
.B(n_1868),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_3317),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_3383),
.A2(n_3348),
.B(n_3363),
.C(n_3323),
.Y(n_3511)
);

INVx3_ASAP7_75t_L g3512 ( 
.A(n_3361),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3304),
.Y(n_3513)
);

OR2x6_ASAP7_75t_L g3514 ( 
.A(n_3379),
.B(n_1718),
.Y(n_3514)
);

O2A1O1Ixp33_ASAP7_75t_L g3515 ( 
.A1(n_3306),
.A2(n_1728),
.B(n_1731),
.C(n_1720),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3327),
.A2(n_1745),
.B(n_1738),
.Y(n_3516)
);

NOR3xp33_ASAP7_75t_L g3517 ( 
.A(n_3291),
.B(n_1815),
.C(n_1764),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3318),
.B(n_1868),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3331),
.A2(n_1749),
.B(n_1747),
.Y(n_3519)
);

AOI221xp5_ASAP7_75t_L g3520 ( 
.A1(n_3309),
.A2(n_3356),
.B1(n_3360),
.B2(n_3354),
.C(n_3371),
.Y(n_3520)
);

CKINVDCx10_ASAP7_75t_R g3521 ( 
.A(n_3275),
.Y(n_3521)
);

NAND3xp33_ASAP7_75t_SL g3522 ( 
.A(n_3284),
.B(n_1877),
.C(n_1929),
.Y(n_3522)
);

OAI22xp5_ASAP7_75t_SL g3523 ( 
.A1(n_3357),
.A2(n_1877),
.B1(n_1929),
.B2(n_1927),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3276),
.A2(n_1930),
.B1(n_1931),
.B2(n_1927),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3276),
.B(n_1750),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3324),
.A2(n_1755),
.B(n_1752),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3245),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_3388),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3452),
.A2(n_1759),
.B(n_1758),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3394),
.B(n_1253),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3400),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3411),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_L g3533 ( 
.A(n_3403),
.B(n_1255),
.Y(n_3533)
);

O2A1O1Ixp5_ASAP7_75t_L g3534 ( 
.A1(n_3489),
.A2(n_1775),
.B(n_1779),
.C(n_1767),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3413),
.B(n_1930),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3419),
.Y(n_3536)
);

NAND3xp33_ASAP7_75t_SL g3537 ( 
.A(n_3395),
.B(n_1934),
.C(n_1933),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3458),
.B(n_1933),
.Y(n_3538)
);

AND2x4_ASAP7_75t_L g3539 ( 
.A(n_3497),
.B(n_1784),
.Y(n_3539)
);

O2A1O1Ixp5_ASAP7_75t_SL g3540 ( 
.A1(n_3512),
.A2(n_1914),
.B(n_1915),
.C(n_1911),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_3402),
.Y(n_3541)
);

INVx3_ASAP7_75t_L g3542 ( 
.A(n_3442),
.Y(n_3542)
);

BUFx12f_ASAP7_75t_L g3543 ( 
.A(n_3418),
.Y(n_3543)
);

AO21x2_ASAP7_75t_L g3544 ( 
.A1(n_3468),
.A2(n_1793),
.B(n_1788),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3415),
.B(n_1935),
.Y(n_3545)
);

BUFx6f_ASAP7_75t_L g3546 ( 
.A(n_3402),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3405),
.B(n_3477),
.Y(n_3547)
);

AOI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3441),
.A2(n_1799),
.B(n_1798),
.Y(n_3548)
);

OA21x2_ASAP7_75t_L g3549 ( 
.A1(n_3453),
.A2(n_1923),
.B(n_1920),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3392),
.A2(n_1805),
.B(n_1800),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3399),
.A2(n_1809),
.B(n_1808),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3398),
.Y(n_3552)
);

AOI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3469),
.A2(n_1817),
.B(n_1810),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3410),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3508),
.A2(n_1827),
.B(n_1825),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3404),
.A2(n_1832),
.B(n_1830),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3412),
.Y(n_3557)
);

A2O1A1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3525),
.A2(n_1837),
.B(n_1842),
.C(n_1836),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3396),
.B(n_1935),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3428),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3527),
.Y(n_3561)
);

INVx1_ASAP7_75t_SL g3562 ( 
.A(n_3393),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3505),
.B(n_1256),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3435),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3511),
.A2(n_1856),
.B(n_1843),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3429),
.A2(n_1869),
.B(n_1864),
.Y(n_3566)
);

INVxp67_ASAP7_75t_L g3567 ( 
.A(n_3406),
.Y(n_3567)
);

OAI21x1_ASAP7_75t_L g3568 ( 
.A1(n_3526),
.A2(n_1872),
.B(n_1871),
.Y(n_3568)
);

NOR4xp25_ASAP7_75t_L g3569 ( 
.A(n_3482),
.B(n_1875),
.C(n_1876),
.D(n_1873),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_SL g3570 ( 
.A(n_3433),
.B(n_1905),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3466),
.A2(n_1882),
.B(n_1879),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3494),
.A2(n_1893),
.B(n_1888),
.Y(n_3572)
);

INVx2_ASAP7_75t_SL g3573 ( 
.A(n_3421),
.Y(n_3573)
);

AOI31xp67_ASAP7_75t_L g3574 ( 
.A1(n_3483),
.A2(n_1008),
.A3(n_1010),
.B(n_1007),
.Y(n_3574)
);

BUFx2_ASAP7_75t_L g3575 ( 
.A(n_3438),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3437),
.Y(n_3576)
);

A2O1A1Ixp33_ASAP7_75t_L g3577 ( 
.A1(n_3509),
.A2(n_1916),
.B(n_1932),
.C(n_1909),
.Y(n_3577)
);

BUFx2_ASAP7_75t_L g3578 ( 
.A(n_3447),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3390),
.A2(n_1016),
.B(n_1013),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_3513),
.A2(n_1020),
.B(n_1018),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3462),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3417),
.A2(n_1027),
.B(n_1026),
.Y(n_3582)
);

AO32x2_ASAP7_75t_L g3583 ( 
.A1(n_3408),
.A2(n_3),
.A3(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_3583)
);

INVx3_ASAP7_75t_L g3584 ( 
.A(n_3439),
.Y(n_3584)
);

AND2x4_ASAP7_75t_L g3585 ( 
.A(n_3414),
.B(n_1029),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3416),
.B(n_1262),
.Y(n_3586)
);

BUFx3_ASAP7_75t_L g3587 ( 
.A(n_3424),
.Y(n_3587)
);

AOI21x1_ASAP7_75t_L g3588 ( 
.A1(n_3485),
.A2(n_1034),
.B(n_1033),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3471),
.B(n_3506),
.Y(n_3589)
);

OAI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3478),
.A2(n_1913),
.B(n_1912),
.Y(n_3590)
);

AO31x2_ASAP7_75t_L g3591 ( 
.A1(n_3504),
.A2(n_3474),
.A3(n_3498),
.B(n_3500),
.Y(n_3591)
);

OR2x6_ASAP7_75t_L g3592 ( 
.A(n_3397),
.B(n_1035),
.Y(n_3592)
);

AO22x2_ASAP7_75t_L g3593 ( 
.A1(n_3409),
.A2(n_5),
.B1(n_1),
.B2(n_3),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3473),
.Y(n_3594)
);

NAND2x1p5_ASAP7_75t_L g3595 ( 
.A(n_3425),
.B(n_1037),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3460),
.B(n_1264),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3486),
.Y(n_3597)
);

INVx1_ASAP7_75t_SL g3598 ( 
.A(n_3434),
.Y(n_3598)
);

INVx2_ASAP7_75t_SL g3599 ( 
.A(n_3521),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3493),
.A2(n_1042),
.B(n_1041),
.Y(n_3600)
);

AOI22xp5_ASAP7_75t_L g3601 ( 
.A1(n_3430),
.A2(n_1267),
.B1(n_1268),
.B2(n_1266),
.Y(n_3601)
);

AND2x4_ASAP7_75t_L g3602 ( 
.A(n_3397),
.B(n_1044),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3510),
.B(n_1904),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3492),
.A2(n_1048),
.B(n_1047),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3422),
.B(n_1269),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_3391),
.A2(n_1053),
.B(n_1049),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_3520),
.A2(n_1058),
.B(n_1054),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3426),
.A2(n_1063),
.B(n_1061),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3449),
.A2(n_3503),
.B(n_3507),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3423),
.B(n_1270),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3420),
.A2(n_1277),
.B1(n_1278),
.B2(n_1272),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3461),
.A2(n_1065),
.B(n_1064),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3432),
.B(n_1903),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3518),
.B(n_1280),
.Y(n_3614)
);

OAI22x1_ASAP7_75t_L g3615 ( 
.A1(n_3459),
.A2(n_3480),
.B1(n_3487),
.B2(n_3444),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_3502),
.B(n_1283),
.Y(n_3616)
);

AOI21x1_ASAP7_75t_L g3617 ( 
.A1(n_3501),
.A2(n_1069),
.B(n_1067),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3464),
.B(n_1284),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3467),
.B(n_1286),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3481),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3457),
.A2(n_3465),
.B(n_3454),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3472),
.Y(n_3622)
);

CKINVDCx16_ASAP7_75t_R g3623 ( 
.A(n_3401),
.Y(n_3623)
);

NAND3x1_ASAP7_75t_L g3624 ( 
.A(n_3479),
.B(n_6),
.C(n_7),
.Y(n_3624)
);

NOR2x1_ASAP7_75t_SL g3625 ( 
.A(n_3425),
.B(n_1071),
.Y(n_3625)
);

AND2x6_ASAP7_75t_L g3626 ( 
.A(n_3389),
.B(n_1072),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3443),
.B(n_1288),
.Y(n_3627)
);

OR2x6_ASAP7_75t_L g3628 ( 
.A(n_3424),
.B(n_1075),
.Y(n_3628)
);

OAI21x1_ASAP7_75t_SL g3629 ( 
.A1(n_3470),
.A2(n_6),
.B(n_8),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3450),
.B(n_1291),
.Y(n_3630)
);

O2A1O1Ixp33_ASAP7_75t_SL g3631 ( 
.A1(n_3499),
.A2(n_11),
.B(n_8),
.C(n_9),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3456),
.B(n_1293),
.Y(n_3632)
);

NAND3xp33_ASAP7_75t_SL g3633 ( 
.A(n_3475),
.B(n_3517),
.C(n_3407),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3495),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3488),
.A2(n_3476),
.B(n_3448),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3484),
.A2(n_1296),
.B(n_1295),
.Y(n_3636)
);

AOI221xp5_ASAP7_75t_L g3637 ( 
.A1(n_3524),
.A2(n_1303),
.B1(n_1305),
.B2(n_1300),
.C(n_1297),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3496),
.B(n_1307),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3620),
.Y(n_3639)
);

OAI21x1_ASAP7_75t_L g3640 ( 
.A1(n_3606),
.A2(n_3519),
.B(n_3516),
.Y(n_3640)
);

BUFx6f_ASAP7_75t_L g3641 ( 
.A(n_3541),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3634),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3579),
.A2(n_3515),
.B(n_3463),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_SL g3644 ( 
.A1(n_3628),
.A2(n_3633),
.B(n_3592),
.Y(n_3644)
);

AO31x2_ASAP7_75t_L g3645 ( 
.A1(n_3565),
.A2(n_3445),
.A3(n_3431),
.B(n_3490),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3607),
.A2(n_3582),
.B(n_3608),
.Y(n_3646)
);

INVx4_ASAP7_75t_L g3647 ( 
.A(n_3541),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3572),
.A2(n_3491),
.B(n_3522),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3609),
.B(n_3451),
.Y(n_3649)
);

INVx3_ASAP7_75t_L g3650 ( 
.A(n_3584),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_SL g3651 ( 
.A1(n_3533),
.A2(n_3523),
.B1(n_3514),
.B2(n_3440),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3589),
.B(n_3446),
.Y(n_3652)
);

NOR2xp67_ASAP7_75t_L g3653 ( 
.A(n_3528),
.B(n_3425),
.Y(n_3653)
);

OAI22xp5_ASAP7_75t_L g3654 ( 
.A1(n_3545),
.A2(n_3455),
.B1(n_3514),
.B2(n_3436),
.Y(n_3654)
);

NAND2x1p5_ASAP7_75t_L g3655 ( 
.A(n_3562),
.B(n_3578),
.Y(n_3655)
);

AND2x2_ASAP7_75t_SL g3656 ( 
.A(n_3623),
.B(n_3427),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3536),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3552),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3576),
.Y(n_3659)
);

INVx3_ASAP7_75t_L g3660 ( 
.A(n_3542),
.Y(n_3660)
);

OAI21xp33_ASAP7_75t_L g3661 ( 
.A1(n_3530),
.A2(n_3455),
.B(n_1310),
.Y(n_3661)
);

INVxp67_ASAP7_75t_L g3662 ( 
.A(n_3575),
.Y(n_3662)
);

NOR4xp25_ASAP7_75t_L g3663 ( 
.A(n_3624),
.B(n_12),
.C(n_9),
.D(n_11),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3554),
.Y(n_3664)
);

O2A1O1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_3621),
.A2(n_1894),
.B(n_1895),
.C(n_1892),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3557),
.Y(n_3666)
);

OAI21x1_ASAP7_75t_SL g3667 ( 
.A1(n_3553),
.A2(n_12),
.B(n_13),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3547),
.B(n_3427),
.Y(n_3668)
);

OAI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3614),
.A2(n_1312),
.B1(n_1314),
.B2(n_1309),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3615),
.A2(n_1316),
.B1(n_1319),
.B2(n_1315),
.Y(n_3670)
);

BUFx8_ASAP7_75t_L g3671 ( 
.A(n_3543),
.Y(n_3671)
);

OAI22x1_ASAP7_75t_L g3672 ( 
.A1(n_3597),
.A2(n_3560),
.B1(n_3561),
.B2(n_3603),
.Y(n_3672)
);

OA21x2_ASAP7_75t_L g3673 ( 
.A1(n_3555),
.A2(n_1324),
.B(n_1320),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3581),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3622),
.B(n_13),
.Y(n_3675)
);

OAI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3588),
.A2(n_3548),
.B(n_3529),
.Y(n_3676)
);

BUFx2_ASAP7_75t_L g3677 ( 
.A(n_3549),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_3638),
.B(n_1325),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3587),
.Y(n_3679)
);

NAND2xp33_ASAP7_75t_SL g3680 ( 
.A(n_3535),
.B(n_3602),
.Y(n_3680)
);

OAI21x1_ASAP7_75t_L g3681 ( 
.A1(n_3600),
.A2(n_15),
.B(n_16),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3531),
.B(n_16),
.Y(n_3682)
);

BUFx3_ASAP7_75t_L g3683 ( 
.A(n_3546),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3537),
.A2(n_1331),
.B1(n_1333),
.B2(n_1326),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3569),
.B(n_1336),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_SL g3686 ( 
.A1(n_3629),
.A2(n_17),
.B(n_18),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3532),
.B(n_17),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3564),
.Y(n_3688)
);

INVxp67_ASAP7_75t_SL g3689 ( 
.A(n_3567),
.Y(n_3689)
);

BUFx2_ASAP7_75t_L g3690 ( 
.A(n_3593),
.Y(n_3690)
);

OAI211xp5_ASAP7_75t_L g3691 ( 
.A1(n_3613),
.A2(n_1902),
.B(n_1906),
.C(n_1900),
.Y(n_3691)
);

AOI22xp33_ASAP7_75t_L g3692 ( 
.A1(n_3593),
.A2(n_1341),
.B1(n_1342),
.B2(n_1337),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3540),
.A2(n_18),
.B(n_19),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3594),
.Y(n_3694)
);

OAI22x1_ASAP7_75t_L g3695 ( 
.A1(n_3601),
.A2(n_1344),
.B1(n_1346),
.B2(n_1343),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3583),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3568),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3610),
.B(n_21),
.Y(n_3698)
);

OAI21x1_ASAP7_75t_L g3699 ( 
.A1(n_3551),
.A2(n_22),
.B(n_23),
.Y(n_3699)
);

AOI22xp33_ASAP7_75t_L g3700 ( 
.A1(n_3616),
.A2(n_1348),
.B1(n_1351),
.B2(n_1347),
.Y(n_3700)
);

BUFx2_ASAP7_75t_L g3701 ( 
.A(n_3546),
.Y(n_3701)
);

O2A1O1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3577),
.A2(n_1891),
.B(n_1896),
.C(n_1890),
.Y(n_3702)
);

OAI22xp5_ASAP7_75t_L g3703 ( 
.A1(n_3538),
.A2(n_1360),
.B1(n_1361),
.B2(n_1353),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_SL g3704 ( 
.A1(n_3566),
.A2(n_22),
.B(n_23),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3617),
.A2(n_24),
.B(n_25),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3583),
.Y(n_3706)
);

OAI21x1_ASAP7_75t_L g3707 ( 
.A1(n_3550),
.A2(n_24),
.B(n_26),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3598),
.Y(n_3708)
);

OAI21x1_ASAP7_75t_L g3709 ( 
.A1(n_3635),
.A2(n_26),
.B(n_27),
.Y(n_3709)
);

OR2x6_ASAP7_75t_L g3710 ( 
.A(n_3628),
.B(n_27),
.Y(n_3710)
);

BUFx3_ASAP7_75t_L g3711 ( 
.A(n_3573),
.Y(n_3711)
);

OAI21x1_ASAP7_75t_L g3712 ( 
.A1(n_3556),
.A2(n_28),
.B(n_29),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3574),
.Y(n_3713)
);

OAI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3563),
.A2(n_1367),
.B(n_1362),
.Y(n_3714)
);

CKINVDCx20_ASAP7_75t_R g3715 ( 
.A(n_3671),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3668),
.B(n_3632),
.Y(n_3716)
);

INVx1_ASAP7_75t_SL g3717 ( 
.A(n_3708),
.Y(n_3717)
);

OA21x2_ASAP7_75t_L g3718 ( 
.A1(n_3705),
.A2(n_3571),
.B(n_3612),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_3711),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3688),
.Y(n_3720)
);

OAI21x1_ASAP7_75t_SL g3721 ( 
.A1(n_3686),
.A2(n_3667),
.B(n_3704),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3641),
.Y(n_3722)
);

OAI21x1_ASAP7_75t_L g3723 ( 
.A1(n_3676),
.A2(n_3580),
.B(n_3604),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3694),
.Y(n_3724)
);

OAI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3646),
.A2(n_3595),
.B(n_3534),
.Y(n_3725)
);

OAI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3665),
.A2(n_3590),
.B(n_3627),
.Y(n_3726)
);

CKINVDCx20_ASAP7_75t_R g3727 ( 
.A(n_3680),
.Y(n_3727)
);

AO21x2_ASAP7_75t_L g3728 ( 
.A1(n_3713),
.A2(n_3544),
.B(n_3631),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3644),
.A2(n_3625),
.B(n_3592),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3642),
.B(n_3586),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3658),
.Y(n_3731)
);

O2A1O1Ixp33_ASAP7_75t_L g3732 ( 
.A1(n_3649),
.A2(n_3619),
.B(n_3618),
.C(n_3558),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3664),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3666),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_SL g3735 ( 
.A1(n_3710),
.A2(n_3559),
.B(n_3596),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3657),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3652),
.B(n_3570),
.Y(n_3737)
);

OA21x2_ASAP7_75t_L g3738 ( 
.A1(n_3709),
.A2(n_3636),
.B(n_3630),
.Y(n_3738)
);

BUFx8_ASAP7_75t_SL g3739 ( 
.A(n_3701),
.Y(n_3739)
);

INVxp67_ASAP7_75t_L g3740 ( 
.A(n_3639),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3689),
.B(n_3659),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3690),
.Y(n_3742)
);

BUFx12f_ASAP7_75t_L g3743 ( 
.A(n_3641),
.Y(n_3743)
);

INVxp67_ASAP7_75t_SL g3744 ( 
.A(n_3677),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3640),
.A2(n_3591),
.B(n_3611),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3674),
.B(n_3605),
.Y(n_3746)
);

OA21x2_ASAP7_75t_L g3747 ( 
.A1(n_3681),
.A2(n_3539),
.B(n_3637),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3690),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3672),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3662),
.B(n_3626),
.Y(n_3750)
);

NAND2x1p5_ASAP7_75t_L g3751 ( 
.A(n_3656),
.B(n_3585),
.Y(n_3751)
);

OAI21x1_ASAP7_75t_L g3752 ( 
.A1(n_3643),
.A2(n_3591),
.B(n_3626),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3697),
.A2(n_3626),
.B(n_28),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3655),
.B(n_3599),
.Y(n_3754)
);

OR2x6_ASAP7_75t_L g3755 ( 
.A(n_3710),
.B(n_29),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3673),
.A2(n_1369),
.B(n_1368),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3693),
.A2(n_30),
.B(n_33),
.Y(n_3757)
);

AOI21x1_ASAP7_75t_L g3758 ( 
.A1(n_3677),
.A2(n_1375),
.B(n_1372),
.Y(n_3758)
);

OAI21x1_ASAP7_75t_L g3759 ( 
.A1(n_3699),
.A2(n_30),
.B(n_33),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3663),
.B(n_1377),
.Y(n_3760)
);

OR2x6_ASAP7_75t_L g3761 ( 
.A(n_3648),
.B(n_34),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3682),
.B(n_1379),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3687),
.B(n_1380),
.Y(n_3763)
);

OA21x2_ASAP7_75t_L g3764 ( 
.A1(n_3712),
.A2(n_1386),
.B(n_1384),
.Y(n_3764)
);

BUFx3_ASAP7_75t_L g3765 ( 
.A(n_3683),
.Y(n_3765)
);

OAI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3670),
.A2(n_1392),
.B(n_1390),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3696),
.Y(n_3767)
);

BUFx2_ASAP7_75t_L g3768 ( 
.A(n_3679),
.Y(n_3768)
);

AND2x4_ASAP7_75t_L g3769 ( 
.A(n_3650),
.B(n_35),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3706),
.B(n_1395),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_3647),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3740),
.B(n_3698),
.Y(n_3772)
);

INVx3_ASAP7_75t_L g3773 ( 
.A(n_3733),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3731),
.Y(n_3774)
);

AO21x2_ASAP7_75t_L g3775 ( 
.A1(n_3758),
.A2(n_3685),
.B(n_3714),
.Y(n_3775)
);

AO21x2_ASAP7_75t_L g3776 ( 
.A1(n_3745),
.A2(n_3707),
.B(n_3653),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3734),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3720),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3724),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_SL g3780 ( 
.A(n_3729),
.B(n_3651),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3742),
.Y(n_3781)
);

OAI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3752),
.A2(n_3673),
.B(n_3654),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3741),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3748),
.Y(n_3784)
);

AO21x2_ASAP7_75t_L g3785 ( 
.A1(n_3749),
.A2(n_3661),
.B(n_3669),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3767),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3723),
.A2(n_3702),
.B(n_3692),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3736),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3768),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3744),
.Y(n_3790)
);

OR2x2_ASAP7_75t_L g3791 ( 
.A(n_3730),
.B(n_3717),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3746),
.Y(n_3792)
);

INVxp67_ASAP7_75t_L g3793 ( 
.A(n_3737),
.Y(n_3793)
);

CKINVDCx5p33_ASAP7_75t_R g3794 ( 
.A(n_3715),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3725),
.A2(n_3660),
.B(n_3675),
.Y(n_3795)
);

AND2x4_ASAP7_75t_L g3796 ( 
.A(n_3750),
.B(n_3645),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3770),
.Y(n_3797)
);

BUFx2_ASAP7_75t_L g3798 ( 
.A(n_3739),
.Y(n_3798)
);

INVxp67_ASAP7_75t_SL g3799 ( 
.A(n_3759),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3765),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3754),
.B(n_3645),
.Y(n_3801)
);

BUFx2_ASAP7_75t_SL g3802 ( 
.A(n_3727),
.Y(n_3802)
);

OR2x6_ASAP7_75t_L g3803 ( 
.A(n_3735),
.B(n_3695),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3761),
.Y(n_3804)
);

AO21x2_ASAP7_75t_L g3805 ( 
.A1(n_3756),
.A2(n_3703),
.B(n_3691),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3716),
.B(n_3678),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3761),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3728),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3722),
.Y(n_3809)
);

OAI21x1_ASAP7_75t_L g3810 ( 
.A1(n_3753),
.A2(n_3684),
.B(n_3700),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3757),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3760),
.B(n_1397),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3721),
.Y(n_3813)
);

HB1xp67_ASAP7_75t_L g3814 ( 
.A(n_3764),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3764),
.Y(n_3815)
);

OR2x2_ASAP7_75t_L g3816 ( 
.A(n_3762),
.B(n_36),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3738),
.Y(n_3817)
);

AOI22xp33_ASAP7_75t_L g3818 ( 
.A1(n_3726),
.A2(n_1399),
.B1(n_1400),
.B2(n_1398),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3738),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3718),
.Y(n_3820)
);

INVx3_ASAP7_75t_L g3821 ( 
.A(n_3743),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3769),
.Y(n_3822)
);

BUFx2_ASAP7_75t_L g3823 ( 
.A(n_3771),
.Y(n_3823)
);

INVxp67_ASAP7_75t_L g3824 ( 
.A(n_3722),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3719),
.Y(n_3825)
);

INVx5_ASAP7_75t_SL g3826 ( 
.A(n_3755),
.Y(n_3826)
);

HB1xp67_ASAP7_75t_L g3827 ( 
.A(n_3747),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3751),
.B(n_37),
.Y(n_3828)
);

CKINVDCx20_ASAP7_75t_R g3829 ( 
.A(n_3763),
.Y(n_3829)
);

OAI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3732),
.A2(n_3766),
.B(n_3755),
.Y(n_3830)
);

NAND3xp33_ASAP7_75t_L g3831 ( 
.A(n_3818),
.B(n_1402),
.C(n_1401),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3786),
.Y(n_3832)
);

AOI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3780),
.A2(n_1413),
.B1(n_1417),
.B2(n_1415),
.Y(n_3833)
);

BUFx3_ASAP7_75t_L g3834 ( 
.A(n_3798),
.Y(n_3834)
);

AOI22xp33_ASAP7_75t_L g3835 ( 
.A1(n_3803),
.A2(n_1874),
.B1(n_1878),
.B2(n_1870),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3777),
.Y(n_3836)
);

AOI22xp33_ASAP7_75t_L g3837 ( 
.A1(n_3803),
.A2(n_1884),
.B1(n_1885),
.B2(n_1881),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3789),
.B(n_3801),
.Y(n_3838)
);

AO21x2_ASAP7_75t_L g3839 ( 
.A1(n_3817),
.A2(n_48),
.B(n_38),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3796),
.A2(n_3805),
.B1(n_3807),
.B2(n_3804),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3783),
.B(n_1412),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3773),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3772),
.B(n_38),
.Y(n_3843)
);

OAI21x1_ASAP7_75t_L g3844 ( 
.A1(n_3782),
.A2(n_3795),
.B(n_3808),
.Y(n_3844)
);

INVxp33_ASAP7_75t_L g3845 ( 
.A(n_3823),
.Y(n_3845)
);

OAI222xp33_ASAP7_75t_L g3846 ( 
.A1(n_3793),
.A2(n_1425),
.B1(n_1421),
.B2(n_1429),
.C1(n_1422),
.C2(n_1420),
.Y(n_3846)
);

OAI211xp5_ASAP7_75t_L g3847 ( 
.A1(n_3812),
.A2(n_1453),
.B(n_1472),
.C(n_1436),
.Y(n_3847)
);

OA21x2_ASAP7_75t_L g3848 ( 
.A1(n_3819),
.A2(n_1435),
.B(n_1430),
.Y(n_3848)
);

INVx3_ASAP7_75t_L g3849 ( 
.A(n_3773),
.Y(n_3849)
);

OAI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_3826),
.A2(n_1441),
.B1(n_1442),
.B2(n_1437),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3796),
.B(n_3813),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3792),
.B(n_1446),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3778),
.Y(n_3853)
);

OAI22xp5_ASAP7_75t_L g3854 ( 
.A1(n_3826),
.A2(n_1449),
.B1(n_1452),
.B2(n_1447),
.Y(n_3854)
);

AOI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3785),
.A2(n_1917),
.B1(n_1919),
.B2(n_1908),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3784),
.B(n_40),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3791),
.B(n_40),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3830),
.A2(n_1460),
.B1(n_1461),
.B2(n_1459),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3777),
.Y(n_3859)
);

AOI22xp5_ASAP7_75t_L g3860 ( 
.A1(n_3775),
.A2(n_1465),
.B1(n_1468),
.B2(n_1464),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3797),
.A2(n_1861),
.B1(n_1862),
.B2(n_1860),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3800),
.B(n_41),
.Y(n_3862)
);

OAI211xp5_ASAP7_75t_L g3863 ( 
.A1(n_3827),
.A2(n_1502),
.B(n_1515),
.C(n_1485),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3778),
.Y(n_3864)
);

OR2x2_ASAP7_75t_L g3865 ( 
.A(n_3838),
.B(n_3790),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3836),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3859),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3834),
.Y(n_3868)
);

AND2x4_ASAP7_75t_L g3869 ( 
.A(n_3851),
.B(n_3781),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3851),
.B(n_3800),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3845),
.B(n_3802),
.Y(n_3871)
);

AND2x4_ASAP7_75t_L g3872 ( 
.A(n_3849),
.B(n_3799),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3832),
.Y(n_3873)
);

OR2x2_ASAP7_75t_L g3874 ( 
.A(n_3842),
.B(n_3779),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_3852),
.B(n_3794),
.Y(n_3875)
);

BUFx6f_ASAP7_75t_L g3876 ( 
.A(n_3862),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3832),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3853),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3864),
.B(n_3788),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3849),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3840),
.B(n_3802),
.Y(n_3881)
);

OAI221xp5_ASAP7_75t_SL g3882 ( 
.A1(n_3855),
.A2(n_3816),
.B1(n_3815),
.B2(n_3814),
.C(n_3828),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3856),
.B(n_3774),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3857),
.B(n_3821),
.Y(n_3884)
);

INVx3_ASAP7_75t_L g3885 ( 
.A(n_3844),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3841),
.B(n_3811),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3839),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3843),
.B(n_3821),
.Y(n_3888)
);

OAI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3858),
.A2(n_3824),
.B1(n_3822),
.B2(n_3809),
.Y(n_3889)
);

NAND2x1p5_ASAP7_75t_L g3890 ( 
.A(n_3848),
.B(n_3825),
.Y(n_3890)
);

BUFx3_ASAP7_75t_L g3891 ( 
.A(n_3839),
.Y(n_3891)
);

AND2x4_ASAP7_75t_L g3892 ( 
.A(n_3860),
.B(n_3825),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3848),
.B(n_3806),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3863),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_L g3895 ( 
.A(n_3833),
.B(n_3829),
.Y(n_3895)
);

NOR2xp33_ASAP7_75t_L g3896 ( 
.A(n_3847),
.B(n_3810),
.Y(n_3896)
);

INVx3_ASAP7_75t_L g3897 ( 
.A(n_3835),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3870),
.B(n_3776),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3873),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3877),
.Y(n_3900)
);

INVxp67_ASAP7_75t_SL g3901 ( 
.A(n_3890),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3893),
.B(n_3837),
.Y(n_3902)
);

INVx2_ASAP7_75t_SL g3903 ( 
.A(n_3868),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3866),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3881),
.B(n_3787),
.Y(n_3905)
);

AOI22xp33_ASAP7_75t_L g3906 ( 
.A1(n_3897),
.A2(n_3831),
.B1(n_3861),
.B2(n_3820),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3867),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3871),
.B(n_3850),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3869),
.B(n_3820),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3878),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3879),
.Y(n_3911)
);

NOR2xp67_ASAP7_75t_L g3912 ( 
.A(n_3885),
.B(n_3854),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3886),
.B(n_3883),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3869),
.B(n_41),
.Y(n_3914)
);

AND2x4_ASAP7_75t_L g3915 ( 
.A(n_3872),
.B(n_43),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3884),
.B(n_42),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3891),
.B(n_1469),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3887),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3888),
.B(n_42),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3874),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3876),
.B(n_44),
.Y(n_3921)
);

OA21x2_ASAP7_75t_L g3922 ( 
.A1(n_3872),
.A2(n_3846),
.B(n_1478),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3896),
.B(n_1476),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3876),
.B(n_46),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3880),
.B(n_46),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3865),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3892),
.B(n_47),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3889),
.B(n_1487),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3875),
.B(n_50),
.Y(n_3929)
);

OR2x2_ASAP7_75t_L g3930 ( 
.A(n_3882),
.B(n_51),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3895),
.B(n_52),
.Y(n_3931)
);

BUFx3_ASAP7_75t_L g3932 ( 
.A(n_3894),
.Y(n_3932)
);

AOI33xp33_ASAP7_75t_L g3933 ( 
.A1(n_3906),
.A2(n_1499),
.A3(n_1491),
.B1(n_1500),
.B2(n_1495),
.B3(n_1488),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3926),
.B(n_52),
.Y(n_3934)
);

OAI33xp33_ASAP7_75t_L g3935 ( 
.A1(n_3930),
.A2(n_1506),
.A3(n_1503),
.B1(n_1507),
.B2(n_1504),
.B3(n_1501),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3903),
.B(n_55),
.Y(n_3936)
);

OR2x2_ASAP7_75t_L g3937 ( 
.A(n_3913),
.B(n_55),
.Y(n_3937)
);

NOR3xp33_ASAP7_75t_SL g3938 ( 
.A(n_3902),
.B(n_1512),
.C(n_1509),
.Y(n_3938)
);

OR2x2_ASAP7_75t_L g3939 ( 
.A(n_3920),
.B(n_56),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3899),
.Y(n_3940)
);

OAI33xp33_ASAP7_75t_L g3941 ( 
.A1(n_3917),
.A2(n_1529),
.A3(n_1516),
.B1(n_1535),
.B2(n_1528),
.B3(n_1513),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3899),
.Y(n_3942)
);

INVx1_ASAP7_75t_SL g3943 ( 
.A(n_3915),
.Y(n_3943)
);

NAND4xp25_ASAP7_75t_SL g3944 ( 
.A(n_3923),
.B(n_59),
.C(n_57),
.D(n_58),
.Y(n_3944)
);

INVx3_ASAP7_75t_L g3945 ( 
.A(n_3915),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3900),
.Y(n_3946)
);

OAI31xp33_ASAP7_75t_L g3947 ( 
.A1(n_3901),
.A2(n_60),
.A3(n_58),
.B(n_59),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3909),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3932),
.Y(n_3949)
);

AOI221xp5_ASAP7_75t_L g3950 ( 
.A1(n_3928),
.A2(n_1539),
.B1(n_1541),
.B2(n_1538),
.C(n_1537),
.Y(n_3950)
);

AOI33xp33_ASAP7_75t_L g3951 ( 
.A1(n_3931),
.A2(n_1557),
.A3(n_1544),
.B1(n_1559),
.B2(n_1555),
.B3(n_1543),
.Y(n_3951)
);

AOI22xp33_ASAP7_75t_L g3952 ( 
.A1(n_3922),
.A2(n_1567),
.B1(n_1568),
.B2(n_1562),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3900),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3904),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_3922),
.A2(n_1573),
.B1(n_1574),
.B2(n_1569),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3905),
.B(n_61),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3907),
.Y(n_3957)
);

OAI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3912),
.A2(n_1601),
.B1(n_1611),
.B2(n_1586),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3914),
.B(n_3911),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3898),
.B(n_62),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3916),
.B(n_62),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3910),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3918),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3918),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3919),
.B(n_63),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3945),
.B(n_3908),
.Y(n_3966)
);

NAND2x1_ASAP7_75t_SL g3967 ( 
.A(n_3945),
.B(n_3927),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3949),
.Y(n_3968)
);

BUFx2_ASAP7_75t_L g3969 ( 
.A(n_3943),
.Y(n_3969)
);

NAND2x1_ASAP7_75t_L g3970 ( 
.A(n_3960),
.B(n_3921),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3959),
.B(n_3924),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3953),
.Y(n_3972)
);

NOR2x1_ASAP7_75t_L g3973 ( 
.A(n_3958),
.B(n_3929),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3935),
.A2(n_3925),
.B1(n_1581),
.B2(n_1584),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3937),
.B(n_63),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3956),
.B(n_1576),
.Y(n_3976)
);

CKINVDCx16_ASAP7_75t_R g3977 ( 
.A(n_3936),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3947),
.B(n_1587),
.Y(n_3978)
);

INVx5_ASAP7_75t_L g3979 ( 
.A(n_3934),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3939),
.B(n_1588),
.Y(n_3980)
);

INVx2_ASAP7_75t_SL g3981 ( 
.A(n_3961),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3965),
.B(n_1590),
.Y(n_3982)
);

OR2x2_ASAP7_75t_L g3983 ( 
.A(n_3948),
.B(n_64),
.Y(n_3983)
);

HB1xp67_ASAP7_75t_L g3984 ( 
.A(n_3963),
.Y(n_3984)
);

OAI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3952),
.A2(n_1889),
.B(n_1886),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3962),
.B(n_64),
.Y(n_3986)
);

INVx1_ASAP7_75t_SL g3987 ( 
.A(n_3954),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3953),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3957),
.B(n_66),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3940),
.B(n_66),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3942),
.B(n_68),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3946),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3955),
.B(n_1596),
.Y(n_3993)
);

HB1xp67_ASAP7_75t_L g3994 ( 
.A(n_3964),
.Y(n_3994)
);

NOR2xp33_ASAP7_75t_SL g3995 ( 
.A(n_3944),
.B(n_1597),
.Y(n_3995)
);

INVxp67_ASAP7_75t_SL g3996 ( 
.A(n_3950),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3951),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3938),
.B(n_69),
.Y(n_3998)
);

HB1xp67_ASAP7_75t_L g3999 ( 
.A(n_3941),
.Y(n_3999)
);

BUFx2_ASAP7_75t_L g4000 ( 
.A(n_3933),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_L g4001 ( 
.A(n_3943),
.B(n_1598),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3945),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3945),
.B(n_69),
.Y(n_4003)
);

INVxp67_ASAP7_75t_L g4004 ( 
.A(n_3945),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3945),
.B(n_70),
.Y(n_4005)
);

INVxp33_ASAP7_75t_L g4006 ( 
.A(n_3959),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3943),
.B(n_71),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3945),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3945),
.B(n_72),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3945),
.B(n_72),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3984),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3967),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3988),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3977),
.B(n_1600),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3966),
.B(n_74),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3979),
.B(n_1603),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3969),
.B(n_75),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3971),
.B(n_76),
.Y(n_4018)
);

OR2x2_ASAP7_75t_L g4019 ( 
.A(n_3981),
.B(n_77),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3979),
.B(n_79),
.Y(n_4020)
);

OR2x2_ASAP7_75t_L g4021 ( 
.A(n_4004),
.B(n_81),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3988),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_SL g4023 ( 
.A1(n_3979),
.A2(n_1605),
.B1(n_1606),
.B2(n_1604),
.Y(n_4023)
);

INVx2_ASAP7_75t_L g4024 ( 
.A(n_4002),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_4006),
.B(n_82),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3972),
.Y(n_4026)
);

INVxp67_ASAP7_75t_L g4027 ( 
.A(n_3973),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_4008),
.Y(n_4028)
);

INVx1_ASAP7_75t_SL g4029 ( 
.A(n_4007),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3994),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3990),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3999),
.B(n_1608),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_3968),
.B(n_82),
.Y(n_4033)
);

INVxp67_ASAP7_75t_L g4034 ( 
.A(n_4003),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3991),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3970),
.B(n_83),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_4000),
.B(n_1609),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3996),
.A2(n_1855),
.B(n_1854),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3986),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_4005),
.B(n_1610),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3989),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_4009),
.B(n_1615),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_4010),
.B(n_84),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_4001),
.B(n_1616),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3992),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3997),
.B(n_1617),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3997),
.B(n_1618),
.Y(n_4047)
);

NAND2x1_ASAP7_75t_L g4048 ( 
.A(n_3983),
.B(n_84),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3987),
.B(n_3980),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3975),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3976),
.Y(n_4051)
);

INVxp67_ASAP7_75t_L g4052 ( 
.A(n_3995),
.Y(n_4052)
);

OR2x6_ASAP7_75t_L g4053 ( 
.A(n_3982),
.B(n_85),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_L g4054 ( 
.A(n_3978),
.B(n_1619),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3998),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3974),
.B(n_1623),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_SL g4057 ( 
.A1(n_3985),
.A2(n_85),
.B(n_86),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3993),
.B(n_86),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3967),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3977),
.B(n_1624),
.Y(n_4060)
);

AND2x4_ASAP7_75t_L g4061 ( 
.A(n_3979),
.B(n_88),
.Y(n_4061)
);

INVx3_ASAP7_75t_L g4062 ( 
.A(n_4002),
.Y(n_4062)
);

INVx2_ASAP7_75t_SL g4063 ( 
.A(n_3967),
.Y(n_4063)
);

OR2x2_ASAP7_75t_L g4064 ( 
.A(n_3969),
.B(n_89),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3977),
.B(n_1625),
.Y(n_4065)
);

INVxp67_ASAP7_75t_L g4066 ( 
.A(n_3969),
.Y(n_4066)
);

OAI211xp5_ASAP7_75t_L g4067 ( 
.A1(n_3967),
.A2(n_1628),
.B(n_1635),
.C(n_1633),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3984),
.Y(n_4068)
);

OR2x2_ASAP7_75t_L g4069 ( 
.A(n_3969),
.B(n_89),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3984),
.Y(n_4070)
);

OR2x2_ASAP7_75t_L g4071 ( 
.A(n_3969),
.B(n_90),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_3969),
.B(n_90),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3977),
.B(n_92),
.Y(n_4073)
);

INVxp67_ASAP7_75t_L g4074 ( 
.A(n_3969),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3977),
.B(n_1627),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_4012),
.B(n_1636),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_4066),
.B(n_93),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_4027),
.A2(n_1638),
.B1(n_1639),
.B2(n_1637),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4061),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_4074),
.B(n_93),
.Y(n_4080)
);

AOI321xp33_ASAP7_75t_L g4081 ( 
.A1(n_4059),
.A2(n_4070),
.A3(n_4068),
.B1(n_4011),
.B2(n_4055),
.C(n_4024),
.Y(n_4081)
);

INVxp33_ASAP7_75t_L g4082 ( 
.A(n_4073),
.Y(n_4082)
);

AND2x4_ASAP7_75t_SL g4083 ( 
.A(n_4061),
.B(n_94),
.Y(n_4083)
);

INVxp67_ASAP7_75t_L g4084 ( 
.A(n_4020),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4021),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4063),
.B(n_1641),
.Y(n_4086)
);

OR2x2_ASAP7_75t_L g4087 ( 
.A(n_4029),
.B(n_95),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_4019),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4017),
.B(n_1645),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_4064),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4069),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_4071),
.B(n_1646),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_4034),
.B(n_95),
.Y(n_4093)
);

INVx2_ASAP7_75t_SL g4094 ( 
.A(n_4062),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4072),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_4052),
.B(n_1647),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_4039),
.B(n_96),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_4015),
.B(n_1648),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4013),
.Y(n_4099)
);

OAI21xp33_ASAP7_75t_L g4100 ( 
.A1(n_4049),
.A2(n_4041),
.B(n_4035),
.Y(n_4100)
);

AOI22xp33_ASAP7_75t_L g4101 ( 
.A1(n_4031),
.A2(n_1652),
.B1(n_1653),
.B2(n_1651),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_4048),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4022),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_4050),
.B(n_96),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4025),
.Y(n_4105)
);

OR2x2_ASAP7_75t_L g4106 ( 
.A(n_4028),
.B(n_97),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4033),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_4030),
.B(n_4014),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4018),
.Y(n_4109)
);

AOI22x1_ASAP7_75t_L g4110 ( 
.A1(n_4036),
.A2(n_1658),
.B1(n_1659),
.B2(n_1655),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_4043),
.Y(n_4111)
);

INVx2_ASAP7_75t_SL g4112 ( 
.A(n_4053),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4026),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4051),
.B(n_1660),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4045),
.Y(n_4115)
);

AO22x1_ASAP7_75t_L g4116 ( 
.A1(n_4032),
.A2(n_4075),
.B1(n_4060),
.B2(n_4065),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4053),
.B(n_1664),
.Y(n_4117)
);

OAI21xp5_ASAP7_75t_SL g4118 ( 
.A1(n_4057),
.A2(n_4067),
.B(n_4023),
.Y(n_4118)
);

OR2x2_ASAP7_75t_L g4119 ( 
.A(n_4037),
.B(n_97),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_4054),
.B(n_1667),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_4046),
.B(n_1669),
.Y(n_4121)
);

INVx1_ASAP7_75t_SL g4122 ( 
.A(n_4058),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_4016),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4047),
.B(n_4040),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4042),
.Y(n_4125)
);

INVx1_ASAP7_75t_SL g4126 ( 
.A(n_4044),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_4038),
.B(n_1670),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_4056),
.A2(n_1672),
.B1(n_1675),
.B2(n_1671),
.Y(n_4128)
);

NAND2x1_ASAP7_75t_SL g4129 ( 
.A(n_4061),
.B(n_98),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_SL g4130 ( 
.A(n_4027),
.B(n_1678),
.Y(n_4130)
);

OAI32xp33_ASAP7_75t_L g4131 ( 
.A1(n_4027),
.A2(n_1685),
.A3(n_1688),
.B1(n_1687),
.B2(n_1684),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4061),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_4027),
.A2(n_1689),
.B1(n_1690),
.B2(n_1679),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_4027),
.A2(n_1699),
.B(n_1694),
.Y(n_4134)
);

INVxp67_ASAP7_75t_L g4135 ( 
.A(n_4073),
.Y(n_4135)
);

INVxp67_ASAP7_75t_L g4136 ( 
.A(n_4073),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4012),
.B(n_1702),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_4027),
.A2(n_1838),
.B(n_1834),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4061),
.Y(n_4139)
);

O2A1O1Ixp33_ASAP7_75t_SL g4140 ( 
.A1(n_4027),
.A2(n_101),
.B(n_98),
.C(n_99),
.Y(n_4140)
);

OAI33xp33_ASAP7_75t_L g4141 ( 
.A1(n_4027),
.A2(n_1712),
.A3(n_1708),
.B1(n_1713),
.B2(n_1709),
.B3(n_1707),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4061),
.Y(n_4142)
);

AOI22xp5_ASAP7_75t_L g4143 ( 
.A1(n_4027),
.A2(n_1717),
.B1(n_1719),
.B2(n_1715),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4061),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4012),
.B(n_1721),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_4027),
.B(n_1722),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4061),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4027),
.B(n_1724),
.Y(n_4148)
);

NAND2x1_ASAP7_75t_SL g4149 ( 
.A(n_4061),
.B(n_101),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4012),
.B(n_1725),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4027),
.B(n_1726),
.Y(n_4151)
);

INVx3_ASAP7_75t_L g4152 ( 
.A(n_4061),
.Y(n_4152)
);

OAI221xp5_ASAP7_75t_SL g4153 ( 
.A1(n_4027),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4027),
.B(n_1730),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4061),
.Y(n_4155)
);

HB1xp67_ASAP7_75t_L g4156 ( 
.A(n_4061),
.Y(n_4156)
);

OAI221xp5_ASAP7_75t_L g4157 ( 
.A1(n_4027),
.A2(n_1853),
.B1(n_1734),
.B2(n_1735),
.C(n_1733),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_4027),
.B(n_1732),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4061),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4061),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4027),
.B(n_1736),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4061),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4082),
.B(n_1739),
.Y(n_4163)
);

OR2x6_ASAP7_75t_L g4164 ( 
.A(n_4112),
.B(n_105),
.Y(n_4164)
);

OAI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_4135),
.A2(n_1744),
.B1(n_1746),
.B2(n_1741),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_4136),
.B(n_1754),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4152),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4156),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4102),
.B(n_1756),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4129),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_4152),
.Y(n_4171)
);

INVx2_ASAP7_75t_SL g4172 ( 
.A(n_4149),
.Y(n_4172)
);

AOI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4094),
.A2(n_1760),
.B1(n_1761),
.B2(n_1757),
.Y(n_4173)
);

NAND2x1p5_ASAP7_75t_L g4174 ( 
.A(n_4079),
.B(n_104),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_4084),
.B(n_1765),
.Y(n_4175)
);

NOR2xp33_ASAP7_75t_L g4176 ( 
.A(n_4132),
.B(n_1766),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_4139),
.B(n_1769),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4142),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4144),
.Y(n_4179)
);

OAI21xp33_ASAP7_75t_L g4180 ( 
.A1(n_4100),
.A2(n_1771),
.B(n_1770),
.Y(n_4180)
);

HB1xp67_ASAP7_75t_L g4181 ( 
.A(n_4147),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4155),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4159),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_4130),
.A2(n_1773),
.B1(n_1776),
.B2(n_1772),
.Y(n_4184)
);

AOI221xp5_ASAP7_75t_L g4185 ( 
.A1(n_4140),
.A2(n_1781),
.B1(n_1782),
.B2(n_1780),
.C(n_1777),
.Y(n_4185)
);

AOI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_4109),
.A2(n_1785),
.B1(n_1789),
.B2(n_1783),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4160),
.B(n_106),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4162),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_4111),
.B(n_1792),
.Y(n_4189)
);

OR2x2_ASAP7_75t_L g4190 ( 
.A(n_4090),
.B(n_106),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4077),
.Y(n_4191)
);

NAND3xp33_ASAP7_75t_L g4192 ( 
.A(n_4081),
.B(n_1863),
.C(n_1859),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4080),
.Y(n_4193)
);

HB1xp67_ASAP7_75t_L g4194 ( 
.A(n_4091),
.Y(n_4194)
);

INVx1_ASAP7_75t_SL g4195 ( 
.A(n_4083),
.Y(n_4195)
);

NAND3xp33_ASAP7_75t_L g4196 ( 
.A(n_4095),
.B(n_1898),
.C(n_1865),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_4098),
.B(n_1795),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4104),
.Y(n_4198)
);

INVxp67_ASAP7_75t_L g4199 ( 
.A(n_4087),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_4106),
.Y(n_4200)
);

OAI21xp33_ASAP7_75t_L g4201 ( 
.A1(n_4105),
.A2(n_1797),
.B(n_1796),
.Y(n_4201)
);

AOI21xp5_ASAP7_75t_L g4202 ( 
.A1(n_4118),
.A2(n_4138),
.B(n_4092),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4097),
.Y(n_4203)
);

NAND2x1_ASAP7_75t_L g4204 ( 
.A(n_4088),
.B(n_110),
.Y(n_4204)
);

INVx2_ASAP7_75t_SL g4205 ( 
.A(n_4093),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4107),
.Y(n_4206)
);

OAI32xp33_ASAP7_75t_L g4207 ( 
.A1(n_4122),
.A2(n_1807),
.A3(n_1811),
.B1(n_1804),
.B2(n_1801),
.Y(n_4207)
);

AOI221xp5_ASAP7_75t_L g4208 ( 
.A1(n_4153),
.A2(n_1814),
.B1(n_1816),
.B2(n_1813),
.C(n_1812),
.Y(n_4208)
);

OAI22xp5_ASAP7_75t_L g4209 ( 
.A1(n_4078),
.A2(n_1819),
.B1(n_1820),
.B2(n_1818),
.Y(n_4209)
);

CKINVDCx14_ASAP7_75t_R g4210 ( 
.A(n_4117),
.Y(n_4210)
);

AOI32xp33_ASAP7_75t_L g4211 ( 
.A1(n_4085),
.A2(n_1823),
.A3(n_1824),
.B1(n_1822),
.B2(n_1821),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4116),
.B(n_1828),
.Y(n_4212)
);

OAI22xp5_ASAP7_75t_L g4213 ( 
.A1(n_4143),
.A2(n_1844),
.B1(n_1846),
.B2(n_1833),
.Y(n_4213)
);

AOI32xp33_ASAP7_75t_L g4214 ( 
.A1(n_4133),
.A2(n_1907),
.A3(n_1921),
.B1(n_1857),
.B2(n_1851),
.Y(n_4214)
);

AOI22xp5_ASAP7_75t_L g4215 ( 
.A1(n_4126),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_4215)
);

OAI211xp5_ASAP7_75t_SL g4216 ( 
.A1(n_4108),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4076),
.B(n_114),
.Y(n_4217)
);

AOI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_4125),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.Y(n_4218)
);

OAI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_4134),
.A2(n_116),
.B(n_117),
.Y(n_4219)
);

A2O1A1Ixp33_ASAP7_75t_L g4220 ( 
.A1(n_4119),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_4220)
);

OR2x2_ASAP7_75t_L g4221 ( 
.A(n_4123),
.B(n_120),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4099),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4137),
.B(n_122),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4103),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4145),
.B(n_122),
.Y(n_4225)
);

O2A1O1Ixp33_ASAP7_75t_L g4226 ( 
.A1(n_4146),
.A2(n_985),
.B(n_986),
.C(n_984),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4124),
.B(n_123),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4150),
.B(n_123),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4114),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4113),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4115),
.Y(n_4231)
);

OA211x2_ASAP7_75t_L g4232 ( 
.A1(n_4096),
.A2(n_128),
.B(n_124),
.C(n_125),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4086),
.B(n_125),
.Y(n_4233)
);

AOI221x1_ASAP7_75t_L g4234 ( 
.A1(n_4148),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_4234)
);

NAND3xp33_ASAP7_75t_L g4235 ( 
.A(n_4151),
.B(n_130),
.C(n_131),
.Y(n_4235)
);

AOI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_4141),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_4236)
);

AOI22xp33_ASAP7_75t_L g4237 ( 
.A1(n_4154),
.A2(n_135),
.B1(n_132),
.B2(n_134),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4089),
.B(n_135),
.Y(n_4238)
);

OAI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_4158),
.A2(n_136),
.B(n_139),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4101),
.B(n_136),
.Y(n_4240)
);

INVx1_ASAP7_75t_SL g4241 ( 
.A(n_4110),
.Y(n_4241)
);

A2O1A1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_4161),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4127),
.B(n_141),
.Y(n_4243)
);

O2A1O1Ixp33_ASAP7_75t_L g4244 ( 
.A1(n_4131),
.A2(n_986),
.B(n_987),
.C(n_984),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4121),
.B(n_143),
.Y(n_4245)
);

AOI21xp33_ASAP7_75t_L g4246 ( 
.A1(n_4157),
.A2(n_4128),
.B(n_4120),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_4129),
.Y(n_4247)
);

NAND2xp33_ASAP7_75t_L g4248 ( 
.A(n_4102),
.B(n_144),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4156),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4156),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4079),
.B(n_144),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4152),
.B(n_145),
.Y(n_4252)
);

AOI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_4112),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4152),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4152),
.B(n_146),
.Y(n_4255)
);

OAI21xp33_ASAP7_75t_L g4256 ( 
.A1(n_4082),
.A2(n_147),
.B(n_148),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4082),
.B(n_149),
.Y(n_4257)
);

HB1xp67_ASAP7_75t_L g4258 ( 
.A(n_4102),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4152),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_4082),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_4152),
.B(n_151),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_4152),
.B(n_152),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_4152),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4156),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4152),
.Y(n_4265)
);

AOI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4112),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_4082),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4156),
.Y(n_4268)
);

OAI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_4112),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4152),
.B(n_156),
.Y(n_4270)
);

NAND2xp33_ASAP7_75t_L g4271 ( 
.A(n_4102),
.B(n_157),
.Y(n_4271)
);

AOI21xp33_ASAP7_75t_L g4272 ( 
.A1(n_4082),
.A2(n_988),
.B(n_983),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4156),
.Y(n_4273)
);

AND2x4_ASAP7_75t_L g4274 ( 
.A(n_4152),
.B(n_158),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4082),
.B(n_159),
.Y(n_4275)
);

OAI32xp33_ASAP7_75t_L g4276 ( 
.A1(n_4102),
.A2(n_163),
.A3(n_165),
.B1(n_162),
.B2(n_164),
.Y(n_4276)
);

OAI21xp33_ASAP7_75t_L g4277 ( 
.A1(n_4082),
.A2(n_160),
.B(n_162),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4082),
.B(n_165),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4156),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4152),
.Y(n_4280)
);

NAND3xp33_ASAP7_75t_L g4281 ( 
.A(n_4081),
.B(n_166),
.C(n_167),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4152),
.B(n_170),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4156),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4152),
.Y(n_4284)
);

OAI221xp5_ASAP7_75t_L g4285 ( 
.A1(n_4081),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.C(n_174),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4156),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4152),
.B(n_171),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4156),
.Y(n_4288)
);

OAI22xp33_ASAP7_75t_L g4289 ( 
.A1(n_4130),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_4289)
);

OAI32xp33_ASAP7_75t_L g4290 ( 
.A1(n_4102),
.A2(n_180),
.A3(n_184),
.B1(n_179),
.B2(n_181),
.Y(n_4290)
);

AOI22xp33_ASAP7_75t_L g4291 ( 
.A1(n_4082),
.A2(n_180),
.B1(n_177),
.B2(n_179),
.Y(n_4291)
);

AOI22xp5_ASAP7_75t_L g4292 ( 
.A1(n_4112),
.A2(n_186),
.B1(n_177),
.B2(n_185),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4156),
.Y(n_4293)
);

OR2x2_ASAP7_75t_L g4294 ( 
.A(n_4079),
.B(n_185),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4152),
.B(n_186),
.Y(n_4295)
);

AOI211xp5_ASAP7_75t_L g4296 ( 
.A1(n_4153),
.A2(n_191),
.B(n_188),
.C(n_189),
.Y(n_4296)
);

AOI322xp5_ASAP7_75t_L g4297 ( 
.A1(n_4112),
.A2(n_195),
.A3(n_194),
.B1(n_192),
.B2(n_188),
.C1(n_189),
.C2(n_193),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_4082),
.B(n_196),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4152),
.B(n_196),
.Y(n_4299)
);

AOI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4112),
.A2(n_201),
.B1(n_198),
.B2(n_200),
.Y(n_4300)
);

NAND3xp33_ASAP7_75t_L g4301 ( 
.A(n_4081),
.B(n_200),
.C(n_202),
.Y(n_4301)
);

NOR3xp33_ASAP7_75t_L g4302 ( 
.A(n_4100),
.B(n_203),
.C(n_204),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4082),
.B(n_204),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4156),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_4152),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4156),
.Y(n_4306)
);

AOI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_4112),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_4307)
);

OR2x2_ASAP7_75t_L g4308 ( 
.A(n_4079),
.B(n_205),
.Y(n_4308)
);

OAI32xp33_ASAP7_75t_L g4309 ( 
.A1(n_4102),
.A2(n_210),
.A3(n_214),
.B1(n_208),
.B2(n_212),
.Y(n_4309)
);

OR2x2_ASAP7_75t_L g4310 ( 
.A(n_4079),
.B(n_206),
.Y(n_4310)
);

INVxp67_ASAP7_75t_L g4311 ( 
.A(n_4102),
.Y(n_4311)
);

A2O1A1Ixp33_ASAP7_75t_L g4312 ( 
.A1(n_4081),
.A2(n_212),
.B(n_208),
.C(n_210),
.Y(n_4312)
);

O2A1O1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_4312),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_4313)
);

INVx3_ASAP7_75t_L g4314 ( 
.A(n_4274),
.Y(n_4314)
);

INVx2_ASAP7_75t_SL g4315 ( 
.A(n_4181),
.Y(n_4315)
);

AOI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_4281),
.A2(n_981),
.B1(n_982),
.B2(n_980),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4172),
.B(n_216),
.Y(n_4317)
);

AOI221x1_ASAP7_75t_L g4318 ( 
.A1(n_4301),
.A2(n_222),
.B1(n_217),
.B2(n_221),
.C(n_224),
.Y(n_4318)
);

AOI221xp5_ASAP7_75t_L g4319 ( 
.A1(n_4285),
.A2(n_990),
.B1(n_991),
.B2(n_989),
.C(n_988),
.Y(n_4319)
);

OAI32xp33_ASAP7_75t_L g4320 ( 
.A1(n_4170),
.A2(n_239),
.A3(n_247),
.B1(n_231),
.B2(n_222),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4258),
.Y(n_4321)
);

AOI21xp33_ASAP7_75t_SL g4322 ( 
.A1(n_4247),
.A2(n_994),
.B(n_993),
.Y(n_4322)
);

AOI221x1_ASAP7_75t_L g4323 ( 
.A1(n_4168),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.C(n_227),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4195),
.B(n_225),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_4248),
.A2(n_226),
.B(n_227),
.Y(n_4325)
);

OAI211xp5_ASAP7_75t_SL g4326 ( 
.A1(n_4199),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_4326)
);

INVxp67_ASAP7_75t_L g4327 ( 
.A(n_4164),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4167),
.Y(n_4328)
);

AOI22xp33_ASAP7_75t_L g4329 ( 
.A1(n_4210),
.A2(n_232),
.B1(n_228),
.B2(n_229),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4171),
.Y(n_4330)
);

NOR3xp33_ASAP7_75t_L g4331 ( 
.A(n_4246),
.B(n_232),
.C(n_233),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4254),
.B(n_234),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_4185),
.B(n_234),
.Y(n_4333)
);

INVxp67_ASAP7_75t_L g4334 ( 
.A(n_4164),
.Y(n_4334)
);

OA21x2_ASAP7_75t_L g4335 ( 
.A1(n_4192),
.A2(n_235),
.B(n_236),
.Y(n_4335)
);

OAI321xp33_ASAP7_75t_L g4336 ( 
.A1(n_4311),
.A2(n_237),
.A3(n_240),
.B1(n_235),
.B2(n_236),
.C(n_238),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4249),
.A2(n_242),
.B1(n_238),
.B2(n_241),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4259),
.B(n_243),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4263),
.Y(n_4339)
);

OAI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4302),
.A2(n_246),
.B(n_245),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4265),
.Y(n_4341)
);

OR2x2_ASAP7_75t_L g4342 ( 
.A(n_4280),
.B(n_244),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4284),
.B(n_244),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4305),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4250),
.Y(n_4345)
);

INVxp67_ASAP7_75t_L g4346 ( 
.A(n_4194),
.Y(n_4346)
);

OAI21xp33_ASAP7_75t_L g4347 ( 
.A1(n_4264),
.A2(n_245),
.B(n_246),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4268),
.B(n_973),
.Y(n_4348)
);

INVx2_ASAP7_75t_SL g4349 ( 
.A(n_4274),
.Y(n_4349)
);

INVxp33_ASAP7_75t_L g4350 ( 
.A(n_4174),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4273),
.B(n_4279),
.Y(n_4351)
);

AOI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_4283),
.A2(n_975),
.B1(n_976),
.B2(n_974),
.Y(n_4352)
);

AOI221xp5_ASAP7_75t_L g4353 ( 
.A1(n_4202),
.A2(n_977),
.B1(n_978),
.B2(n_974),
.C(n_973),
.Y(n_4353)
);

INVx2_ASAP7_75t_SL g4354 ( 
.A(n_4204),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4286),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4288),
.B(n_247),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4293),
.B(n_249),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4304),
.B(n_249),
.Y(n_4358)
);

INVxp67_ASAP7_75t_L g4359 ( 
.A(n_4271),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_4306),
.B(n_250),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4252),
.Y(n_4361)
);

AOI32xp33_ASAP7_75t_L g4362 ( 
.A1(n_4296),
.A2(n_254),
.A3(n_250),
.B1(n_253),
.B2(n_255),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_4212),
.A2(n_253),
.B(n_255),
.Y(n_4363)
);

OR2x2_ASAP7_75t_L g4364 ( 
.A(n_4178),
.B(n_257),
.Y(n_4364)
);

OAI22xp33_ASAP7_75t_L g4365 ( 
.A1(n_4234),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4365)
);

AOI222xp33_ASAP7_75t_L g4366 ( 
.A1(n_4179),
.A2(n_261),
.B1(n_263),
.B2(n_258),
.C1(n_259),
.C2(n_262),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4255),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4261),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4262),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4270),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4182),
.B(n_261),
.Y(n_4371)
);

NOR2xp33_ASAP7_75t_L g4372 ( 
.A(n_4256),
.B(n_262),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4282),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_4205),
.B(n_264),
.Y(n_4374)
);

OAI211xp5_ASAP7_75t_L g4375 ( 
.A1(n_4183),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_4375)
);

OAI322xp33_ASAP7_75t_L g4376 ( 
.A1(n_4188),
.A2(n_272),
.A3(n_270),
.B1(n_268),
.B2(n_266),
.C1(n_267),
.C2(n_269),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4229),
.A2(n_275),
.B1(n_270),
.B2(n_274),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4287),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4277),
.B(n_275),
.Y(n_4379)
);

AOI22xp33_ASAP7_75t_L g4380 ( 
.A1(n_4241),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_4380)
);

OAI221xp5_ASAP7_75t_SL g4381 ( 
.A1(n_4297),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.C(n_282),
.Y(n_4381)
);

OAI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4215),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_4382)
);

AOI211xp5_ASAP7_75t_L g4383 ( 
.A1(n_4276),
.A2(n_295),
.B(n_303),
.C(n_283),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4257),
.B(n_286),
.Y(n_4384)
);

OR4x1_ASAP7_75t_L g4385 ( 
.A(n_4206),
.B(n_288),
.C(n_286),
.D(n_287),
.Y(n_4385)
);

NAND4xp25_ASAP7_75t_L g4386 ( 
.A(n_4191),
.B(n_290),
.C(n_287),
.D(n_288),
.Y(n_4386)
);

OAI32xp33_ASAP7_75t_SL g4387 ( 
.A1(n_4235),
.A2(n_4196),
.A3(n_4193),
.B1(n_4203),
.B2(n_4230),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4198),
.B(n_4295),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4299),
.Y(n_4389)
);

AOI22xp33_ASAP7_75t_L g4390 ( 
.A1(n_4200),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4275),
.B(n_291),
.Y(n_4391)
);

AOI32xp33_ASAP7_75t_L g4392 ( 
.A1(n_4216),
.A2(n_296),
.A3(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4187),
.Y(n_4393)
);

AOI322xp5_ASAP7_75t_L g4394 ( 
.A1(n_4236),
.A2(n_301),
.A3(n_300),
.B1(n_298),
.B2(n_296),
.C1(n_297),
.C2(n_299),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4251),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4278),
.B(n_300),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4303),
.B(n_302),
.Y(n_4397)
);

OAI21xp5_ASAP7_75t_SL g4398 ( 
.A1(n_4226),
.A2(n_302),
.B(n_303),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_SL g4399 ( 
.A1(n_4169),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4294),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4308),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4260),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_4402)
);

INVx1_ASAP7_75t_SL g4403 ( 
.A(n_4310),
.Y(n_4403)
);

AOI22xp5_ASAP7_75t_L g4404 ( 
.A1(n_4298),
.A2(n_982),
.B1(n_989),
.B2(n_980),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4189),
.B(n_308),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4163),
.B(n_309),
.Y(n_4406)
);

A2O1A1Ixp33_ASAP7_75t_L g4407 ( 
.A1(n_4244),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4190),
.Y(n_4408)
);

INVx2_ASAP7_75t_SL g4409 ( 
.A(n_4221),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4227),
.Y(n_4410)
);

OAI21xp33_ASAP7_75t_L g4411 ( 
.A1(n_4231),
.A2(n_311),
.B(n_313),
.Y(n_4411)
);

A2O1A1Ixp33_ASAP7_75t_L g4412 ( 
.A1(n_4290),
.A2(n_316),
.B(n_313),
.C(n_315),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_4208),
.B(n_4289),
.Y(n_4413)
);

OAI31xp33_ASAP7_75t_L g4414 ( 
.A1(n_4220),
.A2(n_318),
.A3(n_315),
.B(n_317),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4176),
.A2(n_4180),
.B1(n_4201),
.B2(n_4269),
.Y(n_4415)
);

OAI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_4242),
.A2(n_319),
.B(n_318),
.Y(n_4416)
);

AOI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4175),
.A2(n_969),
.B1(n_971),
.B2(n_968),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4166),
.B(n_317),
.Y(n_4418)
);

INVx1_ASAP7_75t_SL g4419 ( 
.A(n_4233),
.Y(n_4419)
);

NAND2x1p5_ASAP7_75t_L g4420 ( 
.A(n_4253),
.B(n_321),
.Y(n_4420)
);

OR2x6_ASAP7_75t_L g4421 ( 
.A(n_4217),
.B(n_320),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4223),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4211),
.B(n_320),
.Y(n_4423)
);

INVx3_ASAP7_75t_SL g4424 ( 
.A(n_4240),
.Y(n_4424)
);

INVx1_ASAP7_75t_SL g4425 ( 
.A(n_4225),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_4228),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_L g4427 ( 
.A(n_4272),
.B(n_324),
.Y(n_4427)
);

OAI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4219),
.A2(n_326),
.B(n_325),
.Y(n_4428)
);

OR2x2_ASAP7_75t_L g4429 ( 
.A(n_4177),
.B(n_324),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4238),
.Y(n_4430)
);

INVxp33_ASAP7_75t_L g4431 ( 
.A(n_4243),
.Y(n_4431)
);

AOI222xp33_ASAP7_75t_L g4432 ( 
.A1(n_4346),
.A2(n_4359),
.B1(n_4334),
.B2(n_4327),
.C1(n_4321),
.C2(n_4413),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4354),
.B(n_4314),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4314),
.Y(n_4434)
);

OAI21xp5_ASAP7_75t_SL g4435 ( 
.A1(n_4350),
.A2(n_4292),
.B(n_4266),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4315),
.Y(n_4436)
);

AOI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4349),
.A2(n_4224),
.B1(n_4222),
.B2(n_4232),
.Y(n_4437)
);

NOR2xp33_ASAP7_75t_L g4438 ( 
.A(n_4424),
.B(n_4197),
.Y(n_4438)
);

AOI31xp33_ASAP7_75t_L g4439 ( 
.A1(n_4383),
.A2(n_4239),
.A3(n_4291),
.B(n_4267),
.Y(n_4439)
);

AOI211x1_ASAP7_75t_L g4440 ( 
.A1(n_4365),
.A2(n_4309),
.B(n_4207),
.C(n_4165),
.Y(n_4440)
);

AOI221xp5_ASAP7_75t_L g4441 ( 
.A1(n_4387),
.A2(n_4237),
.B1(n_4213),
.B2(n_4214),
.C(n_4300),
.Y(n_4441)
);

NOR3xp33_ASAP7_75t_L g4442 ( 
.A(n_4351),
.B(n_4245),
.C(n_4209),
.Y(n_4442)
);

NOR3xp33_ASAP7_75t_L g4443 ( 
.A(n_4333),
.B(n_4173),
.C(n_4186),
.Y(n_4443)
);

OAI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_4316),
.A2(n_4307),
.B1(n_4218),
.B2(n_4184),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4324),
.Y(n_4445)
);

NOR3xp33_ASAP7_75t_L g4446 ( 
.A(n_4395),
.B(n_325),
.C(n_326),
.Y(n_4446)
);

NAND3xp33_ASAP7_75t_SL g4447 ( 
.A(n_4403),
.B(n_329),
.C(n_328),
.Y(n_4447)
);

AOI211xp5_ASAP7_75t_L g4448 ( 
.A1(n_4381),
.A2(n_996),
.B(n_993),
.C(n_330),
.Y(n_4448)
);

AOI222xp33_ASAP7_75t_L g4449 ( 
.A1(n_4345),
.A2(n_330),
.B1(n_332),
.B2(n_327),
.C1(n_329),
.C2(n_331),
.Y(n_4449)
);

AOI221xp5_ASAP7_75t_L g4450 ( 
.A1(n_4313),
.A2(n_332),
.B1(n_327),
.B2(n_331),
.C(n_333),
.Y(n_4450)
);

NOR3xp33_ASAP7_75t_SL g4451 ( 
.A(n_4328),
.B(n_333),
.C(n_334),
.Y(n_4451)
);

INVxp67_ASAP7_75t_SL g4452 ( 
.A(n_4374),
.Y(n_4452)
);

OAI211xp5_ASAP7_75t_L g4453 ( 
.A1(n_4318),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_4453)
);

OR2x2_ASAP7_75t_L g4454 ( 
.A(n_4330),
.B(n_336),
.Y(n_4454)
);

AOI22xp5_ASAP7_75t_L g4455 ( 
.A1(n_4319),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_4455)
);

AOI221xp5_ASAP7_75t_L g4456 ( 
.A1(n_4398),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.C(n_342),
.Y(n_4456)
);

AND2x4_ASAP7_75t_L g4457 ( 
.A(n_4393),
.B(n_340),
.Y(n_4457)
);

NAND2xp33_ASAP7_75t_SL g4458 ( 
.A(n_4409),
.B(n_342),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_4407),
.A2(n_343),
.B(n_344),
.Y(n_4459)
);

AOI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4422),
.A2(n_347),
.B1(n_343),
.B2(n_345),
.Y(n_4460)
);

AOI221xp5_ASAP7_75t_L g4461 ( 
.A1(n_4339),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.C(n_351),
.Y(n_4461)
);

AOI211xp5_ASAP7_75t_L g4462 ( 
.A1(n_4341),
.A2(n_964),
.B(n_966),
.C(n_963),
.Y(n_4462)
);

OAI211xp5_ASAP7_75t_L g4463 ( 
.A1(n_4323),
.A2(n_353),
.B(n_349),
.C(n_352),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4322),
.B(n_352),
.Y(n_4464)
);

AOI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_4363),
.A2(n_354),
.B(n_355),
.Y(n_4465)
);

AOI21xp33_ASAP7_75t_L g4466 ( 
.A1(n_4431),
.A2(n_356),
.B(n_357),
.Y(n_4466)
);

AOI322xp5_ASAP7_75t_L g4467 ( 
.A1(n_4331),
.A2(n_968),
.A3(n_362),
.B1(n_359),
.B2(n_361),
.C1(n_356),
.C2(n_357),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4348),
.B(n_359),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_4348),
.Y(n_4469)
);

INVxp67_ASAP7_75t_SL g4470 ( 
.A(n_4420),
.Y(n_4470)
);

AND2x4_ASAP7_75t_L g4471 ( 
.A(n_4355),
.B(n_360),
.Y(n_4471)
);

OAI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_4380),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_4472)
);

AOI22xp5_ASAP7_75t_L g4473 ( 
.A1(n_4344),
.A2(n_366),
.B1(n_363),
.B2(n_365),
.Y(n_4473)
);

NAND4xp25_ASAP7_75t_L g4474 ( 
.A(n_4419),
.B(n_369),
.C(n_366),
.D(n_368),
.Y(n_4474)
);

NAND4xp25_ASAP7_75t_SL g4475 ( 
.A(n_4362),
.B(n_370),
.C(n_368),
.D(n_369),
.Y(n_4475)
);

NAND3xp33_ASAP7_75t_SL g4476 ( 
.A(n_4414),
.B(n_373),
.C(n_372),
.Y(n_4476)
);

OAI211xp5_ASAP7_75t_L g4477 ( 
.A1(n_4392),
.A2(n_375),
.B(n_371),
.C(n_374),
.Y(n_4477)
);

OAI221xp5_ASAP7_75t_L g4478 ( 
.A1(n_4340),
.A2(n_377),
.B1(n_371),
.B2(n_376),
.C(n_378),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_SL g4479 ( 
.A(n_4336),
.B(n_377),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4325),
.A2(n_378),
.B(n_379),
.Y(n_4480)
);

AOI211xp5_ASAP7_75t_SL g4481 ( 
.A1(n_4400),
.A2(n_383),
.B(n_380),
.C(n_382),
.Y(n_4481)
);

AOI221xp5_ASAP7_75t_L g4482 ( 
.A1(n_4401),
.A2(n_385),
.B1(n_380),
.B2(n_383),
.C(n_386),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_SL g4483 ( 
.A(n_4412),
.B(n_385),
.Y(n_4483)
);

AOI222xp33_ASAP7_75t_L g4484 ( 
.A1(n_4353),
.A2(n_391),
.B1(n_393),
.B2(n_387),
.C1(n_388),
.C2(n_392),
.Y(n_4484)
);

AOI21xp33_ASAP7_75t_L g4485 ( 
.A1(n_4388),
.A2(n_4408),
.B(n_4410),
.Y(n_4485)
);

AOI21xp33_ASAP7_75t_L g4486 ( 
.A1(n_4425),
.A2(n_387),
.B(n_388),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4396),
.Y(n_4487)
);

AOI211xp5_ASAP7_75t_L g4488 ( 
.A1(n_4382),
.A2(n_971),
.B(n_972),
.C(n_967),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4394),
.B(n_391),
.Y(n_4489)
);

NAND3xp33_ASAP7_75t_L g4490 ( 
.A(n_4366),
.B(n_393),
.C(n_394),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4418),
.B(n_4399),
.Y(n_4491)
);

NOR2xp33_ASAP7_75t_L g4492 ( 
.A(n_4347),
.B(n_394),
.Y(n_4492)
);

AOI221xp5_ASAP7_75t_L g4493 ( 
.A1(n_4376),
.A2(n_4320),
.B1(n_4416),
.B2(n_4367),
.C(n_4368),
.Y(n_4493)
);

OAI211xp5_ASAP7_75t_SL g4494 ( 
.A1(n_4361),
.A2(n_399),
.B(n_396),
.C(n_398),
.Y(n_4494)
);

AOI221x1_ASAP7_75t_L g4495 ( 
.A1(n_4356),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.C(n_401),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4428),
.A2(n_401),
.B(n_402),
.Y(n_4496)
);

AOI222xp33_ASAP7_75t_L g4497 ( 
.A1(n_4369),
.A2(n_404),
.B1(n_406),
.B2(n_402),
.C1(n_403),
.C2(n_405),
.Y(n_4497)
);

NOR2xp33_ASAP7_75t_L g4498 ( 
.A(n_4411),
.B(n_404),
.Y(n_4498)
);

O2A1O1Ixp5_ASAP7_75t_SL g4499 ( 
.A1(n_4370),
.A2(n_4378),
.B(n_4389),
.C(n_4373),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_SL g4500 ( 
.A(n_4317),
.B(n_407),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4421),
.B(n_407),
.Y(n_4501)
);

AOI221xp5_ASAP7_75t_L g4502 ( 
.A1(n_4326),
.A2(n_411),
.B1(n_408),
.B2(n_410),
.C(n_412),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4342),
.Y(n_4503)
);

AOI222xp33_ASAP7_75t_L g4504 ( 
.A1(n_4402),
.A2(n_412),
.B1(n_414),
.B2(n_410),
.C1(n_411),
.C2(n_413),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_4415),
.A2(n_421),
.B1(n_413),
.B2(n_416),
.Y(n_4505)
);

AOI22xp5_ASAP7_75t_L g4506 ( 
.A1(n_4430),
.A2(n_427),
.B1(n_421),
.B2(n_422),
.Y(n_4506)
);

OAI21xp33_ASAP7_75t_L g4507 ( 
.A1(n_4426),
.A2(n_427),
.B(n_428),
.Y(n_4507)
);

NAND4xp25_ASAP7_75t_L g4508 ( 
.A(n_4357),
.B(n_431),
.C(n_429),
.D(n_430),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4364),
.Y(n_4509)
);

OAI22xp33_ASAP7_75t_L g4510 ( 
.A1(n_4386),
.A2(n_432),
.B1(n_429),
.B2(n_431),
.Y(n_4510)
);

AOI32xp33_ASAP7_75t_L g4511 ( 
.A1(n_4372),
.A2(n_435),
.A3(n_433),
.B1(n_434),
.B2(n_436),
.Y(n_4511)
);

AOI221x1_ASAP7_75t_L g4512 ( 
.A1(n_4358),
.A2(n_437),
.B1(n_433),
.B2(n_434),
.C(n_438),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4384),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_4332),
.B(n_438),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4391),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_4337),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_L g4517 ( 
.A1(n_4335),
.A2(n_444),
.B1(n_439),
.B2(n_441),
.Y(n_4517)
);

OAI21xp33_ASAP7_75t_L g4518 ( 
.A1(n_4360),
.A2(n_444),
.B(n_445),
.Y(n_4518)
);

NAND4xp25_ASAP7_75t_L g4519 ( 
.A(n_4338),
.B(n_449),
.C(n_446),
.D(n_447),
.Y(n_4519)
);

OAI21xp33_ASAP7_75t_L g4520 ( 
.A1(n_4343),
.A2(n_446),
.B(n_447),
.Y(n_4520)
);

NAND3xp33_ASAP7_75t_L g4521 ( 
.A(n_4335),
.B(n_449),
.C(n_450),
.Y(n_4521)
);

NAND3xp33_ASAP7_75t_L g4522 ( 
.A(n_4375),
.B(n_450),
.C(n_452),
.Y(n_4522)
);

INVx2_ASAP7_75t_SL g4523 ( 
.A(n_4421),
.Y(n_4523)
);

OAI21xp33_ASAP7_75t_SL g4524 ( 
.A1(n_4371),
.A2(n_452),
.B(n_453),
.Y(n_4524)
);

AOI221xp5_ASAP7_75t_L g4525 ( 
.A1(n_4385),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.C(n_458),
.Y(n_4525)
);

AOI21xp33_ASAP7_75t_L g4526 ( 
.A1(n_4423),
.A2(n_455),
.B(n_457),
.Y(n_4526)
);

OAI222xp33_ASAP7_75t_L g4527 ( 
.A1(n_4352),
.A2(n_992),
.B1(n_978),
.B2(n_990),
.C1(n_977),
.C2(n_464),
.Y(n_4527)
);

NOR2xp33_ASAP7_75t_L g4528 ( 
.A(n_4397),
.B(n_459),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4379),
.B(n_459),
.Y(n_4529)
);

OAI21xp5_ASAP7_75t_L g4530 ( 
.A1(n_4427),
.A2(n_461),
.B(n_464),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4329),
.B(n_465),
.Y(n_4531)
);

AOI321xp33_ASAP7_75t_L g4532 ( 
.A1(n_4390),
.A2(n_470),
.A3(n_472),
.B1(n_466),
.B2(n_467),
.C(n_471),
.Y(n_4532)
);

OA22x2_ASAP7_75t_L g4533 ( 
.A1(n_4404),
.A2(n_472),
.B1(n_466),
.B2(n_470),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4405),
.B(n_4406),
.Y(n_4534)
);

OAI22xp5_ASAP7_75t_L g4535 ( 
.A1(n_4377),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4429),
.Y(n_4536)
);

OAI221xp5_ASAP7_75t_SL g4537 ( 
.A1(n_4417),
.A2(n_477),
.B1(n_474),
.B2(n_476),
.C(n_479),
.Y(n_4537)
);

AOI311xp33_ASAP7_75t_L g4538 ( 
.A1(n_4321),
.A2(n_481),
.A3(n_477),
.B(n_479),
.C(n_483),
.Y(n_4538)
);

AOI222xp33_ASAP7_75t_L g4539 ( 
.A1(n_4346),
.A2(n_485),
.B1(n_489),
.B2(n_481),
.C1(n_483),
.C2(n_487),
.Y(n_4539)
);

OAI21xp33_ASAP7_75t_L g4540 ( 
.A1(n_4350),
.A2(n_487),
.B(n_489),
.Y(n_4540)
);

OAI221xp5_ASAP7_75t_L g4541 ( 
.A1(n_4327),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.C(n_493),
.Y(n_4541)
);

A2O1A1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_4313),
.A2(n_495),
.B(n_492),
.C(n_494),
.Y(n_4542)
);

NAND3x2_ASAP7_75t_L g4543 ( 
.A(n_4321),
.B(n_494),
.C(n_496),
.Y(n_4543)
);

AOI322xp5_ASAP7_75t_L g4544 ( 
.A1(n_4413),
.A2(n_502),
.A3(n_501),
.B1(n_498),
.B2(n_496),
.C1(n_497),
.C2(n_499),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4314),
.Y(n_4545)
);

OAI21xp33_ASAP7_75t_L g4546 ( 
.A1(n_4350),
.A2(n_497),
.B(n_498),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4327),
.A2(n_499),
.B(n_503),
.Y(n_4547)
);

OAI22xp5_ASAP7_75t_L g4548 ( 
.A1(n_4359),
.A2(n_508),
.B1(n_503),
.B2(n_507),
.Y(n_4548)
);

NOR2xp33_ASAP7_75t_L g4549 ( 
.A(n_4354),
.B(n_507),
.Y(n_4549)
);

AOI21xp5_ASAP7_75t_L g4550 ( 
.A1(n_4354),
.A2(n_509),
.B(n_511),
.Y(n_4550)
);

AOI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_4354),
.A2(n_511),
.B(n_514),
.Y(n_4551)
);

AND4x1_ASAP7_75t_L g4552 ( 
.A(n_4323),
.B(n_516),
.C(n_514),
.D(n_515),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_4354),
.B(n_519),
.Y(n_4553)
);

AOI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_4354),
.A2(n_520),
.B(n_521),
.Y(n_4554)
);

NOR2xp33_ASAP7_75t_L g4555 ( 
.A(n_4354),
.B(n_520),
.Y(n_4555)
);

OAI21xp5_ASAP7_75t_L g4556 ( 
.A1(n_4327),
.A2(n_522),
.B(n_523),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_4354),
.A2(n_522),
.B(n_524),
.Y(n_4557)
);

O2A1O1Ixp5_ASAP7_75t_L g4558 ( 
.A1(n_4350),
.A2(n_530),
.B(n_525),
.C(n_529),
.Y(n_4558)
);

NOR3xp33_ASAP7_75t_L g4559 ( 
.A(n_4327),
.B(n_529),
.C(n_530),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_4350),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_4560)
);

AOI221xp5_ASAP7_75t_L g4561 ( 
.A1(n_4387),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.C(n_535),
.Y(n_4561)
);

NOR3xp33_ASAP7_75t_L g4562 ( 
.A(n_4327),
.B(n_534),
.C(n_535),
.Y(n_4562)
);

NAND3xp33_ASAP7_75t_SL g4563 ( 
.A(n_4350),
.B(n_537),
.C(n_539),
.Y(n_4563)
);

NOR4xp25_ASAP7_75t_L g4564 ( 
.A(n_4327),
.B(n_542),
.C(n_540),
.D(n_541),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4354),
.A2(n_540),
.B(n_541),
.Y(n_4565)
);

OR2x2_ASAP7_75t_L g4566 ( 
.A(n_4349),
.B(n_542),
.Y(n_4566)
);

AOI21xp5_ASAP7_75t_L g4567 ( 
.A1(n_4354),
.A2(n_543),
.B(n_544),
.Y(n_4567)
);

AOI221xp5_ASAP7_75t_L g4568 ( 
.A1(n_4387),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.C(n_546),
.Y(n_4568)
);

OAI221xp5_ASAP7_75t_SL g4569 ( 
.A1(n_4327),
.A2(n_548),
.B1(n_545),
.B2(n_547),
.C(n_549),
.Y(n_4569)
);

AOI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4327),
.A2(n_553),
.B1(n_549),
.B2(n_552),
.Y(n_4570)
);

AOI221x1_ASAP7_75t_L g4571 ( 
.A1(n_4331),
.A2(n_556),
.B1(n_552),
.B2(n_554),
.C(n_557),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_4354),
.A2(n_557),
.B(n_558),
.Y(n_4572)
);

NAND4xp25_ASAP7_75t_L g4573 ( 
.A(n_4351),
.B(n_967),
.C(n_560),
.D(n_558),
.Y(n_4573)
);

NAND3xp33_ASAP7_75t_L g4574 ( 
.A(n_4346),
.B(n_559),
.C(n_561),
.Y(n_4574)
);

AOI22xp33_ASAP7_75t_L g4575 ( 
.A1(n_4350),
.A2(n_562),
.B1(n_559),
.B2(n_561),
.Y(n_4575)
);

OAI221xp5_ASAP7_75t_L g4576 ( 
.A1(n_4327),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.C(n_566),
.Y(n_4576)
);

O2A1O1Ixp33_ASAP7_75t_SL g4577 ( 
.A1(n_4365),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_4577)
);

AOI22xp33_ASAP7_75t_L g4578 ( 
.A1(n_4350),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_4578)
);

OAI211xp5_ASAP7_75t_L g4579 ( 
.A1(n_4318),
.A2(n_570),
.B(n_568),
.C(n_569),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4359),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.Y(n_4580)
);

INVx2_ASAP7_75t_SL g4581 ( 
.A(n_4469),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4433),
.Y(n_4582)
);

AOI21xp33_ASAP7_75t_L g4583 ( 
.A1(n_4432),
.A2(n_4523),
.B(n_4470),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4436),
.B(n_571),
.Y(n_4584)
);

OAI21xp5_ASAP7_75t_L g4585 ( 
.A1(n_4499),
.A2(n_573),
.B(n_574),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4434),
.B(n_574),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4545),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4566),
.Y(n_4588)
);

OAI22xp5_ASAP7_75t_L g4589 ( 
.A1(n_4437),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_4589)
);

INVx1_ASAP7_75t_SL g4590 ( 
.A(n_4458),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4481),
.B(n_575),
.Y(n_4591)
);

NAND3xp33_ASAP7_75t_SL g4592 ( 
.A(n_4552),
.B(n_576),
.C(n_578),
.Y(n_4592)
);

AOI32xp33_ASAP7_75t_L g4593 ( 
.A1(n_4561),
.A2(n_581),
.A3(n_578),
.B1(n_580),
.B2(n_582),
.Y(n_4593)
);

AOI321xp33_ASAP7_75t_L g4594 ( 
.A1(n_4438),
.A2(n_584),
.A3(n_587),
.B1(n_580),
.B2(n_581),
.C(n_585),
.Y(n_4594)
);

OAI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4455),
.A2(n_590),
.B1(n_587),
.B2(n_588),
.Y(n_4595)
);

O2A1O1Ixp33_ASAP7_75t_SL g4596 ( 
.A1(n_4463),
.A2(n_592),
.B(n_588),
.C(n_590),
.Y(n_4596)
);

AOI21xp33_ASAP7_75t_L g4597 ( 
.A1(n_4439),
.A2(n_966),
.B(n_592),
.Y(n_4597)
);

AOI21xp33_ASAP7_75t_R g4598 ( 
.A1(n_4487),
.A2(n_593),
.B(n_594),
.Y(n_4598)
);

O2A1O1Ixp33_ASAP7_75t_L g4599 ( 
.A1(n_4479),
.A2(n_596),
.B(n_593),
.C(n_595),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4564),
.B(n_596),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4501),
.Y(n_4601)
);

AOI321xp33_ASAP7_75t_L g4602 ( 
.A1(n_4485),
.A2(n_964),
.A3(n_600),
.B1(n_603),
.B2(n_597),
.C(n_598),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4553),
.Y(n_4603)
);

O2A1O1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_4577),
.A2(n_4542),
.B(n_4447),
.C(n_4453),
.Y(n_4604)
);

OAI322xp33_ASAP7_75t_L g4605 ( 
.A1(n_4483),
.A2(n_605),
.A3(n_604),
.B1(n_600),
.B2(n_597),
.C1(n_598),
.C2(n_602),
.Y(n_4605)
);

NOR2xp67_ASAP7_75t_L g4606 ( 
.A(n_4521),
.B(n_602),
.Y(n_4606)
);

OAI221xp5_ASAP7_75t_L g4607 ( 
.A1(n_4568),
.A2(n_608),
.B1(n_604),
.B2(n_607),
.C(n_609),
.Y(n_4607)
);

OAI221xp5_ASAP7_75t_L g4608 ( 
.A1(n_4435),
.A2(n_611),
.B1(n_608),
.B2(n_610),
.C(n_612),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4468),
.Y(n_4609)
);

AOI21xp5_ASAP7_75t_L g4610 ( 
.A1(n_4465),
.A2(n_610),
.B(n_611),
.Y(n_4610)
);

OAI321xp33_ASAP7_75t_L g4611 ( 
.A1(n_4493),
.A2(n_614),
.A3(n_616),
.B1(n_612),
.B2(n_613),
.C(n_615),
.Y(n_4611)
);

A2O1A1Ixp33_ASAP7_75t_L g4612 ( 
.A1(n_4558),
.A2(n_963),
.B(n_617),
.C(n_613),
.Y(n_4612)
);

AOI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4475),
.A2(n_618),
.B1(n_616),
.B2(n_617),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4457),
.Y(n_4614)
);

NOR2xp33_ASAP7_75t_SL g4615 ( 
.A(n_4569),
.B(n_620),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4549),
.B(n_621),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_SL g4617 ( 
.A(n_4452),
.B(n_962),
.Y(n_4617)
);

OAI221xp5_ASAP7_75t_L g4618 ( 
.A1(n_4524),
.A2(n_624),
.B1(n_621),
.B2(n_623),
.C(n_625),
.Y(n_4618)
);

OAI211xp5_ASAP7_75t_L g4619 ( 
.A1(n_4579),
.A2(n_629),
.B(n_624),
.C(n_627),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4451),
.B(n_627),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4555),
.B(n_630),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4457),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4471),
.Y(n_4623)
);

OAI21xp33_ASAP7_75t_L g4624 ( 
.A1(n_4491),
.A2(n_630),
.B(n_631),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4503),
.B(n_632),
.Y(n_4625)
);

OAI21xp33_ASAP7_75t_SL g4626 ( 
.A1(n_4441),
.A2(n_632),
.B(n_633),
.Y(n_4626)
);

AOI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4444),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.C(n_637),
.Y(n_4627)
);

NOR2xp67_ASAP7_75t_L g4628 ( 
.A(n_4563),
.B(n_635),
.Y(n_4628)
);

AOI222xp33_ASAP7_75t_L g4629 ( 
.A1(n_4476),
.A2(n_639),
.B1(n_642),
.B2(n_636),
.C1(n_638),
.C2(n_640),
.Y(n_4629)
);

AOI21xp5_ASAP7_75t_L g4630 ( 
.A1(n_4550),
.A2(n_638),
.B(n_642),
.Y(n_4630)
);

AOI22xp5_ASAP7_75t_L g4631 ( 
.A1(n_4477),
.A2(n_648),
.B1(n_643),
.B2(n_647),
.Y(n_4631)
);

OAI22xp5_ASAP7_75t_SL g4632 ( 
.A1(n_4440),
.A2(n_4517),
.B1(n_4522),
.B2(n_4490),
.Y(n_4632)
);

OAI22xp5_ASAP7_75t_L g4633 ( 
.A1(n_4543),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_4633)
);

AOI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_4443),
.A2(n_652),
.B1(n_649),
.B2(n_650),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4471),
.Y(n_4635)
);

AOI22xp5_ASAP7_75t_L g4636 ( 
.A1(n_4442),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_4636)
);

OAI21xp33_ASAP7_75t_SL g4637 ( 
.A1(n_4509),
.A2(n_653),
.B(n_655),
.Y(n_4637)
);

OAI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4448),
.A2(n_661),
.B1(n_656),
.B2(n_659),
.Y(n_4638)
);

AOI322xp5_ASAP7_75t_L g4639 ( 
.A1(n_4489),
.A2(n_656),
.A3(n_659),
.B1(n_662),
.B2(n_663),
.C1(n_665),
.C2(n_666),
.Y(n_4639)
);

NOR2xp33_ASAP7_75t_L g4640 ( 
.A(n_4573),
.B(n_662),
.Y(n_4640)
);

O2A1O1Ixp33_ASAP7_75t_L g4641 ( 
.A1(n_4527),
.A2(n_670),
.B(n_667),
.C(n_668),
.Y(n_4641)
);

OAI221xp5_ASAP7_75t_SL g4642 ( 
.A1(n_4445),
.A2(n_671),
.B1(n_667),
.B2(n_668),
.C(n_672),
.Y(n_4642)
);

OAI21xp5_ASAP7_75t_SL g4643 ( 
.A1(n_4459),
.A2(n_671),
.B(n_672),
.Y(n_4643)
);

AOI221xp5_ASAP7_75t_L g4644 ( 
.A1(n_4525),
.A2(n_676),
.B1(n_674),
.B2(n_675),
.C(n_677),
.Y(n_4644)
);

OAI22xp5_ASAP7_75t_L g4645 ( 
.A1(n_4560),
.A2(n_677),
.B1(n_674),
.B2(n_676),
.Y(n_4645)
);

AOI21xp33_ASAP7_75t_L g4646 ( 
.A1(n_4534),
.A2(n_678),
.B(n_679),
.Y(n_4646)
);

OAI211xp5_ASAP7_75t_L g4647 ( 
.A1(n_4571),
.A2(n_681),
.B(n_679),
.C(n_680),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4454),
.Y(n_4648)
);

NOR2xp33_ASAP7_75t_L g4649 ( 
.A(n_4540),
.B(n_682),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4551),
.B(n_684),
.Y(n_4650)
);

AOI221xp5_ASAP7_75t_L g4651 ( 
.A1(n_4526),
.A2(n_688),
.B1(n_685),
.B2(n_686),
.C(n_689),
.Y(n_4651)
);

OAI31xp33_ASAP7_75t_L g4652 ( 
.A1(n_4494),
.A2(n_690),
.A3(n_688),
.B(n_689),
.Y(n_4652)
);

AOI22xp5_ASAP7_75t_L g4653 ( 
.A1(n_4510),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4464),
.Y(n_4654)
);

HB1xp67_ASAP7_75t_L g4655 ( 
.A(n_4533),
.Y(n_4655)
);

AOI322xp5_ASAP7_75t_L g4656 ( 
.A1(n_4456),
.A2(n_692),
.A3(n_693),
.B1(n_695),
.B2(n_696),
.C1(n_698),
.C2(n_699),
.Y(n_4656)
);

AOI221xp5_ASAP7_75t_L g4657 ( 
.A1(n_4450),
.A2(n_4502),
.B1(n_4472),
.B2(n_4516),
.C(n_4486),
.Y(n_4657)
);

HB1xp67_ASAP7_75t_L g4658 ( 
.A(n_4547),
.Y(n_4658)
);

OAI221xp5_ASAP7_75t_L g4659 ( 
.A1(n_4511),
.A2(n_698),
.B1(n_695),
.B2(n_696),
.C(n_700),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4554),
.B(n_700),
.Y(n_4660)
);

AOI21xp33_ASAP7_75t_SL g4661 ( 
.A1(n_4484),
.A2(n_701),
.B(n_702),
.Y(n_4661)
);

NOR2x1_ASAP7_75t_L g4662 ( 
.A(n_4474),
.B(n_701),
.Y(n_4662)
);

OAI211xp5_ASAP7_75t_SL g4663 ( 
.A1(n_4536),
.A2(n_706),
.B(n_702),
.C(n_704),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4513),
.Y(n_4664)
);

AOI22xp33_ASAP7_75t_SL g4665 ( 
.A1(n_4515),
.A2(n_707),
.B1(n_704),
.B2(n_706),
.Y(n_4665)
);

O2A1O1Ixp5_ASAP7_75t_SL g4666 ( 
.A1(n_4500),
.A2(n_710),
.B(n_708),
.C(n_709),
.Y(n_4666)
);

OAI221xp5_ASAP7_75t_L g4667 ( 
.A1(n_4532),
.A2(n_4530),
.B1(n_4488),
.B2(n_4546),
.C(n_4556),
.Y(n_4667)
);

NOR3x1_ASAP7_75t_L g4668 ( 
.A(n_4478),
.B(n_708),
.C(n_710),
.Y(n_4668)
);

INVxp33_ASAP7_75t_SL g4669 ( 
.A(n_4655),
.Y(n_4669)
);

OAI21xp5_ASAP7_75t_SL g4670 ( 
.A1(n_4583),
.A2(n_4496),
.B(n_4480),
.Y(n_4670)
);

NOR2x1_ASAP7_75t_L g4671 ( 
.A(n_4585),
.B(n_4592),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4596),
.A2(n_4565),
.B(n_4557),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4614),
.Y(n_4673)
);

AOI22xp5_ASAP7_75t_L g4674 ( 
.A1(n_4632),
.A2(n_4562),
.B1(n_4559),
.B2(n_4492),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4622),
.Y(n_4675)
);

A2O1A1Ixp33_ASAP7_75t_L g4676 ( 
.A1(n_4604),
.A2(n_4544),
.B(n_4572),
.C(n_4567),
.Y(n_4676)
);

OAI21xp5_ASAP7_75t_L g4677 ( 
.A1(n_4628),
.A2(n_4574),
.B(n_4514),
.Y(n_4677)
);

AOI211xp5_ASAP7_75t_SL g4678 ( 
.A1(n_4611),
.A2(n_4537),
.B(n_4466),
.C(n_4518),
.Y(n_4678)
);

OAI211xp5_ASAP7_75t_L g4679 ( 
.A1(n_4626),
.A2(n_4512),
.B(n_4495),
.C(n_4539),
.Y(n_4679)
);

OAI211xp5_ASAP7_75t_SL g4680 ( 
.A1(n_4582),
.A2(n_4467),
.B(n_4520),
.C(n_4504),
.Y(n_4680)
);

AOI21x1_ASAP7_75t_L g4681 ( 
.A1(n_4623),
.A2(n_4635),
.B(n_4600),
.Y(n_4681)
);

OA211x2_ASAP7_75t_L g4682 ( 
.A1(n_4617),
.A2(n_4507),
.B(n_4498),
.C(n_4528),
.Y(n_4682)
);

AOI211x1_ASAP7_75t_SL g4683 ( 
.A1(n_4589),
.A2(n_4535),
.B(n_4505),
.C(n_4548),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_SL g4684 ( 
.A(n_4602),
.B(n_4538),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4581),
.Y(n_4685)
);

AOI221xp5_ASAP7_75t_L g4686 ( 
.A1(n_4597),
.A2(n_4446),
.B1(n_4461),
.B2(n_4482),
.C(n_4580),
.Y(n_4686)
);

AOI21xp5_ASAP7_75t_L g4687 ( 
.A1(n_4610),
.A2(n_4529),
.B(n_4531),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4584),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4620),
.Y(n_4689)
);

OAI22xp33_ASAP7_75t_L g4690 ( 
.A1(n_4615),
.A2(n_4508),
.B1(n_4570),
.B2(n_4519),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4625),
.Y(n_4691)
);

AOI221xp5_ASAP7_75t_L g4692 ( 
.A1(n_4661),
.A2(n_4576),
.B1(n_4541),
.B2(n_4578),
.C(n_4575),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4599),
.A2(n_4462),
.B(n_4449),
.Y(n_4693)
);

AOI211xp5_ASAP7_75t_L g4694 ( 
.A1(n_4647),
.A2(n_4473),
.B(n_4506),
.C(n_4497),
.Y(n_4694)
);

AOI22xp33_ASAP7_75t_L g4695 ( 
.A1(n_4590),
.A2(n_4460),
.B1(n_716),
.B2(n_711),
.Y(n_4695)
);

O2A1O1Ixp5_ASAP7_75t_SL g4696 ( 
.A1(n_4587),
.A2(n_716),
.B(n_711),
.C(n_713),
.Y(n_4696)
);

NOR2x1_ASAP7_75t_SL g4697 ( 
.A(n_4619),
.B(n_717),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4601),
.Y(n_4698)
);

AOI211xp5_ASAP7_75t_SL g4699 ( 
.A1(n_4606),
.A2(n_723),
.B(n_719),
.C(n_721),
.Y(n_4699)
);

NOR2x1_ASAP7_75t_L g4700 ( 
.A(n_4591),
.B(n_721),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4588),
.B(n_961),
.Y(n_4701)
);

AOI21xp33_ASAP7_75t_L g4702 ( 
.A1(n_4667),
.A2(n_723),
.B(n_724),
.Y(n_4702)
);

AOI221xp5_ASAP7_75t_L g4703 ( 
.A1(n_4598),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.C(n_728),
.Y(n_4703)
);

O2A1O1Ixp5_ASAP7_75t_L g4704 ( 
.A1(n_4664),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_4704)
);

NOR4xp25_ASAP7_75t_SL g4705 ( 
.A(n_4643),
.B(n_731),
.C(n_728),
.D(n_730),
.Y(n_4705)
);

AOI22xp33_ASAP7_75t_SL g4706 ( 
.A1(n_4658),
.A2(n_733),
.B1(n_730),
.B2(n_732),
.Y(n_4706)
);

NOR2x1_ASAP7_75t_L g4707 ( 
.A(n_4605),
.B(n_732),
.Y(n_4707)
);

INVx3_ASAP7_75t_L g4708 ( 
.A(n_4648),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4639),
.B(n_4593),
.Y(n_4709)
);

OAI322xp33_ASAP7_75t_L g4710 ( 
.A1(n_4654),
.A2(n_733),
.A3(n_734),
.B1(n_735),
.B2(n_736),
.C1(n_737),
.C2(n_738),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4650),
.Y(n_4711)
);

OA21x2_ASAP7_75t_L g4712 ( 
.A1(n_4586),
.A2(n_734),
.B(n_735),
.Y(n_4712)
);

OR2x2_ASAP7_75t_L g4713 ( 
.A(n_4660),
.B(n_737),
.Y(n_4713)
);

AOI21xp33_ASAP7_75t_L g4714 ( 
.A1(n_4641),
.A2(n_739),
.B(n_740),
.Y(n_4714)
);

OAI21xp5_ASAP7_75t_L g4715 ( 
.A1(n_4637),
.A2(n_739),
.B(n_740),
.Y(n_4715)
);

NAND3xp33_ASAP7_75t_L g4716 ( 
.A(n_4629),
.B(n_741),
.C(n_742),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4616),
.Y(n_4717)
);

OAI21xp5_ASAP7_75t_L g4718 ( 
.A1(n_4612),
.A2(n_743),
.B(n_744),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4621),
.Y(n_4719)
);

O2A1O1Ixp33_ASAP7_75t_L g4720 ( 
.A1(n_4663),
.A2(n_4607),
.B(n_4638),
.C(n_4642),
.Y(n_4720)
);

INVx2_ASAP7_75t_L g4721 ( 
.A(n_4609),
.Y(n_4721)
);

OAI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4613),
.A2(n_748),
.B1(n_743),
.B2(n_747),
.Y(n_4722)
);

INVx1_ASAP7_75t_SL g4723 ( 
.A(n_4662),
.Y(n_4723)
);

AOI22xp5_ASAP7_75t_L g4724 ( 
.A1(n_4640),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.Y(n_4724)
);

AOI22xp5_ASAP7_75t_L g4725 ( 
.A1(n_4624),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_4725)
);

AOI221xp5_ASAP7_75t_L g4726 ( 
.A1(n_4657),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.C(n_755),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4681),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4712),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4699),
.A2(n_4631),
.B1(n_4653),
.B2(n_4659),
.Y(n_4729)
);

OAI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4669),
.A2(n_4608),
.B1(n_4636),
.B2(n_4618),
.Y(n_4730)
);

HB1xp67_ASAP7_75t_L g4731 ( 
.A(n_4712),
.Y(n_4731)
);

O2A1O1Ixp33_ASAP7_75t_SL g4732 ( 
.A1(n_4676),
.A2(n_4594),
.B(n_4633),
.C(n_4646),
.Y(n_4732)
);

AOI211xp5_ASAP7_75t_L g4733 ( 
.A1(n_4714),
.A2(n_4644),
.B(n_4595),
.C(n_4645),
.Y(n_4733)
);

OAI211xp5_ASAP7_75t_L g4734 ( 
.A1(n_4670),
.A2(n_4627),
.B(n_4652),
.C(n_4630),
.Y(n_4734)
);

OAI221xp5_ASAP7_75t_SL g4735 ( 
.A1(n_4674),
.A2(n_4603),
.B1(n_4656),
.B2(n_4651),
.C(n_4634),
.Y(n_4735)
);

XOR2x2_ASAP7_75t_L g4736 ( 
.A(n_4671),
.B(n_4649),
.Y(n_4736)
);

O2A1O1Ixp33_ASAP7_75t_L g4737 ( 
.A1(n_4704),
.A2(n_4666),
.B(n_4665),
.C(n_4668),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4701),
.Y(n_4738)
);

OAI21xp33_ASAP7_75t_SL g4739 ( 
.A1(n_4684),
.A2(n_753),
.B(n_754),
.Y(n_4739)
);

OAI21xp5_ASAP7_75t_SL g4740 ( 
.A1(n_4683),
.A2(n_756),
.B(n_757),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4697),
.Y(n_4741)
);

AOI221xp5_ASAP7_75t_L g4742 ( 
.A1(n_4690),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.C(n_759),
.Y(n_4742)
);

OAI21xp5_ASAP7_75t_L g4743 ( 
.A1(n_4672),
.A2(n_758),
.B(n_759),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4708),
.B(n_760),
.Y(n_4744)
);

OAI211xp5_ASAP7_75t_L g4745 ( 
.A1(n_4715),
.A2(n_763),
.B(n_761),
.C(n_762),
.Y(n_4745)
);

AO22x2_ASAP7_75t_L g4746 ( 
.A1(n_4673),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.Y(n_4746)
);

OR3x1_ASAP7_75t_L g4747 ( 
.A(n_4680),
.B(n_766),
.C(n_767),
.Y(n_4747)
);

OAI211xp5_ASAP7_75t_SL g4748 ( 
.A1(n_4723),
.A2(n_4675),
.B(n_4689),
.C(n_4709),
.Y(n_4748)
);

AOI22xp5_ASAP7_75t_L g4749 ( 
.A1(n_4685),
.A2(n_770),
.B1(n_767),
.B2(n_769),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4708),
.Y(n_4750)
);

OA22x2_ASAP7_75t_L g4751 ( 
.A1(n_4677),
.A2(n_773),
.B1(n_769),
.B2(n_770),
.Y(n_4751)
);

AOI22xp5_ASAP7_75t_L g4752 ( 
.A1(n_4692),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_4752)
);

AOI221xp5_ASAP7_75t_L g4753 ( 
.A1(n_4702),
.A2(n_777),
.B1(n_774),
.B2(n_776),
.C(n_778),
.Y(n_4753)
);

OAI221xp5_ASAP7_75t_L g4754 ( 
.A1(n_4695),
.A2(n_4686),
.B1(n_4679),
.B2(n_4694),
.C(n_4718),
.Y(n_4754)
);

CKINVDCx16_ASAP7_75t_R g4755 ( 
.A(n_4705),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4713),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4700),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4706),
.B(n_777),
.Y(n_4758)
);

XNOR2x1_ASAP7_75t_L g4759 ( 
.A(n_4682),
.B(n_779),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4688),
.Y(n_4760)
);

AOI21xp33_ASAP7_75t_L g4761 ( 
.A1(n_4720),
.A2(n_781),
.B(n_782),
.Y(n_4761)
);

A2O1A1Ixp33_ASAP7_75t_SL g4762 ( 
.A1(n_4727),
.A2(n_4698),
.B(n_4721),
.C(n_4719),
.Y(n_4762)
);

AOI221xp5_ASAP7_75t_L g4763 ( 
.A1(n_4732),
.A2(n_4740),
.B1(n_4729),
.B2(n_4761),
.C(n_4754),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4728),
.Y(n_4764)
);

INVxp67_ASAP7_75t_L g4765 ( 
.A(n_4731),
.Y(n_4765)
);

AND2x4_ASAP7_75t_L g4766 ( 
.A(n_4741),
.B(n_4691),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4751),
.Y(n_4767)
);

AOI22xp5_ASAP7_75t_L g4768 ( 
.A1(n_4747),
.A2(n_4707),
.B1(n_4716),
.B2(n_4722),
.Y(n_4768)
);

AOI22xp5_ASAP7_75t_L g4769 ( 
.A1(n_4748),
.A2(n_4703),
.B1(n_4711),
.B2(n_4726),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4759),
.Y(n_4770)
);

NOR2xp33_ASAP7_75t_L g4771 ( 
.A(n_4755),
.B(n_4725),
.Y(n_4771)
);

NOR2x1_ASAP7_75t_L g4772 ( 
.A(n_4757),
.B(n_4710),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4746),
.Y(n_4773)
);

O2A1O1Ixp33_ASAP7_75t_L g4774 ( 
.A1(n_4750),
.A2(n_4717),
.B(n_4687),
.C(n_4678),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4746),
.Y(n_4775)
);

NOR2xp67_ASAP7_75t_L g4776 ( 
.A(n_4739),
.B(n_4724),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4744),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4758),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4736),
.Y(n_4779)
);

XNOR2x1_ASAP7_75t_L g4780 ( 
.A(n_4772),
.B(n_4770),
.Y(n_4780)
);

NAND4xp75_ASAP7_75t_L g4781 ( 
.A(n_4763),
.B(n_4743),
.C(n_4760),
.D(n_4738),
.Y(n_4781)
);

OAI22xp5_ASAP7_75t_L g4782 ( 
.A1(n_4769),
.A2(n_4752),
.B1(n_4735),
.B2(n_4733),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4773),
.Y(n_4783)
);

NAND4xp75_ASAP7_75t_L g4784 ( 
.A(n_4771),
.B(n_4742),
.C(n_4753),
.D(n_4756),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4775),
.Y(n_4785)
);

INVx2_ASAP7_75t_SL g4786 ( 
.A(n_4766),
.Y(n_4786)
);

NOR2xp67_ASAP7_75t_L g4787 ( 
.A(n_4765),
.B(n_4745),
.Y(n_4787)
);

AND2x4_ASAP7_75t_L g4788 ( 
.A(n_4767),
.B(n_4693),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4764),
.Y(n_4789)
);

NAND3xp33_ASAP7_75t_L g4790 ( 
.A(n_4774),
.B(n_4730),
.C(n_4734),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4768),
.Y(n_4791)
);

OAI221xp5_ASAP7_75t_L g4792 ( 
.A1(n_4786),
.A2(n_4762),
.B1(n_4737),
.B2(n_4779),
.C(n_4776),
.Y(n_4792)
);

NOR2xp33_ASAP7_75t_SL g4793 ( 
.A(n_4787),
.B(n_4778),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4780),
.A2(n_4777),
.B(n_4749),
.Y(n_4794)
);

OAI21xp33_ASAP7_75t_SL g4795 ( 
.A1(n_4781),
.A2(n_4696),
.B(n_781),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4783),
.B(n_783),
.Y(n_4796)
);

AOI22xp5_ASAP7_75t_L g4797 ( 
.A1(n_4788),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_4797)
);

A2O1A1Ixp33_ASAP7_75t_L g4798 ( 
.A1(n_4790),
.A2(n_4785),
.B(n_4789),
.C(n_4791),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4784),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4782),
.Y(n_4800)
);

OA22x2_ASAP7_75t_L g4801 ( 
.A1(n_4797),
.A2(n_789),
.B1(n_787),
.B2(n_788),
.Y(n_4801)
);

INVx2_ASAP7_75t_SL g4802 ( 
.A(n_4796),
.Y(n_4802)
);

XNOR2xp5_ASAP7_75t_L g4803 ( 
.A(n_4792),
.B(n_787),
.Y(n_4803)
);

NAND3x1_ASAP7_75t_L g4804 ( 
.A(n_4794),
.B(n_788),
.C(n_789),
.Y(n_4804)
);

BUFx2_ASAP7_75t_L g4805 ( 
.A(n_4804),
.Y(n_4805)
);

NAND4xp75_ASAP7_75t_L g4806 ( 
.A(n_4802),
.B(n_4799),
.C(n_4800),
.D(n_4795),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4801),
.Y(n_4807)
);

OAI31xp33_ASAP7_75t_L g4808 ( 
.A1(n_4805),
.A2(n_4798),
.A3(n_4803),
.B(n_4793),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4808),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4809),
.Y(n_4810)
);

AO21x2_ASAP7_75t_L g4811 ( 
.A1(n_4810),
.A2(n_4807),
.B(n_4806),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4811),
.B(n_790),
.Y(n_4812)
);

AOI21xp5_ASAP7_75t_L g4813 ( 
.A1(n_4812),
.A2(n_790),
.B(n_791),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4813),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4813),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.Y(n_4815)
);

NAND3xp33_ASAP7_75t_L g4816 ( 
.A(n_4814),
.B(n_795),
.C(n_797),
.Y(n_4816)
);

NAND2x2_ASAP7_75t_L g4817 ( 
.A(n_4815),
.B(n_797),
.Y(n_4817)
);

AOI22xp5_ASAP7_75t_L g4818 ( 
.A1(n_4816),
.A2(n_804),
.B1(n_800),
.B2(n_803),
.Y(n_4818)
);

AOI211xp5_ASAP7_75t_L g4819 ( 
.A1(n_4818),
.A2(n_4817),
.B(n_804),
.C(n_800),
.Y(n_4819)
);


endmodule