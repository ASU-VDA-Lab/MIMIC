module real_jpeg_15796_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_617, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_617;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_611;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_120;
wire n_155;
wire n_572;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_614),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_0),
.B(n_615),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_1),
.A2(n_57),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_1),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_1),
.A2(n_365),
.B1(n_396),
.B2(n_399),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_1),
.A2(n_365),
.B1(n_536),
.B2(n_539),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_1),
.A2(n_365),
.B1(n_547),
.B2(n_549),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_101),
.B1(n_110),
.B2(n_121),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_110),
.B1(n_239),
.B2(n_244),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_2),
.A2(n_110),
.B1(n_349),
.B2(n_353),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_3),
.A2(n_357),
.B1(n_358),
.B2(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_3),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_3),
.A2(n_357),
.B1(n_421),
.B2(n_424),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_3),
.A2(n_357),
.B1(n_513),
.B2(n_518),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_3),
.A2(n_354),
.B1(n_357),
.B2(n_569),
.Y(n_568)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_4),
.Y(n_227)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_4),
.Y(n_384)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_6),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_6),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_6),
.A2(n_297),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_6),
.A2(n_297),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_6),
.A2(n_297),
.B1(n_523),
.B2(n_525),
.Y(n_522)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_7),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_8),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_8),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_8),
.A2(n_255),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_8),
.A2(n_255),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_8),
.A2(n_255),
.B1(n_483),
.B2(n_488),
.Y(n_482)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_9),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_9),
.B(n_62),
.Y(n_434)
);

OAI32xp33_ASAP7_75t_L g474 ( 
.A1(n_9),
.A2(n_70),
.A3(n_404),
.B1(n_475),
.B2(n_478),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_9),
.B(n_94),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_9),
.A2(n_221),
.B1(n_381),
.B2(n_568),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_9),
.A2(n_331),
.B1(n_587),
.B2(n_588),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_65),
.B1(n_97),
.B2(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_65),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_65),
.B1(n_229),
.B2(n_234),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

BUFx4f_ASAP7_75t_L g352 ( 
.A(n_11),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_50),
.B1(n_56),
.B2(n_60),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_60),
.B1(n_119),
.B2(n_124),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_60),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_12),
.A2(n_60),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_13),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_14),
.A2(n_136),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_14),
.A2(n_136),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g342 ( 
.A1(n_14),
.A2(n_136),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_16),
.A2(n_108),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_16),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_16),
.A2(n_183),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_16),
.A2(n_183),
.B1(n_375),
.B2(n_377),
.Y(n_374)
);

OAI22x1_ASAP7_75t_SL g426 ( 
.A1(n_16),
.A2(n_183),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_17),
.Y(n_156)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_17),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_17),
.Y(n_379)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_17),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g359 ( 
.A(n_19),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_19),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_170),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_168),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_66),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_49),
.B1(n_61),
.B2(n_63),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_25),
.A2(n_49),
.B1(n_61),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_25),
.A2(n_61),
.B1(n_131),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_25),
.A2(n_37),
.B1(n_180),
.B2(n_253),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g293 ( 
.A1(n_25),
.A2(n_37),
.B1(n_253),
.B2(n_294),
.Y(n_293)
);

OAI22x1_ASAP7_75t_SL g386 ( 
.A1(n_25),
.A2(n_61),
.B1(n_294),
.B2(n_364),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_26),
.A2(n_62),
.B1(n_107),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_26),
.A2(n_62),
.B1(n_356),
.B2(n_363),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_26),
.A2(n_62),
.B1(n_356),
.B2(n_401),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_34),
.B(n_37),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_34),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_35),
.Y(n_333)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22x1_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_43),
.Y(n_127)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_45),
.Y(n_215)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_56),
.B(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g296 ( 
.A(n_59),
.Y(n_296)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_66),
.B(n_173),
.Y(n_613)
);

FAx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_105),
.CI(n_115),
.CON(n_66),
.SN(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_94),
.B(n_95),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_68),
.A2(n_94),
.B1(n_210),
.B2(n_216),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_68),
.A2(n_94),
.B1(n_316),
.B2(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_68),
.A2(n_94),
.B1(n_395),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_96),
.B1(n_118),
.B2(n_128),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_69),
.A2(n_118),
.B1(n_128),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_69),
.A2(n_128),
.B1(n_211),
.B2(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_69),
.A2(n_128),
.B1(n_315),
.B2(n_321),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_69),
.A2(n_128),
.B1(n_301),
.B2(n_321),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_69),
.A2(n_128),
.B1(n_420),
.B2(n_586),
.Y(n_585)
);

AO21x2_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_87),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_76),
.Y(n_317)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_78),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_86),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_88),
.Y(n_376)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_92),
.Y(n_208)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_92),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_93),
.Y(n_406)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_104),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_104),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_129),
.C(n_137),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_117),
.B1(n_137),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_121),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_122),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_123),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_126),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_126),
.Y(n_399)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_127),
.Y(n_398)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_127),
.Y(n_592)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_137),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_178),
.C(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_137),
.B(n_186),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_151),
.B(n_163),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_138),
.A2(n_151),
.B1(n_163),
.B2(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_138),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_138),
.A2(n_151),
.B1(n_403),
.B2(n_411),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_138),
.A2(n_151),
.B1(n_510),
.B2(n_512),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_138),
.A2(n_151),
.B1(n_512),
.B2(n_535),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_138),
.A2(n_151),
.B1(n_465),
.B2(n_535),
.Y(n_594)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_139),
.A2(n_203),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_139),
.A2(n_237),
.B1(n_270),
.B2(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_139),
.A2(n_237),
.B1(n_464),
.B2(n_471),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_139),
.B(n_331),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_146),
.B2(n_149),
.Y(n_140)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_145),
.Y(n_284)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_145),
.Y(n_354)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_145),
.Y(n_428)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_145),
.Y(n_487)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_148),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_148),
.Y(n_548)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_148),
.Y(n_565)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_150),
.Y(n_504)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_151),
.B(n_269),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_160),
.B2(n_162),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_156),
.Y(n_470)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_160),
.Y(n_498)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_167),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21x1_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_188),
.B(n_612),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_184),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_177),
.B1(n_178),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_308),
.B(n_609),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_258),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_192),
.A2(n_610),
.B(n_611),
.Y(n_609)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_193),
.B(n_196),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_217),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_200),
.A2(n_201),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_204),
.Y(n_511)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_206),
.Y(n_466)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_217),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_249),
.B1(n_257),
.B2(n_617),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_218),
.A2(n_219),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_251),
.B1(n_252),
.B2(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_220),
.A2(n_236),
.B1(n_257),
.B2(n_446),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_226),
.B(n_228),
.Y(n_220)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_221),
.A2(n_341),
.B1(n_346),
.B2(n_348),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_221),
.A2(n_281),
.B1(n_348),
.B2(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_221),
.A2(n_290),
.B1(n_522),
.B2(n_530),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_221),
.A2(n_546),
.B1(n_568),
.B2(n_572),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_224),
.Y(n_347)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_225),
.Y(n_497)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_227),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_231),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_232),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_236),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_243),
.Y(n_410)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_254),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_305),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_259),
.B(n_305),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_261),
.B(n_265),
.Y(n_440)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_266),
.B(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_292),
.C(n_300),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_267),
.B(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_276),
.B(n_278),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_268),
.B(n_276),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_278),
.B(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_289),
.B2(n_291),
.Y(n_278)
);

AOI22x1_ASAP7_75t_SL g425 ( 
.A1(n_279),
.A2(n_342),
.B1(n_426),
.B2(n_432),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_279),
.A2(n_382),
.B1(n_426),
.B2(n_482),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_279),
.A2(n_545),
.B1(n_552),
.B2(n_553),
.Y(n_544)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_293),
.B(n_300),
.Y(n_444)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_455),
.B(n_604),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_438),
.C(n_450),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_388),
.B(n_412),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_311),
.B(n_388),
.C(n_606),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_368),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_312),
.B(n_369),
.C(n_371),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_328),
.C(n_355),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_314),
.B(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_340),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_340),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_338),
.B2(n_339),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_SL g401 ( 
.A1(n_330),
.A2(n_331),
.B(n_358),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_331),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_331),
.B(n_500),
.Y(n_499)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_331),
.A2(n_499),
.B(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_331),
.B(n_433),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_351),
.Y(n_488)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_352),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_352),
.Y(n_524)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_385),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_380),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_374),
.Y(n_411)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_378),
.Y(n_540)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_381),
.Y(n_552)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_386),
.B(n_387),
.C(n_449),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_393),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_390),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_392),
.B(n_393),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_400),
.C(n_402),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_402),
.Y(n_415)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_415),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_435),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_413),
.B(n_435),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.C(n_417),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_417),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.C(n_434),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx2_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_434),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_436),
.Y(n_437)
);

A2O1A1O1Ixp25_ASAP7_75t_L g604 ( 
.A1(n_438),
.A2(n_450),
.B(n_605),
.C(n_607),
.D(n_608),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_441),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_439),
.B(n_441),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.C(n_447),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_442),
.A2(n_443),
.B1(n_445),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_445),
.Y(n_453)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_451),
.B(n_454),
.Y(n_607)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_489),
.B(n_603),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_457),
.B(n_459),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.C(n_472),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_460),
.A2(n_461),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_463),
.A2(n_472),
.B1(n_473),
.B2(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_480),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_474),
.A2(n_480),
.B1(n_481),
.B2(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_474),
.Y(n_582)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_479),
.Y(n_500)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_596),
.B(n_602),
.Y(n_489)
);

AOI21x1_ASAP7_75t_SL g490 ( 
.A1(n_491),
.A2(n_578),
.B(n_595),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_542),
.B(n_577),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_520),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_493),
.B(n_520),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_508),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_494),
.A2(n_508),
.B1(n_509),
.B2(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

OAI32xp33_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_497),
.A3(n_498),
.B1(n_499),
.B2(n_501),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_517),
.Y(n_538)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_531),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_521),
.B(n_533),
.C(n_541),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_522),
.Y(n_553)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_533),
.B1(n_534),
.B2(n_541),
.Y(n_531)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_532),
.Y(n_541)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_543),
.A2(n_556),
.B(n_576),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_554),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_544),
.B(n_554),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_557),
.A2(n_570),
.B(n_575),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_567),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_566),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_574),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_574),
.Y(n_575)
);

INVx6_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_580),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_579),
.B(n_580),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_583),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_581),
.B(n_584),
.C(n_594),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_584),
.A2(n_585),
.B1(n_593),
.B2(n_594),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_SL g596 ( 
.A(n_597),
.B(n_601),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_597),
.B(n_601),
.Y(n_602)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);


endmodule