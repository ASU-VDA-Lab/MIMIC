module real_jpeg_13056_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_0),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_0),
.A2(n_44),
.B1(n_46),
.B2(n_61),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_43),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_84),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_6),
.A2(n_44),
.B1(n_46),
.B2(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_84),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_7),
.A2(n_44),
.B1(n_46),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_7),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_7),
.B(n_34),
.C(n_49),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_82),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_117),
.B(n_170),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_64),
.B(n_81),
.C(n_197),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_7),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_7),
.B(n_58),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_44),
.B1(n_46),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_166),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_166),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_166),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_9),
.A2(n_44),
.B1(n_46),
.B2(n_126),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_126),
.Y(n_245)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_44),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_12),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_12),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_15),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_329)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_16),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_20),
.B(n_340),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_18),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_18),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_18),
.A2(n_44),
.B1(n_46),
.B2(n_73),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_73),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_18),
.A2(n_64),
.B1(n_65),
.B2(n_73),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_335),
.B(n_338),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_327),
.B(n_331),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_314),
.B(n_326),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_142),
.B(n_311),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_129),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_104),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_26),
.B(n_104),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_74),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_27),
.B(n_75),
.C(n_90),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_56),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_28),
.A2(n_29),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_30),
.A2(n_31),
.B1(n_56),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_30),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_32),
.A2(n_36),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_32),
.B(n_171),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_32),
.A2(n_36),
.B1(n_116),
.B2(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_33),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_36),
.B(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_38),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_55),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_42),
.A2(n_47),
.B1(n_55),
.B2(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_46),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_44),
.B(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_46),
.A2(n_80),
.B(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_55),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_47),
.B(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_47),
.A2(n_55),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_47),
.A2(n_55),
.B1(n_121),
.B2(n_248),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_53),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_51),
.A2(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_51),
.B(n_154),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_51),
.A2(n_167),
.B(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_55),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B(n_67),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_62),
.B1(n_69),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_59),
.A2(n_69),
.B(n_154),
.C(n_241),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_59),
.A2(n_64),
.A3(n_66),
.B1(n_242),
.B2(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_72),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_69),
.B1(n_93),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_62),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_62),
.A2(n_67),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_62),
.A2(n_69),
.B1(n_125),
.B2(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_63),
.B(n_65),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_68),
.A2(n_222),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_68),
.A2(n_222),
.B1(n_321),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_68),
.A2(n_222),
.B(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_90),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_76),
.B(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_83),
.B1(n_85),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_77),
.A2(n_85),
.B1(n_98),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_77),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_77),
.A2(n_85),
.B1(n_217),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_77),
.A2(n_203),
.B(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_82),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_78),
.B(n_204),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_78),
.A2(n_82),
.B(n_318),
.Y(n_317)
);

NOR2x1_ASAP7_75t_R g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_82),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_85),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_85),
.A2(n_123),
.B(n_218),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_88),
.A2(n_155),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_103),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_92),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_95),
.C(n_100),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_92),
.B(n_133),
.C(n_140),
.Y(n_325)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_100),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_100),
.B(n_134),
.C(n_138),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_111),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_110),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_111),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.C(n_124),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_112),
.A2(n_113),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_114),
.A2(n_119),
.B1(n_120),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_114),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_117),
.A2(n_118),
.B1(n_199),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_117),
.A2(n_118),
.B1(n_225),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_118),
.A2(n_176),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_118),
.B(n_154),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_118),
.A2(n_184),
.B(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_122),
.B(n_124),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_128),
.B(n_240),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_129),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_130),
.B(n_141),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_135),
.Y(n_320)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_139),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_305),
.B(n_310),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_293),
.B(n_304),
.Y(n_143)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_261),
.A3(n_286),
.B1(n_291),
.B2(n_292),
.C(n_343),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_234),
.B(n_260),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_211),
.B(n_233),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_192),
.B(n_210),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_172),
.B(n_191),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_150),
.B(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_169),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_180),
.B(n_190),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_178),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_205),
.C(n_209),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_198),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_226),
.B2(n_227),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_229),
.C(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_220),
.C(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_236),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_250),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_251),
.C(n_252),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_243),
.B2(n_249),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_244),
.C(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_272),
.C(n_275),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_264),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_270),
.C(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_280),
.C(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_283),
.C(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_303),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_336),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule