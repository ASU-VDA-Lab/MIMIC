module real_jpeg_7008_n_21 (n_17, n_8, n_0, n_93, n_2, n_10, n_9, n_12, n_92, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_94, n_1, n_20, n_19, n_16, n_15, n_13, n_21);

input n_17;
input n_8;
input n_0;
input n_93;
input n_2;
input n_10;
input n_9;
input n_12;
input n_92;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_94;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

INVx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_18),
.B(n_81),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_18),
.C(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_6),
.A2(n_20),
.B(n_33),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_20),
.C(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_9),
.A2(n_13),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_11),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_16),
.C(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_11),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_29),
.B(n_92),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.C(n_94),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_15),
.B(n_27),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_15),
.C(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_26),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_32),
.A2(n_39),
.B(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_61),
.C(n_62),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI311xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_83),
.A3(n_85),
.B1(n_86),
.C1(n_87),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.C(n_42),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_80),
.B(n_82),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_75),
.B(n_79),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B(n_73),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_65),
.B(n_69),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_64),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_59),
.B(n_63),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_56),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_77),
.C(n_78),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_93),
.Y(n_55)
);


endmodule