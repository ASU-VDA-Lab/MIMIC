module fake_jpeg_7444_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.C(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_2),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_41),
.B1(n_51),
.B2(n_33),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_25),
.B1(n_17),
.B2(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_37),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_43),
.C(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_68),
.B1(n_38),
.B2(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_77),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_29),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_59),
.B1(n_69),
.B2(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_54),
.B1(n_52),
.B2(n_67),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_81),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_66),
.B(n_34),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_39),
.B1(n_49),
.B2(n_15),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_39),
.B(n_34),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_87),
.B(n_80),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_102),
.C(n_88),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_70),
.C(n_83),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_82),
.B(n_74),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_92),
.B(n_95),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_72),
.B(n_39),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_80),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_102),
.C(n_99),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_95),
.B1(n_84),
.B2(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_107),
.B1(n_29),
.B2(n_5),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_115),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_92),
.B(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_104),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_108),
.C(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_115),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_119),
.C(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_4),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_6),
.C1(n_3),
.C2(n_4),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_116),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_129),
.B1(n_5),
.B2(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.Y(n_133)
);


endmodule