module real_jpeg_12483_n_17 (n_5, n_4, n_8, n_0, n_12, n_327, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_327;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_84),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_4),
.A2(n_60),
.B1(n_65),
.B2(n_84),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_84),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_113),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_60),
.B1(n_65),
.B2(n_113),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_113),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_8),
.A2(n_52),
.B1(n_60),
.B2(n_65),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_76),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_9),
.A2(n_60),
.B1(n_65),
.B2(n_76),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_10),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_10),
.A2(n_60),
.B1(n_65),
.B2(n_179),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_179),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_179),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_12),
.A2(n_44),
.B1(n_60),
.B2(n_65),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_13),
.B(n_60),
.C(n_64),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_31),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_138),
.B(n_183),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_27),
.B(n_30),
.C(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_167),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_13),
.B(n_53),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_13),
.B(n_40),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_14),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_14),
.A2(n_60),
.B1(n_65),
.B2(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_147),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_15),
.A2(n_36),
.B1(n_60),
.B2(n_65),
.Y(n_103)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_77),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_37),
.B1(n_54),
.B2(n_55),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_24),
.A2(n_31),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_24),
.B(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_26),
.A2(n_32),
.B(n_167),
.Y(n_210)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_28),
.B(n_48),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g266 ( 
.A1(n_30),
.A2(n_41),
.A3(n_49),
.B1(n_254),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_31),
.B(n_217),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_33),
.B(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_46),
.B1(n_47),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_41),
.A2(n_46),
.B(n_167),
.C(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_45),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_47),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_46),
.A2(n_47),
.B1(n_146),
.B2(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_83),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_47),
.B(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_47),
.A2(n_110),
.B(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_70),
.C(n_74),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_70),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_81),
.B1(n_86),
.B2(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_66),
.B(n_68),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_66),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_66),
.B1(n_106),
.B2(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_58),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_58),
.A2(n_66),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_58),
.A2(n_66),
.B1(n_142),
.B2(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_69),
.B1(n_108),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_59),
.A2(n_178),
.B(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_59),
.B(n_167),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_59),
.A2(n_180),
.B(n_259),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_65),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_66),
.B(n_169),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_73),
.B1(n_88),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_71),
.A2(n_73),
.B1(n_117),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_71),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_71),
.A2(n_73),
.B1(n_230),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_71),
.A2(n_216),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_73),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_73),
.A2(n_144),
.B(n_231),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_85),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_78),
.A2(n_82),
.B1(n_121),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_85),
.B(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_155),
.B(n_323),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_150),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_125),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_94),
.B(n_125),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_114),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_115),
.C(n_120),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B(n_109),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_97),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_109),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_100),
.A2(n_101),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_100),
.B(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_100),
.A2(n_101),
.B1(n_137),
.B2(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_101),
.B(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_116),
.B(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_119),
.A2(n_168),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_131),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_132),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.C(n_145),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_133),
.A2(n_134),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_135),
.A2(n_140),
.B1(n_141),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_135),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_138),
.A2(n_139),
.B1(n_212),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_138),
.A2(n_139),
.B1(n_237),
.B2(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_139),
.A2(n_189),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_167),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_139),
.A2(n_197),
.B(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_143),
.B(n_145),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_149),
.B(n_252),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_150),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_151),
.B(n_154),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_317),
.B(n_322),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_305),
.B(n_316),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_273),
.A3(n_298),
.B1(n_303),
.B2(n_304),
.C(n_327),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_246),
.B(n_272),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_224),
.B(n_245),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_205),
.B(n_223),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_185),
.B(n_204),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_165),
.B1(n_170),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_181),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_177),
.C(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_193),
.B(n_203),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_191),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_198),
.B(n_202),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_218),
.C(n_222),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_211),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_238),
.B2(n_239),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_241),
.C(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_248),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_262),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_263),
.C(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_255),
.B2(n_261),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_256),
.C(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_288),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.C(n_287),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_276),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_282),
.C(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_292),
.C(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_315),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_315),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);


endmodule