module fake_netlist_6_4347_n_1955 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1955);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1955;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_154),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_113),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_100),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_33),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_88),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_38),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_96),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_168),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_97),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_71),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g237 ( 
.A(n_201),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_133),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_65),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_56),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_31),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_59),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_145),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_161),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_115),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_194),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_34),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_9),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_25),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_172),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_67),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_8),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_186),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_108),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_103),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_22),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_149),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_1),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_76),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_191),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_175),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_98),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_187),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_176),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_73),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_35),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_20),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_70),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_132),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_122),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_102),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_20),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_146),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_183),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_66),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_141),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_94),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_36),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_137),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_174),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_89),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_163),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_80),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_84),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_19),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_48),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_17),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_33),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_124),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_184),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_162),
.Y(n_319)
);

BUFx2_ASAP7_75t_SL g320 ( 
.A(n_104),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_189),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_56),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_30),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_148),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_12),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_67),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_111),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_155),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_24),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_5),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_81),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_197),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_202),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_126),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_140),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_45),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_43),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_48),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_193),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_170),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_22),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_29),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_129),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_169),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_91),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_8),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_76),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_72),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_55),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_116),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_95),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_62),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_65),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_109),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_125),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_178),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_158),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_93),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_166),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_44),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_30),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_17),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_61),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_117),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_110),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_64),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_153),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_135),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_54),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_150),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_3),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_44),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_14),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_60),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_105),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_123),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_182),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_112),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_177),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_57),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_54),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_165),
.Y(n_384)
);

BUFx2_ASAP7_75t_SL g385 ( 
.A(n_45),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_121),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_171),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_152),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_92),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_50),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_29),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_139),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_36),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_118),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_21),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_143),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_205),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_190),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_142),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_79),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_62),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_40),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_7),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_138),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_185),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_344),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_287),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_258),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_287),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_287),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_211),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_287),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_206),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_366),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_207),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_366),
.B(n_1),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_208),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_346),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_229),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_286),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_210),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_292),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_291),
.B(n_305),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_213),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_218),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_219),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_214),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_289),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_223),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_226),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_228),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_230),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_368),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_401),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_231),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_235),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_238),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_372),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_240),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_373),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_289),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_389),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_250),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_252),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_255),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_209),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_371),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_378),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_358),
.B(n_4),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_215),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_241),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_227),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_400),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_358),
.B(n_9),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_291),
.B(n_11),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_217),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_305),
.B(n_11),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_214),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_267),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_332),
.B(n_12),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_301),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_334),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_386),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_269),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_271),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_209),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_224),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_365),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_273),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_214),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_358),
.B(n_13),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_237),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_274),
.Y(n_490)
);

BUFx6f_ASAP7_75t_SL g491 ( 
.A(n_216),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_224),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_234),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_234),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_259),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_212),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_279),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_332),
.B(n_14),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_280),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_236),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_222),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_281),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_236),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_389),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_233),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_259),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_268),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_285),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_242),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_212),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

AND3x2_ASAP7_75t_L g512 ( 
.A(n_418),
.B(n_248),
.C(n_221),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_424),
.A2(n_312),
.B1(n_314),
.B2(n_323),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_415),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_268),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_442),
.B(n_242),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_413),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_412),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_466),
.B(n_221),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_417),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_457),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_466),
.B(n_248),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_419),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_426),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

NAND2x1_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_379),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_425),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_429),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_489),
.B(n_298),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_421),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_430),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_434),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_421),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_436),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_437),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_444),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_458),
.B(n_243),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_445),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_496),
.B(n_220),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_438),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_446),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_457),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_448),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_504),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_416),
.A2(n_370),
.B1(n_313),
.B2(n_257),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_504),
.B(n_243),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_447),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_504),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_439),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_439),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_510),
.B(n_220),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_450),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_510),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_463),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_483),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_464),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_433),
.B(n_302),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_478),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_443),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_427),
.A2(n_403),
.B1(n_247),
.B2(n_395),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_582),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_521),
.A2(n_502),
.B1(n_406),
.B2(n_467),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_543),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_583),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_517),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_451),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_453),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_577),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_530),
.B(n_469),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_534),
.B(n_455),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_534),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_530),
.B(n_469),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_546),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_385),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_546),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

BUFx4f_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

INVxp33_ASAP7_75t_SL g622 ( 
.A(n_585),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_593),
.B(n_385),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_527),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_574),
.B(n_468),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_571),
.B(n_471),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_577),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_525),
.Y(n_629)
);

AO22x2_ASAP7_75t_L g630 ( 
.A1(n_569),
.A2(n_498),
.B1(n_477),
.B2(n_247),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_540),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_565),
.B(n_459),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_379),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_521),
.A2(n_480),
.B1(n_479),
.B2(n_461),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_545),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_460),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_519),
.B(n_476),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_563),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_586),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_532),
.B(n_481),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_525),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_522),
.B(n_495),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_567),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_587),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_522),
.B(n_482),
.Y(n_646)
);

INVx4_ASAP7_75t_SL g647 ( 
.A(n_535),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_535),
.B(n_261),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_524),
.B(n_320),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_520),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_586),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_511),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_535),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_590),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_526),
.A2(n_486),
.B1(n_497),
.B2(n_490),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_525),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_561),
.B(n_472),
.Y(n_657)
);

INVx4_ASAP7_75t_SL g658 ( 
.A(n_525),
.Y(n_658)
);

BUFx4f_ASAP7_75t_L g659 ( 
.A(n_525),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_536),
.B(n_499),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_520),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_525),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_520),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_533),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_525),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_533),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_541),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_526),
.A2(n_508),
.B1(n_485),
.B2(n_449),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_511),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_514),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_590),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_427),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_569),
.B(n_474),
.C(n_475),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_524),
.B(n_488),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_549),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_514),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_557),
.B(n_488),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_515),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_554),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_585),
.A2(n_449),
.B1(n_367),
.B2(n_263),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_537),
.B(n_487),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_531),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_554),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_553),
.B(n_491),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_561),
.B(n_261),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_531),
.A2(n_491),
.B1(n_470),
.B2(n_465),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_557),
.B(n_452),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_515),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_561),
.B(n_578),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_516),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_539),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_539),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_554),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_537),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_516),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_550),
.B(n_381),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_554),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_518),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_556),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_578),
.B(n_307),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_SL g703 ( 
.A(n_578),
.B(n_491),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_554),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_518),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_551),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_551),
.Y(n_708)
);

BUFx8_ASAP7_75t_SL g709 ( 
.A(n_560),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_512),
.A2(n_300),
.B1(n_245),
.B2(n_403),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_523),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_554),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_528),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_528),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_512),
.B(n_328),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_564),
.B(n_573),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_529),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_579),
.B(n_506),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_554),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_303),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_551),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_558),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_538),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_550),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_542),
.B(n_408),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_581),
.B(n_379),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_580),
.A2(n_325),
.B1(n_245),
.B2(n_249),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_581),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_513),
.B(n_246),
.C(n_239),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_581),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_225),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_550),
.B(n_381),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_513),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_544),
.B(n_308),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_544),
.B(n_260),
.C(n_256),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_548),
.Y(n_736)
);

AND2x2_ASAP7_75t_SL g737 ( 
.A(n_580),
.B(n_225),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_548),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_552),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_552),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_691),
.A2(n_317),
.B1(n_405),
.B2(n_398),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_625),
.B(n_484),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_691),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_691),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_653),
.B(n_555),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_660),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_602),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_660),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_689),
.B(n_550),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_602),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_596),
.B(n_232),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_653),
.B(n_555),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_657),
.A2(n_340),
.B1(n_277),
.B2(n_360),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_678),
.B(n_559),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_678),
.B(n_559),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_612),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_599),
.B(n_264),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_678),
.B(n_562),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_594),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_620),
.B(n_379),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_612),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_595),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_600),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_596),
.B(n_232),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_675),
.B(n_244),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_620),
.A2(n_340),
.B1(n_244),
.B2(n_251),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_601),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_641),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_626),
.B(n_562),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_674),
.B(n_266),
.C(n_265),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_620),
.B(n_379),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_689),
.B(n_588),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_657),
.B(n_588),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_605),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_627),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_649),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_603),
.B(n_576),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_604),
.B(n_576),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_687),
.B(n_387),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_694),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_651),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_709),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_566),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_706),
.B(n_581),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_706),
.B(n_581),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_740),
.B(n_581),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_641),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_736),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_709),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_643),
.B(n_588),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_740),
.B(n_592),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_738),
.B(n_646),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_687),
.A2(n_648),
.B1(n_737),
.B2(n_630),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_652),
.B(n_592),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_647),
.B(n_387),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_670),
.B(n_592),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_608),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_671),
.B(n_592),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_677),
.B(n_592),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_618),
.B(n_275),
.C(n_270),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_647),
.B(n_387),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_647),
.B(n_702),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_622),
.B(n_276),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_614),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_616),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_679),
.B(n_581),
.Y(n_810)
);

NOR2x1p5_ASAP7_75t_L g811 ( 
.A(n_599),
.B(n_278),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_682),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_690),
.B(n_591),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_692),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_650),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_697),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_737),
.B(n_387),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_700),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_684),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_650),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_705),
.B(n_592),
.Y(n_821)
);

AO221x1_ASAP7_75t_L g822 ( 
.A1(n_630),
.A2(n_681),
.B1(n_251),
.B2(n_284),
.C(n_277),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_711),
.B(n_592),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_713),
.B(n_591),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_714),
.B(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_591),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_649),
.A2(n_345),
.B1(n_309),
.B2(n_404),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_622),
.B(n_282),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_728),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_649),
.A2(n_339),
.B1(n_310),
.B2(n_399),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_695),
.A2(n_693),
.B(n_659),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_723),
.B(n_591),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_609),
.A2(n_570),
.B(n_558),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_591),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_616),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_662),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_636),
.B(n_253),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_687),
.B(n_253),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_662),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_637),
.B(n_640),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_649),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_720),
.B(n_284),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_696),
.B(n_484),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_630),
.B(n_492),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_661),
.B(n_283),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_L g846 ( 
.A(n_687),
.B(n_293),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_664),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_664),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_734),
.B(n_293),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_731),
.B(n_262),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_665),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_687),
.A2(n_331),
.B1(n_297),
.B2(n_306),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_687),
.A2(n_331),
.B1(n_297),
.B2(n_306),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_665),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_718),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_668),
.B(n_216),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_631),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_731),
.B(n_333),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_667),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_607),
.B(n_492),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_607),
.B(n_290),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_724),
.B(n_311),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_613),
.B(n_295),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_724),
.B(n_318),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_613),
.B(n_493),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_683),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_648),
.B(n_317),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_648),
.B(n_321),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_648),
.B(n_321),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_707),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_708),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_654),
.B(n_493),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_721),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_611),
.B(n_324),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_606),
.Y(n_876)
);

OAI22xp33_ASAP7_75t_L g877 ( 
.A1(n_615),
.A2(n_360),
.B1(n_327),
.B2(n_343),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_615),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_655),
.B(n_296),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_611),
.B(n_324),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_698),
.B(n_732),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_722),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_611),
.B(n_617),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_633),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_597),
.B(n_319),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_617),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_617),
.B(n_327),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_621),
.B(n_343),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_606),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_715),
.B(n_335),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_615),
.A2(n_405),
.B1(n_398),
.B2(n_347),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_621),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_794),
.B(n_676),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_774),
.A2(n_703),
.B1(n_716),
.B2(n_732),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_840),
.B(n_673),
.C(n_634),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_845),
.B(n_733),
.C(n_729),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_778),
.B(n_686),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_774),
.A2(n_703),
.B1(n_698),
.B2(n_733),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_861),
.A2(n_725),
.B(n_735),
.C(n_710),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_831),
.A2(n_659),
.B(n_633),
.Y(n_902)
);

O2A1O1Ixp5_ASAP7_75t_L g903 ( 
.A1(n_760),
.A2(n_621),
.B(n_598),
.C(n_619),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_779),
.B(n_623),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_834),
.A2(n_619),
.B(n_598),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_792),
.B(n_623),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_819),
.B(n_668),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_792),
.B(n_623),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_773),
.B(n_623),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_780),
.A2(n_619),
.B(n_598),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_802),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_749),
.B(n_676),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_799),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_883),
.A2(n_642),
.B(n_629),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_817),
.A2(n_663),
.B(n_642),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_744),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_892),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_873),
.B(n_676),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_863),
.A2(n_388),
.B(n_347),
.C(n_384),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_817),
.A2(n_767),
.B(n_877),
.C(n_753),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_881),
.A2(n_701),
.B1(n_688),
.B2(n_669),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_802),
.Y(n_922)
);

NAND2x1_ASAP7_75t_L g923 ( 
.A(n_876),
.B(n_889),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_837),
.B(n_663),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_802),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_795),
.A2(n_701),
.B1(n_727),
.B2(n_392),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_855),
.B(n_624),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_873),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_760),
.A2(n_680),
.B(n_666),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_812),
.B(n_635),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_807),
.B(n_828),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_747),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_772),
.A2(n_680),
.B(n_666),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_881),
.A2(n_680),
.B1(n_685),
.B2(n_628),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_879),
.A2(n_685),
.B(n_336),
.C(n_326),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_802),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_881),
.A2(n_865),
.B(n_860),
.C(n_755),
.Y(n_937)
);

NOR2x1p5_ASAP7_75t_SL g938 ( 
.A(n_893),
.B(n_558),
.Y(n_938)
);

AOI22x1_ASAP7_75t_L g939 ( 
.A1(n_884),
.A2(n_685),
.B1(n_730),
.B2(n_712),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_843),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_747),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_890),
.A2(n_726),
.B(n_364),
.C(n_294),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_856),
.A2(n_315),
.B(n_299),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_843),
.B(n_635),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_802),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_754),
.A2(n_712),
.B(n_704),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_782),
.B(n_606),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_782),
.B(n_606),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_742),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_750),
.Y(n_950)
);

AOI22x1_ASAP7_75t_SL g951 ( 
.A1(n_784),
.A2(n_631),
.B1(n_645),
.B2(n_644),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_SL g952 ( 
.A(n_878),
.B(n_672),
.Y(n_952)
);

OAI321xp33_ASAP7_75t_L g953 ( 
.A1(n_891),
.A2(n_395),
.A3(n_249),
.B1(n_254),
.B2(n_336),
.C(n_326),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_799),
.Y(n_954)
);

CKINVDCx10_ASAP7_75t_R g955 ( 
.A(n_784),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_758),
.A2(n_699),
.B(n_704),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_860),
.A2(n_304),
.B(n_288),
.C(n_254),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_801),
.B(n_638),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_770),
.A2(n_699),
.B(n_712),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_782),
.B(n_656),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_865),
.B(n_656),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_786),
.A2(n_719),
.B(n_656),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_787),
.A2(n_719),
.B(n_575),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_788),
.A2(n_570),
.B(n_572),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_842),
.A2(n_288),
.B(n_300),
.C(n_304),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_759),
.B(n_658),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_793),
.A2(n_570),
.B(n_572),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_742),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_809),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_746),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_809),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_885),
.B(n_638),
.C(n_645),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_771),
.A2(n_375),
.B(n_330),
.Y(n_973)
);

OAI321xp33_ASAP7_75t_L g974 ( 
.A1(n_885),
.A2(n_391),
.A3(n_382),
.B1(n_272),
.B2(n_390),
.C(n_349),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_804),
.B(n_644),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_762),
.B(n_658),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_749),
.B(n_352),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_748),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_766),
.B(n_494),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_763),
.B(n_658),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_878),
.B(n_672),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_741),
.A2(n_320),
.B1(n_369),
.B2(n_377),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_750),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_790),
.B(n_259),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_772),
.A2(n_575),
.B(n_355),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_849),
.A2(n_376),
.B(n_272),
.C(n_349),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_857),
.B(n_494),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_766),
.B(n_500),
.Y(n_988)
);

BUFx4f_ASAP7_75t_L g989 ( 
.A(n_777),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_785),
.A2(n_380),
.B(n_356),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_890),
.A2(n_382),
.B(n_322),
.C(n_325),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_768),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_844),
.B(n_500),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_829),
.A2(n_397),
.B(n_359),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_835),
.B(n_316),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_844),
.A2(n_376),
.B(n_322),
.C(n_390),
.Y(n_996)
);

BUFx4f_ASAP7_75t_L g997 ( 
.A(n_777),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_751),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_775),
.B(n_337),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_838),
.A2(n_394),
.B(n_396),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_777),
.B(n_841),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_765),
.A2(n_391),
.B(n_357),
.C(n_341),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_765),
.A2(n_374),
.B(n_338),
.C(n_342),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_751),
.Y(n_1004)
);

AND2x2_ASAP7_75t_SL g1005 ( 
.A(n_846),
.B(n_503),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_776),
.B(n_348),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_781),
.B(n_783),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_814),
.B(n_350),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_756),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_816),
.B(n_354),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_796),
.A2(n_509),
.B(n_462),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_818),
.B(n_393),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_745),
.A2(n_462),
.B(n_456),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_751),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_761),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_752),
.A2(n_454),
.B(n_402),
.Y(n_1016)
);

OAI321xp33_ASAP7_75t_L g1017 ( 
.A1(n_827),
.A2(n_216),
.A3(n_383),
.B1(n_363),
.B2(n_362),
.C(n_23),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_757),
.B(n_15),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_808),
.B(n_862),
.Y(n_1019)
);

AO32x1_ASAP7_75t_L g1020 ( 
.A1(n_822),
.A2(n_15),
.A3(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_806),
.A2(n_198),
.B(n_173),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_833),
.A2(n_167),
.B(n_157),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_797),
.A2(n_136),
.B(n_134),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_808),
.B(n_16),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_862),
.B(n_864),
.C(n_857),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_797),
.A2(n_131),
.B(n_130),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_798),
.A2(n_127),
.B(n_120),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_809),
.B(n_101),
.Y(n_1028)
);

AOI222xp33_ASAP7_75t_L g1029 ( 
.A1(n_822),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.C1(n_26),
.C2(n_27),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_761),
.A2(n_90),
.B(n_87),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_764),
.B(n_26),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_764),
.B(n_28),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_864),
.B(n_830),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_769),
.A2(n_86),
.B(n_85),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_809),
.A2(n_82),
.B1(n_78),
.B2(n_32),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_769),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_789),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_800),
.A2(n_37),
.B(n_41),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_803),
.A2(n_37),
.B(n_41),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_809),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_789),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_810),
.A2(n_42),
.B(n_46),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_777),
.A2(n_75),
.B1(n_49),
.B2(n_50),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_764),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_841),
.A2(n_75),
.B1(n_53),
.B2(n_55),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_791),
.B(n_52),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_813),
.A2(n_57),
.B(n_58),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_791),
.B(n_58),
.C(n_61),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_821),
.A2(n_63),
.B(n_64),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_823),
.A2(n_63),
.B(n_66),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_841),
.B(n_867),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_875),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_868),
.A2(n_74),
.B(n_69),
.C(n_70),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_815),
.B(n_68),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_824),
.A2(n_68),
.B(n_69),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_852),
.B(n_72),
.C(n_74),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_815),
.B(n_854),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_820),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_853),
.A2(n_886),
.B1(n_869),
.B2(n_893),
.Y(n_1059)
);

OAI321xp33_ASAP7_75t_L g1060 ( 
.A1(n_880),
.A2(n_887),
.A3(n_888),
.B1(n_858),
.B2(n_850),
.C(n_825),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_826),
.A2(n_832),
.B(n_805),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_886),
.B(n_876),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_820),
.A2(n_874),
.B(n_836),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_876),
.B(n_889),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_811),
.B(n_839),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_848),
.A2(n_871),
.B(n_882),
.C(n_851),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_931),
.B(n_839),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_928),
.B(n_847),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_963),
.A2(n_962),
.B(n_1063),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_937),
.B(n_859),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_899),
.B(n_866),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_940),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_927),
.B(n_870),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_918),
.B(n_872),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_1033),
.A2(n_920),
.B(n_897),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_911),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_901),
.A2(n_1019),
.B(n_904),
.C(n_909),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_961),
.B(n_906),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_908),
.B(n_993),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1001),
.B(n_979),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_913),
.Y(n_1081)
);

AOI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_974),
.A2(n_1017),
.B(n_1029),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_992),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_895),
.B(n_1007),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_947),
.A2(n_948),
.B(n_960),
.Y(n_1085)
);

AOI21xp33_ASAP7_75t_L g1086 ( 
.A1(n_926),
.A2(n_991),
.B(n_1031),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1052),
.B(n_949),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_946),
.A2(n_959),
.B(n_956),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_979),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_903),
.A2(n_985),
.B(n_1051),
.C(n_919),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_977),
.A2(n_894),
.B(n_935),
.C(n_1034),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1060),
.A2(n_1059),
.B(n_915),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_968),
.B(n_944),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_954),
.B(n_975),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_934),
.A2(n_946),
.B(n_959),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_930),
.B(n_958),
.Y(n_1096)
);

AOI221x1_ASAP7_75t_L g1097 ( 
.A1(n_896),
.A2(n_1025),
.B1(n_1042),
.B2(n_1050),
.C(n_1039),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_907),
.B(n_900),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_921),
.B(n_981),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_924),
.A2(n_1054),
.B(n_1024),
.C(n_933),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_898),
.B(n_916),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_929),
.A2(n_1064),
.B(n_1057),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_917),
.B(n_999),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_987),
.B(n_988),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_911),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1062),
.A2(n_1005),
.B(n_980),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_957),
.A2(n_1002),
.A3(n_1053),
.B(n_1049),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_966),
.A2(n_976),
.B(n_1004),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_932),
.B(n_941),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_1018),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_998),
.A2(n_925),
.B(n_936),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_950),
.B(n_983),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1066),
.A2(n_964),
.B(n_967),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1014),
.B(n_989),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1009),
.B(n_1015),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1037),
.B(n_1058),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_969),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1036),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_923),
.A2(n_1041),
.B(n_925),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_936),
.B(n_1065),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_988),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_1032),
.A2(n_953),
.B(n_996),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_989),
.A2(n_997),
.B(n_1028),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_952),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_969),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_971),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1023),
.A2(n_1026),
.B(n_990),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_997),
.A2(n_971),
.B(n_922),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1006),
.B(n_1010),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1021),
.A2(n_1027),
.B(n_1011),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_912),
.A2(n_994),
.B(n_978),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_1013),
.B(n_942),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_971),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_970),
.B(n_922),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_945),
.A2(n_1012),
.B(n_1000),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_972),
.B(n_984),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_943),
.B(n_973),
.C(n_1046),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1016),
.A2(n_1008),
.B(n_995),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1035),
.A2(n_982),
.B(n_1056),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_938),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_965),
.Y(n_1141)
);

CKINVDCx12_ASAP7_75t_R g1142 ( 
.A(n_955),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_951),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1038),
.A2(n_1055),
.A3(n_1050),
.B(n_1049),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1038),
.A2(n_1055),
.B(n_1047),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1003),
.B(n_986),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1044),
.B(n_1043),
.C(n_1045),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1040),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1048),
.B(n_1020),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1020),
.A2(n_937),
.B(n_902),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1001),
.B(n_766),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_931),
.B(n_937),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_931),
.B(n_855),
.Y(n_1154)
);

AOI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_931),
.A2(n_1033),
.B(n_753),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_931),
.B(n_937),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_992),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_SL g1159 ( 
.A1(n_931),
.A2(n_840),
.B(n_879),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_907),
.B(n_635),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_911),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_931),
.B(n_937),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_937),
.A2(n_902),
.B(n_774),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_940),
.Y(n_1166)
);

BUFx4f_ASAP7_75t_L g1167 ( 
.A(n_1001),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_932),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_969),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_931),
.B(n_937),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_940),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_931),
.B(n_937),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_931),
.B(n_918),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_913),
.Y(n_1176)
);

AO22x1_ASAP7_75t_L g1177 ( 
.A1(n_931),
.A2(n_840),
.B1(n_896),
.B2(n_733),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_931),
.A2(n_840),
.B1(n_1033),
.B2(n_896),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_914),
.A2(n_939),
.B(n_963),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_902),
.A2(n_937),
.A3(n_935),
.B(n_919),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_R g1181 ( 
.A(n_940),
.B(n_784),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_SL g1182 ( 
.A1(n_1021),
.A2(n_1022),
.B(n_1030),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_L g1183 ( 
.A(n_901),
.B(n_937),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_910),
.A2(n_620),
.B(n_653),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_937),
.A2(n_902),
.B(n_774),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1001),
.B(n_766),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_932),
.Y(n_1187)
);

AOI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_931),
.A2(n_1033),
.B(n_753),
.Y(n_1188)
);

AOI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_931),
.A2(n_1033),
.B(n_753),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_992),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_940),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_902),
.A2(n_937),
.A3(n_935),
.B(n_919),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_931),
.B(n_937),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_931),
.A2(n_1033),
.B(n_920),
.C(n_901),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_L g1195 ( 
.A1(n_902),
.A2(n_905),
.B(n_1061),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_931),
.A2(n_1033),
.B(n_920),
.C(n_901),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1160),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_1159),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1155),
.A2(n_1189),
.B1(n_1188),
.B2(n_1156),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1099),
.A2(n_1075),
.B1(n_1149),
.B2(n_1154),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_1104),
.Y(n_1202)
);

AND2x6_ASAP7_75t_L g1203 ( 
.A(n_1149),
.B(n_1153),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1125),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1079),
.B(n_1071),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1177),
.B(n_1073),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1083),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1184),
.A2(n_1183),
.B(n_1182),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1158),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1190),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1079),
.B(n_1071),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_1167),
.B(n_1149),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1075),
.B(n_1138),
.C(n_1097),
.Y(n_1214)
);

INVx3_ASAP7_75t_SL g1215 ( 
.A(n_1110),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1142),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1165),
.A2(n_1185),
.B(n_1151),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1096),
.B(n_1175),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1167),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1103),
.B(n_1093),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1136),
.A2(n_1098),
.B(n_1191),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1093),
.B(n_1166),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1172),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1093),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1080),
.B(n_1089),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1087),
.B(n_1121),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1087),
.B(n_1074),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1125),
.Y(n_1228)
);

INVx5_ASAP7_75t_L g1229 ( 
.A(n_1125),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1143),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1164),
.A2(n_1171),
.B(n_1193),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1081),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1124),
.B(n_1080),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1168),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1089),
.B(n_1176),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1181),
.Y(n_1236)
);

OR2x6_ASAP7_75t_SL g1237 ( 
.A(n_1147),
.B(n_1173),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1152),
.B(n_1186),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1126),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1173),
.B(n_1193),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1067),
.B(n_1078),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1067),
.B(n_1078),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1094),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1077),
.A2(n_1092),
.B(n_1100),
.Y(n_1244)
);

BUFx4f_ASAP7_75t_SL g1245 ( 
.A(n_1143),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1152),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1126),
.Y(n_1247)
);

AOI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1148),
.A2(n_1084),
.B(n_1086),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1120),
.B(n_1186),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1163),
.B(n_1117),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1114),
.B(n_1120),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1082),
.B(n_1163),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1187),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1084),
.A2(n_1101),
.B1(n_1070),
.B2(n_1150),
.Y(n_1254)
);

CKINVDCx8_ASAP7_75t_R g1255 ( 
.A(n_1143),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1133),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1117),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1169),
.B(n_1076),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1086),
.A2(n_1122),
.B1(n_1137),
.B2(n_1139),
.C(n_1150),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1091),
.B(n_1146),
.C(n_1141),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1134),
.Y(n_1262)
);

NAND2x1_ASAP7_75t_L g1263 ( 
.A(n_1076),
.B(n_1105),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1118),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1134),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1133),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1122),
.A2(n_1070),
.B1(n_1140),
.B2(n_1115),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1109),
.A2(n_1116),
.B1(n_1115),
.B2(n_1112),
.Y(n_1268)
);

OR2x2_ASAP7_75t_SL g1269 ( 
.A(n_1133),
.B(n_1116),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1112),
.B(n_1131),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1095),
.A2(n_1135),
.B(n_1102),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1106),
.B(n_1085),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1163),
.B(n_1105),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1163),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1119),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1123),
.B(n_1128),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1111),
.B(n_1195),
.Y(n_1277)
);

AOI221xp5_ASAP7_75t_L g1278 ( 
.A1(n_1090),
.A2(n_1113),
.B1(n_1108),
.B2(n_1107),
.C(n_1144),
.Y(n_1278)
);

INVx3_ASAP7_75t_SL g1279 ( 
.A(n_1107),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_SL g1280 ( 
.A(n_1180),
.B(n_1192),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_SL g1281 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_1180),
.C(n_1192),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1107),
.A2(n_1180),
.B(n_1192),
.C(n_1144),
.Y(n_1282)
);

OR2x2_ASAP7_75t_SL g1283 ( 
.A(n_1127),
.B(n_1130),
.Y(n_1283)
);

AO32x1_ASAP7_75t_L g1284 ( 
.A1(n_1157),
.A2(n_1161),
.A3(n_1179),
.B1(n_1174),
.B2(n_1170),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1069),
.B(n_1088),
.Y(n_1285)
);

OR2x6_ASAP7_75t_L g1286 ( 
.A(n_1132),
.B(n_1162),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1080),
.B(n_1089),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1154),
.B(n_928),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1129),
.A2(n_931),
.B1(n_1188),
.B2(n_1155),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1083),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1081),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_1194),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_1194),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1083),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1083),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1297)
);

AND2x6_ASAP7_75t_L g1298 ( 
.A(n_1149),
.B(n_1153),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1083),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1167),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1081),
.Y(n_1301)
);

AND2x6_ASAP7_75t_L g1302 ( 
.A(n_1149),
.B(n_1153),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1129),
.B(n_1178),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1160),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1072),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_1194),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1154),
.B(n_928),
.Y(n_1308)
);

OAI31xp33_ASAP7_75t_L g1309 ( 
.A1(n_1129),
.A2(n_1159),
.A3(n_931),
.B(n_1155),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1167),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1081),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1072),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1083),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1093),
.B(n_1001),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_931),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1178),
.B(n_928),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1129),
.A2(n_1159),
.B(n_1188),
.C(n_1155),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1093),
.B(n_1001),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1159),
.B(n_931),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1072),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1159),
.A2(n_1129),
.B(n_931),
.C(n_1155),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1129),
.A2(n_931),
.B1(n_1188),
.B2(n_1155),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1129),
.A2(n_931),
.B1(n_1188),
.B2(n_1155),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1103),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1080),
.B(n_1089),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_1194),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1129),
.A2(n_931),
.B1(n_1159),
.B2(n_1178),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1081),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1129),
.A2(n_840),
.B(n_931),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1178),
.B(n_1194),
.Y(n_1331)
);

NOR2x1_ASAP7_75t_SL g1332 ( 
.A(n_1163),
.B(n_1001),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1129),
.A2(n_931),
.B1(n_1188),
.B2(n_1155),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1165),
.A2(n_1185),
.B(n_1151),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1072),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1159),
.B(n_931),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1083),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1129),
.B2(n_1194),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1207),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1228),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1303),
.A2(n_1289),
.B1(n_1333),
.B2(n_1324),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1237),
.B(n_1199),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1320),
.A2(n_1336),
.B1(n_1338),
.B2(n_1307),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1211),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1203),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1290),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1198),
.B(n_1293),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1219),
.B(n_1300),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1295),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1232),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1197),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1228),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1335),
.Y(n_1354)
);

CKINVDCx11_ASAP7_75t_R g1355 ( 
.A(n_1255),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1296),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1210),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1313),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1323),
.A2(n_1309),
.B1(n_1292),
.B2(n_1327),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1291),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1330),
.A2(n_1328),
.B1(n_1201),
.B2(n_1206),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1199),
.B(n_1318),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1321),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1198),
.B(n_1293),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1335),
.Y(n_1366)
);

CKINVDCx6p67_ASAP7_75t_R g1367 ( 
.A(n_1215),
.Y(n_1367)
);

BUFx2_ASAP7_75t_R g1368 ( 
.A(n_1304),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1337),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1276),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1276),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1297),
.B(n_1306),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1264),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1230),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1316),
.A2(n_1338),
.B1(n_1307),
.B2(n_1292),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1234),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1309),
.A2(n_1294),
.B1(n_1327),
.B2(n_1331),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1305),
.Y(n_1378)
);

BUFx2_ASAP7_75t_R g1379 ( 
.A(n_1266),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1294),
.A2(n_1252),
.B1(n_1213),
.B2(n_1200),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1301),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1329),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1297),
.A2(n_1306),
.B1(n_1331),
.B2(n_1315),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1253),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1218),
.A2(n_1302),
.B1(n_1298),
.B2(n_1203),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1219),
.B(n_1300),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1317),
.A2(n_1322),
.B1(n_1269),
.B2(n_1221),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1203),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1312),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1315),
.A2(n_1203),
.B1(n_1302),
.B2(n_1298),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1252),
.A2(n_1200),
.B1(n_1298),
.B2(n_1302),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1298),
.A2(n_1302),
.B1(n_1214),
.B2(n_1261),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1202),
.A2(n_1308),
.B1(n_1288),
.B2(n_1220),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1214),
.A2(n_1334),
.B1(n_1217),
.B2(n_1325),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1262),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1228),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1314),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1223),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_R g1399 ( 
.A1(n_1226),
.A2(n_1311),
.B1(n_1224),
.B2(n_1245),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_SL g1400 ( 
.A(n_1287),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1205),
.A2(n_1212),
.B1(n_1241),
.B2(n_1242),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1260),
.A2(n_1240),
.B1(n_1231),
.B2(n_1334),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1208),
.B(n_1314),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1265),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1217),
.A2(n_1325),
.B1(n_1227),
.B2(n_1310),
.Y(n_1405)
);

BUFx2_ASAP7_75t_R g1406 ( 
.A(n_1236),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1222),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1310),
.A2(n_1233),
.B1(n_1231),
.B2(n_1244),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1265),
.Y(n_1409)
);

BUFx2_ASAP7_75t_R g1410 ( 
.A(n_1246),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1229),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1216),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1251),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_R g1414 ( 
.A(n_1229),
.B(n_1258),
.Y(n_1414)
);

BUFx8_ASAP7_75t_SL g1415 ( 
.A(n_1225),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1275),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1238),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1249),
.B(n_1251),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1229),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1238),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1235),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1287),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1256),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1254),
.A2(n_1278),
.B(n_1272),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1267),
.A2(n_1243),
.B1(n_1238),
.B2(n_1314),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1225),
.Y(n_1426)
);

AO21x1_ASAP7_75t_L g1427 ( 
.A1(n_1244),
.A2(n_1248),
.B(n_1254),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1279),
.B(n_1225),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1326),
.B(n_1248),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1263),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1268),
.A2(n_1270),
.B(n_1271),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1280),
.B(n_1319),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1319),
.A2(n_1280),
.B1(n_1277),
.B2(n_1285),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1274),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1259),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1204),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1282),
.B(n_1332),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1285),
.A2(n_1259),
.B1(n_1258),
.B2(n_1247),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1204),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1204),
.A2(n_1239),
.B1(n_1247),
.B2(n_1257),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1273),
.A2(n_1250),
.B1(n_1283),
.B2(n_1239),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1239),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1250),
.A2(n_1273),
.B1(n_1257),
.B2(n_1247),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_R g1444 ( 
.A1(n_1281),
.A2(n_1257),
.B1(n_1284),
.B2(n_1286),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1286),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1284),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1237),
.B(n_1199),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1232),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1207),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1210),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1203),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_931),
.B2(n_1155),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1330),
.A2(n_1159),
.B1(n_1129),
.B2(n_1178),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1207),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_931),
.B2(n_1155),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1255),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1228),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_1159),
.B2(n_931),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1210),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1228),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1207),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1207),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1219),
.B(n_1300),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_931),
.B2(n_1155),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_931),
.B2(n_1155),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1276),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1210),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1216),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1207),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1203),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1228),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1232),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1230),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1303),
.A2(n_1129),
.B1(n_931),
.B2(n_1155),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1335),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1328),
.A2(n_1159),
.B1(n_1178),
.B2(n_1129),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_1232),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1276),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1403),
.B(n_1424),
.Y(n_1479)
);

BUFx4f_ASAP7_75t_SL g1480 ( 
.A(n_1374),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1427),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1427),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1346),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1366),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1452),
.B(n_1455),
.Y(n_1488)
);

CKINVDCx6p67_ASAP7_75t_R g1489 ( 
.A(n_1355),
.Y(n_1489)
);

BUFx4f_ASAP7_75t_SL g1490 ( 
.A(n_1374),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1364),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1447),
.B(n_1432),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1403),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1404),
.Y(n_1495)
);

BUFx4f_ASAP7_75t_SL g1496 ( 
.A(n_1412),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1446),
.A2(n_1431),
.B(n_1402),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1447),
.B(n_1365),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1431),
.A2(n_1392),
.B(n_1377),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1444),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1429),
.B(n_1348),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1416),
.A2(n_1371),
.B(n_1370),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1409),
.Y(n_1503)
);

AO21x1_ASAP7_75t_L g1504 ( 
.A1(n_1375),
.A2(n_1476),
.B(n_1453),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1362),
.A2(n_1387),
.B(n_1441),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1437),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1437),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1401),
.B(n_1424),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1365),
.B(n_1394),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1416),
.A2(n_1478),
.B(n_1466),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1355),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1344),
.A2(n_1464),
.B1(n_1474),
.B2(n_1465),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1450),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1459),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1420),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1360),
.B(n_1418),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1348),
.B(n_1372),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1357),
.Y(n_1518)
);

INVxp33_ASAP7_75t_L g1519 ( 
.A(n_1378),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1418),
.B(n_1380),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1359),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1433),
.A2(n_1390),
.B(n_1383),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1467),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1388),
.B(n_1451),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1413),
.B(n_1372),
.Y(n_1526)
);

AO21x1_ASAP7_75t_SL g1527 ( 
.A1(n_1385),
.A2(n_1342),
.B(n_1458),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1369),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1373),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1445),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1445),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1425),
.A2(n_1339),
.B(n_1340),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1371),
.B(n_1466),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1478),
.B(n_1428),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1393),
.B(n_1451),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1420),
.Y(n_1536)
);

CKINVDCx6p67_ASAP7_75t_R g1537 ( 
.A(n_1456),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1470),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1470),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1345),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1407),
.B(n_1354),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1420),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1347),
.A2(n_1454),
.B(n_1449),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1350),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1356),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1386),
.B(n_1463),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1358),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1461),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1420),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1408),
.B(n_1405),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1462),
.Y(n_1551)
);

BUFx4f_ASAP7_75t_SL g1552 ( 
.A(n_1412),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1469),
.A2(n_1430),
.B(n_1376),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1384),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1434),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1349),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1349),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1414),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1396),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1396),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1475),
.B(n_1398),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1389),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1426),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1386),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1435),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1426),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_SL g1568 ( 
.A(n_1479),
.B(n_1457),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1506),
.B(n_1417),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1518),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1553),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1521),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1523),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1521),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1498),
.B(n_1463),
.Y(n_1576)
);

NOR2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1505),
.B(n_1367),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1509),
.B(n_1438),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1487),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1543),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1506),
.B(n_1417),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1479),
.B(n_1471),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1481),
.B(n_1491),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1501),
.B(n_1422),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1493),
.B(n_1443),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1504),
.A2(n_1399),
.B1(n_1400),
.B2(n_1473),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1508),
.A2(n_1460),
.B(n_1353),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1483),
.B(n_1423),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1507),
.B(n_1423),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1502),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1525),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1483),
.B(n_1410),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1507),
.B(n_1367),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1486),
.B(n_1442),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1481),
.B(n_1460),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1526),
.B(n_1442),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1502),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1525),
.Y(n_1600)
);

OAI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1512),
.A2(n_1440),
.B(n_1473),
.C(n_1472),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1481),
.B(n_1491),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1496),
.B(n_1552),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1510),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1513),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1514),
.B(n_1351),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1517),
.B(n_1477),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1488),
.A2(n_1471),
.B1(n_1468),
.B2(n_1411),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1495),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1534),
.B(n_1352),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1479),
.B(n_1471),
.Y(n_1612)
);

OAI33xp33_ASAP7_75t_L g1613 ( 
.A1(n_1556),
.A2(n_1406),
.A3(n_1415),
.B1(n_1379),
.B2(n_1352),
.B3(n_1368),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1503),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1485),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1534),
.B(n_1352),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1563),
.B(n_1472),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1555),
.B(n_1351),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1491),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1482),
.B(n_1341),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1588),
.A2(n_1504),
.B1(n_1508),
.B2(n_1550),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1588),
.A2(n_1527),
.B1(n_1499),
.B2(n_1550),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1572),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1613),
.B(n_1480),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1505),
.C(n_1559),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1570),
.B(n_1492),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1609),
.B(n_1549),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1589),
.B(n_1549),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1594),
.A2(n_1520),
.B(n_1500),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1603),
.A2(n_1484),
.B1(n_1500),
.B2(n_1519),
.C(n_1555),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1484),
.C(n_1499),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1573),
.B(n_1556),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1606),
.A2(n_1531),
.B1(n_1530),
.B2(n_1566),
.C(n_1520),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1499),
.C(n_1535),
.Y(n_1634)
);

NAND4xp25_ASAP7_75t_L g1635 ( 
.A(n_1575),
.B(n_1531),
.C(n_1535),
.D(n_1548),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1580),
.B(n_1499),
.C(n_1559),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1594),
.A2(n_1524),
.B(n_1516),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1532),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1572),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1578),
.A2(n_1527),
.B1(n_1522),
.B2(n_1516),
.Y(n_1640)
);

AND2x2_ASAP7_75t_SL g1641 ( 
.A(n_1593),
.B(n_1494),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1532),
.Y(n_1642)
);

AND2x2_ASAP7_75t_SL g1643 ( 
.A(n_1593),
.B(n_1539),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1586),
.B(n_1532),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1585),
.B(n_1479),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1585),
.B(n_1497),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1604),
.A2(n_1524),
.B(n_1567),
.Y(n_1647)
);

AOI211xp5_ASAP7_75t_L g1648 ( 
.A1(n_1595),
.A2(n_1557),
.B(n_1558),
.C(n_1567),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1595),
.A2(n_1537),
.B1(n_1489),
.B2(n_1564),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1577),
.A2(n_1522),
.B(n_1542),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1576),
.B(n_1528),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1602),
.B(n_1497),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1578),
.A2(n_1522),
.B1(n_1489),
.B2(n_1537),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1598),
.B(n_1529),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1620),
.B(n_1497),
.C(n_1558),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1620),
.B(n_1557),
.C(n_1561),
.Y(n_1656)
);

OAI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1607),
.A2(n_1564),
.B1(n_1515),
.B2(n_1536),
.C(n_1549),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1587),
.A2(n_1565),
.B(n_1554),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1568),
.A2(n_1522),
.B1(n_1587),
.B2(n_1600),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1611),
.B(n_1490),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1569),
.A2(n_1583),
.B1(n_1618),
.B2(n_1577),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1617),
.A2(n_1551),
.B1(n_1545),
.B2(n_1547),
.C(n_1548),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1591),
.B(n_1540),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1584),
.A2(n_1539),
.B1(n_1533),
.B2(n_1565),
.C(n_1547),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1596),
.B(n_1546),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1611),
.A2(n_1549),
.B(n_1546),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_L g1668 ( 
.A(n_1579),
.B(n_1561),
.C(n_1560),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1590),
.B(n_1616),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1584),
.A2(n_1515),
.B1(n_1536),
.B2(n_1381),
.C(n_1382),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1584),
.A2(n_1612),
.B1(n_1361),
.B2(n_1381),
.C(n_1382),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1590),
.B(n_1540),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1623),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1639),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1646),
.B(n_1600),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1644),
.B(n_1579),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1638),
.B(n_1574),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1664),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1662),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1642),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1668),
.Y(n_1682)
);

INVx5_ASAP7_75t_L g1683 ( 
.A(n_1645),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1629),
.B(n_1596),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1631),
.B(n_1579),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1632),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1634),
.B(n_1581),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1655),
.B(n_1636),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1672),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1643),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1648),
.B(n_1602),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1656),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1641),
.Y(n_1693)
);

AND2x4_ASAP7_75t_SL g1694 ( 
.A(n_1640),
.B(n_1584),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1628),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1641),
.B(n_1592),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1643),
.B(n_1592),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1635),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1671),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1628),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1663),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1626),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1659),
.B(n_1599),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1605),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1666),
.B(n_1605),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1581),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1621),
.A2(n_1542),
.B(n_1538),
.C(n_1615),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_1658),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1706),
.B(n_1602),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1706),
.B(n_1602),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1706),
.B(n_1619),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1661),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1686),
.B(n_1630),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_R g1719 ( 
.A(n_1701),
.B(n_1703),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1707),
.B(n_1619),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1707),
.B(n_1619),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1674),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1707),
.B(n_1619),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1682),
.B(n_1581),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1692),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1703),
.A2(n_1622),
.B1(n_1627),
.B2(n_1625),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1688),
.B(n_1612),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1704),
.B(n_1633),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1619),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1673),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1682),
.B(n_1582),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1678),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1673),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1703),
.A2(n_1627),
.B(n_1622),
.C(n_1647),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1678),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1640),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1582),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1693),
.B(n_1619),
.Y(n_1740)
);

AOI32xp33_ASAP7_75t_L g1741 ( 
.A1(n_1701),
.A2(n_1624),
.A3(n_1653),
.B1(n_1649),
.B2(n_1660),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1673),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1679),
.B(n_1653),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1683),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1678),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1693),
.B(n_1568),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1675),
.B(n_1612),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1677),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1708),
.B(n_1582),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1678),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1571),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1677),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1675),
.B(n_1612),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1692),
.B(n_1571),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1680),
.Y(n_1755)
);

AND2x2_ASAP7_75t_SL g1756 ( 
.A(n_1688),
.B(n_1597),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1744),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1729),
.B(n_1698),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1719),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1731),
.Y(n_1760)
);

OAI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1727),
.A2(n_1688),
.B(n_1698),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1744),
.B(n_1710),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1731),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1737),
.B(n_1511),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1718),
.B(n_1695),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1734),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1734),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1742),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1756),
.B(n_1705),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1717),
.B(n_1684),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1727),
.B(n_1702),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1705),
.Y(n_1772)
);

NAND2x1_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1710),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1756),
.B(n_1705),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1733),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1742),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1755),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1755),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_1684),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1726),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1738),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1711),
.Y(n_1784)
);

NAND2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1746),
.B(n_1691),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1735),
.B(n_1679),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1676),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1739),
.B(n_1676),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1728),
.B(n_1683),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1748),
.B(n_1679),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1689),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1752),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1683),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1730),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1689),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1733),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1736),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1740),
.B(n_1699),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1749),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1740),
.B(n_1699),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_SL g1801 ( 
.A(n_1741),
.B(n_1690),
.C(n_1691),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1749),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1728),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1801),
.B(n_1701),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1785),
.B(n_1713),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1761),
.A2(n_1741),
.B(n_1728),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1783),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1773),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1764),
.B(n_1468),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1782),
.B(n_1751),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1763),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1770),
.B(n_1701),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1781),
.B(n_1700),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1771),
.A2(n_1758),
.B1(n_1786),
.B2(n_1765),
.C(n_1784),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1713),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1763),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1757),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1766),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1769),
.A2(n_1728),
.B1(n_1694),
.B2(n_1690),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_1714),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1773),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1759),
.A2(n_1769),
.B1(n_1774),
.B2(n_1772),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1772),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1757),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1766),
.Y(n_1825)
);

AND2x4_ASAP7_75t_SL g1826 ( 
.A(n_1774),
.B(n_1728),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1780),
.B(n_1751),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1757),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1794),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1775),
.B(n_1714),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1798),
.B(n_1725),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1775),
.B(n_1715),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1789),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1762),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1712),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1800),
.B(n_1725),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_1715),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1799),
.B(n_1361),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1791),
.B(n_1732),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1802),
.B(n_1700),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1804),
.A2(n_1793),
.B1(n_1694),
.B2(n_1762),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1804),
.A2(n_1637),
.B1(n_1683),
.B2(n_1687),
.Y(n_1843)
);

OAI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1822),
.A2(n_1814),
.B(n_1806),
.Y(n_1844)
);

AOI22x1_ASAP7_75t_L g1845 ( 
.A1(n_1823),
.A2(n_1762),
.B1(n_1792),
.B2(n_1778),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1807),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1829),
.B(n_1795),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_SL g1848 ( 
.A(n_1822),
.B(n_1709),
.C(n_1657),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1811),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1812),
.B(n_1448),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1813),
.B(n_1760),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1811),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1810),
.B(n_1787),
.Y(n_1853)
);

NAND2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1803),
.B(n_1835),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1816),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1835),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1816),
.B(n_1777),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1838),
.B(n_1720),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1826),
.A2(n_1694),
.B1(n_1696),
.B2(n_1709),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1827),
.A2(n_1685),
.B(n_1687),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1803),
.B(n_1683),
.Y(n_1862)
);

OAI31xp33_ASAP7_75t_L g1863 ( 
.A1(n_1826),
.A2(n_1694),
.A3(n_1687),
.B(n_1685),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1818),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1825),
.Y(n_1865)
);

OAI31xp33_ASAP7_75t_L g1866 ( 
.A1(n_1826),
.A2(n_1685),
.A3(n_1696),
.B(n_1670),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1825),
.Y(n_1867)
);

OAI322xp33_ASAP7_75t_L g1868 ( 
.A1(n_1810),
.A2(n_1787),
.A3(n_1788),
.B1(n_1778),
.B2(n_1779),
.C1(n_1754),
.C2(n_1767),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1803),
.A2(n_1696),
.B1(n_1697),
.B2(n_1790),
.Y(n_1869)
);

AOI21x1_ASAP7_75t_L g1870 ( 
.A1(n_1808),
.A2(n_1768),
.B(n_1767),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1854),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_1839),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1849),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1846),
.B(n_1833),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1844),
.B(n_1833),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1854),
.B(n_1835),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1853),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1852),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1858),
.B(n_1838),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1855),
.Y(n_1880)
);

OAI21xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1866),
.A2(n_1827),
.B(n_1821),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1847),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1850),
.B(n_1861),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1870),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1851),
.B(n_1840),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1864),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1845),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1865),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1867),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1842),
.B(n_1834),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1869),
.B(n_1834),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_1809),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1857),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1871),
.B(n_1808),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1881),
.A2(n_1843),
.B(n_1868),
.Y(n_1895)
);

AOI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1881),
.A2(n_1887),
.B(n_1892),
.C(n_1875),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_SL g1897 ( 
.A(n_1871),
.B(n_1821),
.Y(n_1897)
);

AND4x1_ASAP7_75t_L g1898 ( 
.A(n_1876),
.B(n_1863),
.C(n_1859),
.D(n_1819),
.Y(n_1898)
);

O2A1O1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1882),
.A2(n_1860),
.B(n_1862),
.C(n_1857),
.Y(n_1899)
);

AOI31xp33_ASAP7_75t_L g1900 ( 
.A1(n_1877),
.A2(n_1876),
.A3(n_1872),
.B(n_1874),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1890),
.A2(n_1891),
.B(n_1884),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_SL g1902 ( 
.A(n_1880),
.B(n_1817),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1885),
.B(n_1851),
.Y(n_1903)
);

NAND2x1_ASAP7_75t_L g1904 ( 
.A(n_1879),
.B(n_1803),
.Y(n_1904)
);

NAND4xp75_ASAP7_75t_L g1905 ( 
.A(n_1890),
.B(n_1860),
.C(n_1815),
.D(n_1805),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1884),
.A2(n_1815),
.B1(n_1805),
.B2(n_1820),
.Y(n_1906)
);

OAI221xp5_ASAP7_75t_SL g1907 ( 
.A1(n_1891),
.A2(n_1883),
.B1(n_1885),
.B2(n_1879),
.C(n_1893),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1893),
.A2(n_1832),
.B(n_1834),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1880),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1900),
.B(n_1880),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1896),
.B(n_1878),
.C(n_1873),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1895),
.B(n_1878),
.C(n_1873),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_L g1913 ( 
.A(n_1907),
.B(n_1888),
.C(n_1886),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1904),
.Y(n_1914)
);

NAND4xp75_ASAP7_75t_L g1915 ( 
.A(n_1901),
.B(n_1889),
.C(n_1886),
.D(n_1888),
.Y(n_1915)
);

NAND4xp75_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1889),
.C(n_1820),
.D(n_1828),
.Y(n_1916)
);

NAND5xp2_ASAP7_75t_L g1917 ( 
.A(n_1899),
.B(n_1830),
.C(n_1841),
.D(n_1667),
.E(n_1832),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1905),
.B(n_1832),
.C(n_1824),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1903),
.B(n_1832),
.Y(n_1919)
);

NOR3xp33_ASAP7_75t_L g1920 ( 
.A(n_1910),
.B(n_1912),
.C(n_1909),
.Y(n_1920)
);

NAND4xp25_ASAP7_75t_L g1921 ( 
.A(n_1917),
.B(n_1897),
.C(n_1906),
.D(n_1898),
.Y(n_1921)
);

NAND4xp25_ASAP7_75t_L g1922 ( 
.A(n_1913),
.B(n_1897),
.C(n_1902),
.D(n_1817),
.Y(n_1922)
);

O2A1O1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1911),
.A2(n_1914),
.B(n_1918),
.C(n_1919),
.Y(n_1923)
);

NOR4xp25_ASAP7_75t_L g1924 ( 
.A(n_1915),
.B(n_1824),
.C(n_1828),
.D(n_1840),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1916),
.B(n_1830),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1926),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1925),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1920),
.A2(n_1836),
.B1(n_1448),
.B2(n_1779),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1922),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1923),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1924),
.B(n_1831),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1921),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1932),
.A2(n_1837),
.B1(n_1831),
.B2(n_1788),
.C(n_1768),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1930),
.A2(n_1836),
.B1(n_1797),
.B2(n_1776),
.Y(n_1935)
);

OAI222xp33_ASAP7_75t_L g1936 ( 
.A1(n_1931),
.A2(n_1836),
.B1(n_1837),
.B2(n_1754),
.C1(n_1796),
.C2(n_1776),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1928),
.A2(n_1836),
.B(n_1797),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1927),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1933),
.B(n_1796),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1937),
.A2(n_1929),
.B(n_1716),
.Y(n_1940)
);

OR3x2_ASAP7_75t_L g1941 ( 
.A(n_1938),
.B(n_1929),
.C(n_1732),
.Y(n_1941)
);

XOR2x1_ASAP7_75t_SL g1942 ( 
.A(n_1939),
.B(n_1736),
.Y(n_1942)
);

NAND5xp2_ASAP7_75t_L g1943 ( 
.A(n_1934),
.B(n_1616),
.C(n_1697),
.D(n_1747),
.E(n_1753),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1943),
.A2(n_1935),
.B1(n_1936),
.B2(n_1681),
.Y(n_1944)
);

OAI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1944),
.A2(n_1940),
.B(n_1941),
.C(n_1942),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1745),
.B1(n_1750),
.B2(n_1716),
.Y(n_1946)
);

AO22x2_ASAP7_75t_L g1947 ( 
.A1(n_1945),
.A2(n_1722),
.B1(n_1723),
.B2(n_1712),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1947),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1946),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1949),
.A2(n_1721),
.B(n_1720),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1948),
.A2(n_1724),
.B(n_1721),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1951),
.A2(n_1750),
.B1(n_1745),
.B2(n_1722),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1950),
.B1(n_1436),
.B2(n_1439),
.Y(n_1953)
);

OAI221xp5_ASAP7_75t_R g1954 ( 
.A1(n_1953),
.A2(n_1436),
.B1(n_1439),
.B2(n_1681),
.C(n_1415),
.Y(n_1954)
);

AOI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1341),
.B(n_1419),
.C(n_1723),
.Y(n_1955)
);


endmodule