module fake_jpeg_2304_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_70),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_82),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_52),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_54),
.C(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_67),
.B1(n_50),
.B2(n_54),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_100),
.B1(n_104),
.B2(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_56),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_101),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_56),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_50),
.B1(n_66),
.B2(n_49),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_64),
.CI(n_57),
.CON(n_101),
.SN(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_53),
.B1(n_63),
.B2(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_22),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_87),
.B(n_81),
.C(n_65),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_12),
.B(n_13),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_81),
.B1(n_65),
.B2(n_20),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_10),
.Y(n_145)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_18),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_1),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_93),
.C(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_136),
.C(n_129),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_25),
.C(n_46),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_3),
.B(n_5),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_150),
.C(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_27),
.B1(n_44),
.B2(n_43),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_149),
.B1(n_154),
.B2(n_152),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_144),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_145),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_28),
.B(n_39),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_11),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_14),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_31),
.B1(n_37),
.B2(n_36),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_47),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_11),
.B(n_12),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_127),
.B(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_165),
.B1(n_170),
.B2(n_136),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_153),
.C(n_150),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_123),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_164),
.B(n_167),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_146),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_127),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_144),
.B(n_16),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_140),
.B(n_133),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_125),
.B(n_15),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_14),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_166),
.B1(n_157),
.B2(n_176),
.Y(n_185)
);

OAI31xp33_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_188),
.A3(n_155),
.B(n_174),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_159),
.B(n_158),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_182),
.B1(n_187),
.B2(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_173),
.B(n_33),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_17),
.C(n_34),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_35),
.Y(n_194)
);


endmodule