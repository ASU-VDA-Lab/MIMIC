module fake_jpeg_31907_n_498 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_498);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_498;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_71),
.Y(n_101)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_22),
.B(n_10),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_11),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_83),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_11),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_11),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_98),
.Y(n_145)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_22),
.B(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_34),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_56),
.B(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_151),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_46),
.B1(n_25),
.B2(n_45),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_106),
.A2(n_136),
.B1(n_98),
.B2(n_84),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_134),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_31),
.B1(n_18),
.B2(n_32),
.Y(n_131)
);

OA22x2_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_98),
.B1(n_84),
.B2(n_99),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_26),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_53),
.A2(n_46),
.B1(n_25),
.B2(n_45),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_30),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_155),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_75),
.A2(n_24),
.B1(n_45),
.B2(n_25),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_146),
.B1(n_31),
.B2(n_48),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_75),
.A2(n_24),
.B1(n_45),
.B2(n_25),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_52),
.B(n_30),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_99),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_78),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_38),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_162),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_167),
.Y(n_250)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_168),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_44),
.B(n_41),
.C(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_169),
.B(n_170),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_172),
.B(n_177),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_66),
.B1(n_61),
.B2(n_55),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_175),
.B1(n_191),
.B2(n_106),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_142),
.B1(n_147),
.B2(n_117),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_186),
.B1(n_206),
.B2(n_130),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_60),
.B1(n_59),
.B2(n_86),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_89),
.B1(n_88),
.B2(n_80),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_178),
.A2(n_184),
.B1(n_201),
.B2(n_202),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_192),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_103),
.A2(n_67),
.B1(n_27),
.B2(n_44),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_180),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_58),
.C(n_36),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_122),
.C(n_157),
.Y(n_230)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_64),
.B1(n_57),
.B2(n_45),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_109),
.A2(n_32),
.B1(n_28),
.B2(n_41),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_130),
.B1(n_115),
.B2(n_149),
.Y(n_223)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_112),
.A2(n_28),
.B1(n_64),
.B2(n_48),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_197),
.B(n_200),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_210),
.Y(n_217)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_18),
.B1(n_62),
.B2(n_57),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_131),
.A2(n_62),
.B1(n_18),
.B2(n_25),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_103),
.A2(n_18),
.B1(n_47),
.B2(n_12),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_101),
.A2(n_18),
.B1(n_47),
.B2(n_13),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_150),
.A2(n_18),
.B1(n_47),
.B2(n_13),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_121),
.B(n_145),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_100),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_0),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_123),
.A2(n_47),
.B1(n_6),
.B2(n_13),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_0),
.Y(n_241)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_131),
.A2(n_47),
.B(n_6),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_5),
.B(n_16),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_219),
.A2(n_226),
.B1(n_231),
.B2(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_222),
.B(n_165),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_223),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_137),
.B(n_152),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_227),
.A2(n_199),
.B(n_196),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_157),
.B1(n_149),
.B2(n_115),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_122),
.C(n_126),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_5),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_189),
.B(n_186),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_241),
.A2(n_165),
.B1(n_172),
.B2(n_170),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_0),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_166),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_257),
.B1(n_261),
.B2(n_3),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_1),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_176),
.B(n_1),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_214),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_215),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_216),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_163),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_279),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_176),
.C(n_201),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_275),
.C(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_189),
.B1(n_169),
.B2(n_159),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_160),
.B(n_190),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_247),
.B(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_187),
.C(n_185),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_277),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_244),
.B(n_193),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_249),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_237),
.B(n_183),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_290),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_235),
.B(n_194),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_292),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_217),
.B(n_188),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_218),
.A2(n_161),
.B1(n_184),
.B2(n_200),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_301),
.B1(n_224),
.B2(n_228),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_289),
.A2(n_291),
.B(n_245),
.Y(n_318)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_227),
.A2(n_179),
.A3(n_181),
.B1(n_213),
.B2(n_171),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_217),
.B(n_198),
.C(n_208),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_197),
.C(n_168),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_275),
.Y(n_309)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_295),
.B(n_300),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_164),
.B1(n_204),
.B2(n_167),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_259),
.B(n_4),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_302),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_260),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_218),
.A2(n_260),
.B1(n_236),
.B2(n_223),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_226),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_252),
.B(n_14),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_223),
.B1(n_219),
.B2(n_221),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_304),
.A2(n_307),
.B1(n_327),
.B2(n_328),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_319),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_223),
.B1(n_261),
.B2(n_231),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_239),
.B1(n_221),
.B2(n_257),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_308),
.A2(n_317),
.B1(n_320),
.B2(n_336),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_309),
.B(n_294),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_264),
.A2(n_229),
.B1(n_255),
.B2(n_232),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_318),
.A2(n_323),
.B(n_331),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_287),
.A2(n_224),
.B1(n_234),
.B2(n_232),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_336),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_296),
.A2(n_225),
.B1(n_247),
.B2(n_228),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_225),
.B1(n_228),
.B2(n_242),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_216),
.B1(n_256),
.B2(n_250),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_329),
.A2(n_286),
.B1(n_285),
.B2(n_293),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_289),
.A2(n_251),
.B(n_250),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_285),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_335),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_256),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_300),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_262),
.B(n_243),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_262),
.C(n_267),
.Y(n_342)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_350),
.C(n_353),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_284),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_326),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_349),
.Y(n_373)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_348),
.B1(n_368),
.B2(n_371),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_307),
.A2(n_306),
.B1(n_329),
.B2(n_335),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_325),
.B(n_288),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_288),
.Y(n_350)
);

AO22x1_ASAP7_75t_L g352 ( 
.A1(n_318),
.A2(n_340),
.B1(n_336),
.B2(n_317),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_358),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_285),
.C(n_292),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_362),
.B1(n_365),
.B2(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_311),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_273),
.C(n_265),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_363),
.C(n_316),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_276),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_372),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_251),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_361),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_291),
.B1(n_301),
.B2(n_302),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_297),
.Y(n_363)
);

AOI322xp5_ASAP7_75t_L g364 ( 
.A1(n_314),
.A2(n_271),
.A3(n_272),
.B1(n_270),
.B2(n_268),
.C1(n_295),
.C2(n_290),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_364),
.B(n_319),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_280),
.B1(n_274),
.B2(n_281),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_306),
.A2(n_263),
.B1(n_243),
.B2(n_17),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_369),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_316),
.B(n_243),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_243),
.B1(n_15),
.B2(n_16),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_352),
.A2(n_351),
.B1(n_358),
.B2(n_372),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_376),
.A2(n_380),
.B(n_391),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_393),
.C(n_395),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_323),
.C(n_331),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_381),
.B(n_394),
.C(n_397),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_341),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_322),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_387),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g385 ( 
.A1(n_352),
.A2(n_348),
.A3(n_351),
.B1(n_347),
.B2(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_330),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_367),
.A2(n_328),
.B1(n_334),
.B2(n_332),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_391),
.A2(n_355),
.B1(n_362),
.B2(n_354),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_366),
.A2(n_330),
.B(n_334),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_392),
.A2(n_357),
.B(n_346),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_326),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_350),
.B(n_327),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_332),
.C(n_337),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_337),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_400),
.C(n_363),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_313),
.C(n_312),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_389),
.B(n_345),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_401),
.Y(n_435)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_386),
.A2(n_367),
.B1(n_357),
.B2(n_368),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_407),
.A2(n_421),
.B1(n_395),
.B2(n_377),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_378),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_365),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_412),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_380),
.B1(n_382),
.B2(n_373),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_357),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_371),
.B(n_313),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_422),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_310),
.C(n_16),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_423),
.C(n_373),
.Y(n_425)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_419),
.A2(n_424),
.B1(n_402),
.B2(n_413),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_310),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_385),
.A2(n_310),
.B1(n_375),
.B2(n_381),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_399),
.A2(n_392),
.B(n_375),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_397),
.C(n_393),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_406),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_428),
.A2(n_402),
.B1(n_421),
.B2(n_422),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_384),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_433),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_400),
.C(n_394),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_437),
.C(n_418),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_387),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_434),
.A2(n_438),
.B1(n_407),
.B2(n_414),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_404),
.C(n_406),
.Y(n_437)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_448),
.C(n_451),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_428),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_401),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_409),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_454),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_418),
.C(n_416),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_452),
.A2(n_441),
.B1(n_427),
.B2(n_403),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_420),
.B(n_419),
.C(n_412),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_453),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_443),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_424),
.C(n_417),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_458),
.C(n_433),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_440),
.B(n_410),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_434),
.B1(n_425),
.B2(n_442),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_408),
.C(n_405),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_446),
.A2(n_426),
.B1(n_438),
.B2(n_429),
.Y(n_459)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_464),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_449),
.A2(n_415),
.B1(n_411),
.B2(n_439),
.Y(n_461)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_470),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_452),
.A2(n_440),
.B(n_430),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_458),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_448),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_476),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_451),
.C(n_455),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_473),
.B(n_477),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_450),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_462),
.C(n_464),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_477),
.B(n_473),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_453),
.Y(n_479)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_479),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_485),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_475),
.B(n_467),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_467),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_465),
.C(n_466),
.Y(n_490)
);

A2O1A1O1Ixp25_ASAP7_75t_L g489 ( 
.A1(n_486),
.A2(n_480),
.B(n_474),
.C(n_459),
.D(n_465),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_489),
.A2(n_466),
.B(n_483),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_491),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_481),
.C(n_463),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_488),
.Y(n_494)
);

AO21x1_ASAP7_75t_L g495 ( 
.A1(n_494),
.A2(n_493),
.B(n_470),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_481),
.C(n_463),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_496),
.A2(n_456),
.B(n_431),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_456),
.Y(n_498)
);


endmodule