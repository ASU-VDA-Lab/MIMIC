module fake_jpeg_19574_n_288 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_SL g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_24),
.B1(n_31),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_47),
.B1(n_35),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_16),
.B1(n_24),
.B2(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_16),
.B1(n_35),
.B2(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

OR2x4_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_75),
.B1(n_23),
.B2(n_43),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_16),
.A3(n_38),
.B1(n_22),
.B2(n_12),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_36),
.B(n_43),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_34),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_54),
.B1(n_43),
.B2(n_39),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_93),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_89),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_39),
.B1(n_59),
.B2(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_39),
.B1(n_51),
.B2(n_37),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_97),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_63),
.B1(n_81),
.B2(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_21),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_57),
.B1(n_50),
.B2(n_44),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_100),
.B1(n_66),
.B2(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_53),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_36),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_66),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_33),
.B1(n_32),
.B2(n_26),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_96),
.B1(n_93),
.B2(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_18),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_65),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_118),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_80),
.A3(n_74),
.B1(n_68),
.B2(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_122),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_64),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_68),
.C(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_76),
.B1(n_70),
.B2(n_12),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_18),
.B1(n_28),
.B2(n_15),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_125),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_76),
.B1(n_34),
.B2(n_26),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_95),
.B(n_99),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_140),
.B1(n_153),
.B2(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_99),
.B1(n_89),
.B2(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_145),
.B1(n_147),
.B2(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_76),
.B1(n_82),
.B2(n_64),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_101),
.B(n_113),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_23),
.B(n_22),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_14),
.B1(n_34),
.B2(n_29),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_14),
.B1(n_29),
.B2(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_17),
.Y(n_150)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_124),
.B1(n_121),
.B2(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_106),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_124),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_134),
.B1(n_154),
.B2(n_132),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_17),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_15),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_15),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_15),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_178),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_182),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_133),
.B(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_137),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_145),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_152),
.C(n_128),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_187),
.C(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_152),
.C(n_128),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_196),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_132),
.C(n_135),
.D(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_205),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_133),
.B1(n_151),
.B2(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_131),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_204),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_138),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_202),
.B1(n_177),
.B2(n_158),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_137),
.C(n_139),
.Y(n_201)
);

AOI22x1_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_155),
.B1(n_147),
.B2(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_143),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_144),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_202),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_183),
.C(n_162),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_220),
.C(n_221),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_171),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_5),
.C(n_9),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_173),
.B1(n_181),
.B2(n_171),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_183),
.C(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_168),
.C(n_181),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_174),
.B(n_165),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_189),
.B(n_203),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_158),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_224),
.C(n_19),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_200),
.C(n_192),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_20),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_224),
.C(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_5),
.B1(n_9),
.B2(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_239),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_208),
.B(n_217),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_206),
.B(n_218),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_10),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_216),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_248),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_228),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_6),
.B(n_7),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_237),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_259),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_257),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_238),
.B(n_6),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_260),
.B(n_0),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_9),
.C(n_7),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_10),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_248),
.B1(n_243),
.B2(n_2),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_247),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_0),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_0),
.B(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_0),
.B(n_1),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_1),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_278),
.B(n_279),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_1),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_266),
.B(n_3),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_281),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_2),
.B(n_3),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_282),
.Y(n_284)
);

OAI321xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_276),
.C(n_283),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_4),
.B(n_2),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_3),
.Y(n_288)
);


endmodule