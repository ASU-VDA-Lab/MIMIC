module real_aes_17608_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_559;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_729;
wire n_394;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g405 ( .A(n_0), .Y(n_405) );
INVx1_ASAP7_75t_L g648 ( .A(n_1), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_2), .A2(n_160), .B1(n_373), .B2(n_670), .Y(n_777) );
OAI22xp33_ASAP7_75t_SL g790 ( .A1(n_2), .A2(n_160), .B1(n_283), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g863 ( .A(n_3), .Y(n_863) );
OAI211xp5_ASAP7_75t_L g867 ( .A1(n_3), .A2(n_544), .B(n_779), .C(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g1389 ( .A(n_4), .Y(n_1389) );
AOI22xp5_ASAP7_75t_SL g1083 ( .A1(n_5), .A2(n_231), .B1(n_1076), .B2(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g616 ( .A(n_6), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g1296 ( .A1(n_7), .A2(n_179), .B1(n_1297), .B2(n_1298), .C(n_1299), .Y(n_1296) );
INVx1_ASAP7_75t_L g1351 ( .A(n_7), .Y(n_1351) );
INVx1_ASAP7_75t_L g262 ( .A(n_8), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_8), .B(n_272), .Y(n_425) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_8), .B(n_364), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_8), .B(n_208), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_9), .A2(n_190), .B1(n_264), .B2(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_9), .A2(n_190), .B1(n_281), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_10), .A2(n_212), .B1(n_556), .B2(n_560), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_10), .A2(n_49), .B1(n_584), .B2(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g822 ( .A(n_11), .Y(n_822) );
OAI222xp33_ASAP7_75t_L g526 ( .A1(n_12), .A2(n_192), .B1(n_473), .B2(n_527), .C1(n_529), .C2(n_533), .Y(n_526) );
OAI222xp33_ASAP7_75t_L g567 ( .A1(n_12), .A2(n_129), .B1(n_192), .B2(n_568), .C1(n_569), .C2(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g978 ( .A(n_13), .Y(n_978) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_14), .B(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1074 ( .A(n_14), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_14), .B(n_95), .Y(n_1079) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_15), .A2(n_236), .B1(n_525), .B2(n_912), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_15), .A2(n_19), .B1(n_927), .B2(n_930), .Y(n_936) );
OAI22xp5_ASAP7_75t_SL g839 ( .A1(n_16), .A2(n_127), .B1(n_361), .B2(n_505), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_16), .A2(n_127), .B1(n_843), .B2(n_844), .Y(n_842) );
INVx1_ASAP7_75t_L g945 ( .A(n_17), .Y(n_945) );
AO22x2_ASAP7_75t_L g742 ( .A1(n_18), .A2(n_743), .B1(n_798), .B2(n_799), .Y(n_742) );
INVx1_ASAP7_75t_L g798 ( .A(n_18), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_19), .A2(n_163), .B1(n_560), .B2(n_916), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_20), .A2(n_199), .B1(n_283), .B2(n_650), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_20), .A2(n_242), .B1(n_492), .B2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_SL g1098 ( .A1(n_21), .A2(n_118), .B1(n_1076), .B2(n_1084), .Y(n_1098) );
INVx1_ASAP7_75t_L g1386 ( .A(n_22), .Y(n_1386) );
INVx1_ASAP7_75t_L g810 ( .A(n_23), .Y(n_810) );
INVx1_ASAP7_75t_L g545 ( .A(n_24), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_24), .A2(n_212), .B1(n_587), .B2(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g1045 ( .A1(n_25), .A2(n_138), .B1(n_373), .B2(n_786), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_25), .A2(n_239), .B1(n_283), .B2(n_643), .Y(n_1047) );
AOI22xp5_ASAP7_75t_SL g1088 ( .A1(n_26), .A2(n_226), .B1(n_1060), .B2(n_1078), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_27), .A2(n_156), .B1(n_264), .B2(n_373), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_27), .A2(n_156), .B1(n_643), .B2(n_949), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_28), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_29), .A2(n_124), .B1(n_492), .B2(n_670), .Y(n_1366) );
OAI22xp33_ASAP7_75t_SL g1368 ( .A1(n_29), .A2(n_124), .B1(n_283), .B2(n_791), .Y(n_1368) );
INVx1_ASAP7_75t_L g749 ( .A(n_30), .Y(n_749) );
INVx1_ASAP7_75t_L g389 ( .A(n_31), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_32), .A2(n_159), .B1(n_1060), .B2(n_1072), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_33), .A2(n_153), .B1(n_264), .B2(n_373), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_33), .A2(n_153), .B1(n_290), .B2(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g885 ( .A(n_34), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_35), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_36), .Y(n_1026) );
XOR2x2_ASAP7_75t_L g907 ( .A(n_37), .B(n_908), .Y(n_907) );
XNOR2xp5_ASAP7_75t_L g804 ( .A(n_38), .B(n_805), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_39), .A2(n_162), .B1(n_325), .B2(n_643), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_39), .A2(n_41), .B1(n_668), .B2(n_786), .Y(n_986) );
INVx1_ASAP7_75t_L g941 ( .A(n_40), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_41), .A2(n_246), .B1(n_283), .B2(n_322), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_42), .A2(n_161), .B1(n_1076), .B2(n_1078), .Y(n_1075) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_43), .A2(n_79), .B1(n_1072), .B2(n_1076), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_44), .A2(n_90), .B1(n_1076), .B2(n_1094), .Y(n_1164) );
INVx1_ASAP7_75t_L g1364 ( .A(n_45), .Y(n_1364) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_46), .A2(n_117), .B1(n_281), .B2(n_290), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_46), .A2(n_117), .B1(n_264), .B2(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g287 ( .A(n_47), .Y(n_287) );
INVx1_ASAP7_75t_L g303 ( .A(n_47), .Y(n_303) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_48), .A2(n_224), .B1(n_1264), .B2(n_1268), .C(n_1271), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_48), .A2(n_110), .B1(n_1337), .B2(n_1340), .Y(n_1336) );
INVx1_ASAP7_75t_L g546 ( .A(n_49), .Y(n_546) );
INVx1_ASAP7_75t_L g474 ( .A(n_50), .Y(n_474) );
XOR2xp5_ASAP7_75t_L g598 ( .A(n_51), .B(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g1110 ( .A1(n_51), .A2(n_241), .B1(n_1060), .B2(n_1072), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_52), .A2(n_99), .B1(n_786), .B2(n_787), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_52), .A2(n_99), .B1(n_322), .B2(n_325), .Y(n_796) );
INVx1_ASAP7_75t_L g460 ( .A(n_53), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_54), .A2(n_183), .B1(n_697), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_54), .A2(n_189), .B1(n_721), .B2(n_725), .Y(n_727) );
INVx1_ASAP7_75t_L g255 ( .A(n_55), .Y(n_255) );
INVx1_ASAP7_75t_L g813 ( .A(n_56), .Y(n_813) );
INVx2_ASAP7_75t_L g289 ( .A(n_57), .Y(n_289) );
XNOR2x2_ASAP7_75t_L g452 ( .A(n_58), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g605 ( .A(n_59), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_60), .A2(n_207), .B1(n_504), .B2(n_505), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g513 ( .A1(n_60), .A2(n_207), .B1(n_321), .B2(n_323), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_61), .A2(n_223), .B1(n_596), .B2(n_952), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_61), .A2(n_165), .B1(n_551), .B2(n_1002), .Y(n_1003) );
AOI211xp5_ASAP7_75t_L g1281 ( .A1(n_62), .A2(n_967), .B(n_1282), .C(n_1286), .Y(n_1281) );
INVx1_ASAP7_75t_L g1349 ( .A(n_62), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_63), .A2(n_66), .B1(n_1072), .B2(n_1076), .Y(n_1089) );
INVx1_ASAP7_75t_L g977 ( .A(n_64), .Y(n_977) );
INVx1_ASAP7_75t_L g975 ( .A(n_65), .Y(n_975) );
INVx1_ASAP7_75t_L g462 ( .A(n_67), .Y(n_462) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_68), .A2(n_100), .B1(n_218), .B2(n_686), .C1(n_688), .C2(n_689), .Y(n_685) );
OAI222xp33_ASAP7_75t_L g737 ( .A1(n_68), .A2(n_100), .B1(n_218), .B2(n_355), .C1(n_738), .C2(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g891 ( .A(n_69), .Y(n_891) );
INVx1_ASAP7_75t_L g1381 ( .A(n_70), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_71), .A2(n_247), .B1(n_703), .B2(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_71), .A2(n_115), .B1(n_729), .B2(n_730), .Y(n_728) );
XOR2xp5_ASAP7_75t_L g518 ( .A(n_72), .B(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_73), .A2(n_115), .B1(n_710), .B2(n_711), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_73), .A2(n_247), .B1(n_721), .B2(n_725), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g962 ( .A1(n_74), .A2(n_244), .B1(n_711), .B2(n_828), .C(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_74), .A2(n_114), .B1(n_730), .B2(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1363 ( .A(n_75), .Y(n_1363) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_76), .A2(n_196), .B1(n_560), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_76), .A2(n_78), .B1(n_396), .B2(n_933), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g1105 ( .A1(n_77), .A2(n_170), .B1(n_1060), .B2(n_1084), .Y(n_1105) );
AOI222xp33_ASAP7_75t_L g1253 ( .A1(n_77), .A2(n_1254), .B1(n_1352), .B2(n_1355), .C1(n_1399), .C2(n_1401), .Y(n_1253) );
XOR2x2_ASAP7_75t_L g1254 ( .A(n_77), .B(n_1255), .Y(n_1254) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_78), .A2(n_151), .B1(n_525), .B2(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g457 ( .A(n_80), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g493 ( .A1(n_81), .A2(n_494), .B(n_497), .C(n_502), .Y(n_493) );
INVx1_ASAP7_75t_L g512 ( .A(n_81), .Y(n_512) );
INVx1_ASAP7_75t_L g817 ( .A(n_82), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_83), .A2(n_110), .B1(n_1291), .B2(n_1294), .Y(n_1290) );
OAI211xp5_ASAP7_75t_L g1305 ( .A1(n_83), .A2(n_1306), .B(n_1311), .C(n_1326), .Y(n_1305) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_84), .A2(n_242), .B1(n_322), .B2(n_643), .C(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g666 ( .A(n_84), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_85), .A2(n_152), .B1(n_668), .B2(n_786), .Y(n_1365) );
OAI22xp33_ASAP7_75t_L g1374 ( .A1(n_85), .A2(n_152), .B1(n_322), .B2(n_325), .Y(n_1374) );
INVx1_ASAP7_75t_L g397 ( .A(n_86), .Y(n_397) );
INVx1_ASAP7_75t_L g1289 ( .A(n_87), .Y(n_1289) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_88), .Y(n_257) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_88), .B(n_255), .Y(n_1061) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_89), .A2(n_522), .B(n_523), .C(n_534), .Y(n_521) );
INVx1_ASAP7_75t_L g576 ( .A(n_89), .Y(n_576) );
INVx1_ASAP7_75t_L g607 ( .A(n_91), .Y(n_607) );
INVx1_ASAP7_75t_L g1301 ( .A(n_92), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1092 ( .A1(n_93), .A2(n_137), .B1(n_1060), .B2(n_1072), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_94), .A2(n_157), .B1(n_321), .B2(n_844), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_94), .A2(n_157), .B1(n_504), .B2(n_505), .Y(n_871) );
INVx1_ASAP7_75t_L g1063 ( .A(n_95), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_95), .B(n_1074), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_96), .A2(n_168), .B1(n_1060), .B2(n_1072), .Y(n_1085) );
INVx1_ASAP7_75t_L g1284 ( .A(n_97), .Y(n_1284) );
INVx1_ASAP7_75t_L g1300 ( .A(n_98), .Y(n_1300) );
INVx1_ASAP7_75t_L g608 ( .A(n_101), .Y(n_608) );
INVx1_ASAP7_75t_L g765 ( .A(n_102), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_103), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_104), .A2(n_210), .B1(n_650), .B2(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_104), .A2(n_210), .B1(n_504), .B2(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g332 ( .A(n_105), .Y(n_332) );
INVx1_ASAP7_75t_L g413 ( .A(n_105), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_105), .B(n_289), .Y(n_1277) );
INVx1_ASAP7_75t_L g862 ( .A(n_106), .Y(n_862) );
INVx1_ASAP7_75t_L g1379 ( .A(n_107), .Y(n_1379) );
INVx1_ASAP7_75t_L g837 ( .A(n_108), .Y(n_837) );
INVx1_ASAP7_75t_L g679 ( .A(n_109), .Y(n_679) );
INVx1_ASAP7_75t_L g419 ( .A(n_111), .Y(n_419) );
INVx1_ASAP7_75t_L g781 ( .A(n_112), .Y(n_781) );
INVx1_ASAP7_75t_L g1388 ( .A(n_113), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_114), .A2(n_202), .B1(n_711), .B2(n_828), .C(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g880 ( .A(n_116), .Y(n_880) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_119), .B(n_676), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_120), .Y(n_1042) );
INVx1_ASAP7_75t_L g883 ( .A(n_121), .Y(n_883) );
INVx1_ASAP7_75t_L g1163 ( .A(n_122), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_123), .A2(n_132), .B1(n_1274), .B2(n_1278), .Y(n_1273) );
INVxp67_ASAP7_75t_SL g1327 ( .A(n_123), .Y(n_1327) );
INVx1_ASAP7_75t_L g532 ( .A(n_125), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_125), .A2(n_206), .B1(n_322), .B2(n_325), .Y(n_573) );
INVx1_ASAP7_75t_L g763 ( .A(n_126), .Y(n_763) );
AOI31xp33_ASAP7_75t_L g959 ( .A1(n_128), .A2(n_960), .A3(n_971), .B(n_980), .Y(n_959) );
NAND2xp33_ASAP7_75t_SL g996 ( .A(n_128), .B(n_997), .Y(n_996) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_128), .Y(n_1007) );
INVx1_ASAP7_75t_L g524 ( .A(n_129), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_130), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_131), .A2(n_167), .B1(n_1076), .B2(n_1094), .Y(n_1093) );
INVxp67_ASAP7_75t_SL g1318 ( .A(n_132), .Y(n_1318) );
BUFx3_ASAP7_75t_L g285 ( .A(n_133), .Y(n_285) );
INVx1_ASAP7_75t_L g387 ( .A(n_134), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_135), .Y(n_1027) );
INVx1_ASAP7_75t_L g458 ( .A(n_136), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_138), .A2(n_243), .B1(n_322), .B2(n_325), .Y(n_1051) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_139), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_140), .A2(n_198), .B1(n_1076), .B2(n_1084), .Y(n_1111) );
INVx1_ASAP7_75t_L g838 ( .A(n_141), .Y(n_838) );
OAI211xp5_ASAP7_75t_SL g845 ( .A1(n_141), .A2(n_305), .B(n_846), .C(n_848), .Y(n_845) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_142), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_143), .Y(n_541) );
INVx1_ASAP7_75t_L g647 ( .A(n_144), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_145), .A2(n_189), .B1(n_697), .B2(n_700), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_145), .A2(n_183), .B1(n_718), .B2(n_719), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_146), .A2(n_188), .B1(n_851), .B2(n_865), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_146), .A2(n_188), .B1(n_373), .B2(n_670), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_147), .Y(n_1015) );
INVx1_ASAP7_75t_L g760 ( .A(n_148), .Y(n_760) );
INVx1_ASAP7_75t_L g393 ( .A(n_149), .Y(n_393) );
INVx1_ASAP7_75t_L g751 ( .A(n_150), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_151), .A2(n_196), .B1(n_924), .B2(n_925), .Y(n_923) );
INVx1_ASAP7_75t_L g315 ( .A(n_154), .Y(n_315) );
INVx1_ASAP7_75t_L g469 ( .A(n_155), .Y(n_469) );
INVx1_ASAP7_75t_L g969 ( .A(n_158), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_158), .A2(n_223), .B1(n_560), .B2(n_1000), .Y(n_999) );
OA22x2_ASAP7_75t_L g853 ( .A1(n_159), .A2(n_854), .B1(n_903), .B2(n_904), .Y(n_853) );
INVxp67_ASAP7_75t_L g904 ( .A(n_159), .Y(n_904) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_162), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_163), .A2(n_236), .B1(n_927), .B2(n_930), .Y(n_926) );
INVx1_ASAP7_75t_L g620 ( .A(n_164), .Y(n_620) );
INVx1_ASAP7_75t_L g968 ( .A(n_165), .Y(n_968) );
INVx1_ASAP7_75t_L g943 ( .A(n_166), .Y(n_943) );
INVx1_ASAP7_75t_L g539 ( .A(n_169), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_169), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g820 ( .A(n_171), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_172), .B(n_313), .Y(n_646) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_172), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g297 ( .A1(n_173), .A2(n_298), .B(n_305), .C(n_309), .Y(n_297) );
INVx1_ASAP7_75t_L g359 ( .A(n_173), .Y(n_359) );
INVx1_ASAP7_75t_L g782 ( .A(n_174), .Y(n_782) );
OAI211xp5_ASAP7_75t_L g857 ( .A1(n_175), .A2(n_858), .B(n_860), .C(n_861), .Y(n_857) );
INVx1_ASAP7_75t_L g869 ( .A(n_175), .Y(n_869) );
INVx1_ASAP7_75t_L g877 ( .A(n_176), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_177), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_178), .A2(n_234), .B1(n_321), .B2(n_323), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_178), .A2(n_234), .B1(n_361), .B2(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g1345 ( .A(n_179), .Y(n_1345) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
XNOR2xp5_ASAP7_75t_L g1356 ( .A(n_181), .B(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g944 ( .A(n_182), .Y(n_944) );
INVx1_ASAP7_75t_L g818 ( .A(n_184), .Y(n_818) );
INVx1_ASAP7_75t_L g753 ( .A(n_185), .Y(n_753) );
INVx1_ASAP7_75t_L g1287 ( .A(n_186), .Y(n_1287) );
INVx1_ASAP7_75t_L g1043 ( .A(n_187), .Y(n_1043) );
OAI211xp5_ASAP7_75t_L g1048 ( .A1(n_187), .A2(n_416), .B(n_860), .C(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g614 ( .A(n_191), .Y(n_614) );
OAI211xp5_ASAP7_75t_SL g835 ( .A1(n_193), .A2(n_345), .B(n_494), .C(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g849 ( .A(n_193), .Y(n_849) );
INVx1_ASAP7_75t_L g1385 ( .A(n_194), .Y(n_1385) );
INVx1_ASAP7_75t_L g747 ( .A(n_195), .Y(n_747) );
INVx1_ASAP7_75t_L g501 ( .A(n_197), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_197), .A2(n_298), .B(n_305), .C(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_199), .Y(n_663) );
INVx1_ASAP7_75t_L g759 ( .A(n_200), .Y(n_759) );
INVx1_ASAP7_75t_L g940 ( .A(n_201), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_202), .A2(n_244), .B1(n_551), .B2(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1258 ( .A(n_203), .Y(n_1258) );
INVx1_ASAP7_75t_L g890 ( .A(n_204), .Y(n_890) );
INVx1_ASAP7_75t_L g1382 ( .A(n_205), .Y(n_1382) );
INVx1_ASAP7_75t_L g536 ( .A(n_206), .Y(n_536) );
BUFx3_ASAP7_75t_L g272 ( .A(n_208), .Y(n_272) );
INVx1_ASAP7_75t_L g364 ( .A(n_208), .Y(n_364) );
INVx1_ASAP7_75t_L g500 ( .A(n_209), .Y(n_500) );
XOR2x2_ASAP7_75t_L g277 ( .A(n_211), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g604 ( .A(n_213), .Y(n_604) );
INVx1_ASAP7_75t_L g886 ( .A(n_214), .Y(n_886) );
INVx1_ASAP7_75t_L g882 ( .A(n_215), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_216), .A2(n_444), .B(n_655), .C(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1050 ( .A(n_216), .Y(n_1050) );
INVx1_ASAP7_75t_L g407 ( .A(n_217), .Y(n_407) );
INVx1_ASAP7_75t_L g1378 ( .A(n_219), .Y(n_1378) );
INVx1_ASAP7_75t_L g784 ( .A(n_220), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g1360 ( .A1(n_221), .A2(n_655), .B(n_1361), .C(n_1362), .Y(n_1360) );
INVx1_ASAP7_75t_L g1371 ( .A(n_221), .Y(n_1371) );
INVx1_ASAP7_75t_L g337 ( .A(n_222), .Y(n_337) );
INVx1_ASAP7_75t_L g412 ( .A(n_222), .Y(n_412) );
INVx2_ASAP7_75t_L g424 ( .A(n_222), .Y(n_424) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_224), .Y(n_1325) );
AOI22xp5_ASAP7_75t_L g1097 ( .A1(n_225), .A2(n_237), .B1(n_1060), .B2(n_1072), .Y(n_1097) );
INVx1_ASAP7_75t_L g1162 ( .A(n_227), .Y(n_1162) );
INVx1_ASAP7_75t_L g618 ( .A(n_228), .Y(n_618) );
INVx1_ASAP7_75t_L g809 ( .A(n_229), .Y(n_809) );
INVx1_ASAP7_75t_L g475 ( .A(n_230), .Y(n_475) );
INVx1_ASAP7_75t_L g812 ( .A(n_232), .Y(n_812) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_233), .A2(n_551), .B(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g580 ( .A(n_233), .Y(n_580) );
INVx1_ASAP7_75t_L g415 ( .A(n_235), .Y(n_415) );
XNOR2xp5_ASAP7_75t_L g1010 ( .A(n_237), .B(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g319 ( .A(n_238), .Y(n_319) );
OAI211xp5_ASAP7_75t_L g339 ( .A1(n_238), .A2(n_340), .B(n_345), .C(n_350), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_239), .A2(n_243), .B1(n_367), .B2(n_670), .Y(n_1044) );
INVx1_ASAP7_75t_L g681 ( .A(n_240), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_245), .Y(n_530) );
INVx1_ASAP7_75t_L g982 ( .A(n_246), .Y(n_982) );
INVx1_ASAP7_75t_L g467 ( .A(n_248), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_273), .B(n_1056), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_258), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1354 ( .A(n_252), .B(n_261), .Y(n_1354) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_254), .B(n_257), .Y(n_1400) );
INVx1_ASAP7_75t_L g1405 ( .A(n_254), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_257), .B(n_1405), .Y(n_1407) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g378 ( .A(n_261), .B(n_379), .Y(n_378) );
AOI21xp5_ASAP7_75t_SL g520 ( .A1(n_261), .A2(n_521), .B(n_537), .Y(n_520) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g447 ( .A(n_262), .B(n_272), .Y(n_447) );
AND2x4_ASAP7_75t_L g554 ( .A(n_262), .B(n_271), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_263), .A2(n_374), .B1(n_679), .B2(n_681), .Y(n_733) );
AND2x4_ASAP7_75t_SL g1353 ( .A(n_263), .B(n_1354), .Y(n_1353) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_270), .Y(n_264) );
OR2x6_ASAP7_75t_L g362 ( .A(n_265), .B(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_L g540 ( .A(n_265), .Y(n_540) );
OR2x2_ASAP7_75t_L g786 ( .A(n_265), .B(n_363), .Y(n_786) );
INVx1_ASAP7_75t_L g1398 ( .A(n_265), .Y(n_1398) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx4f_ASAP7_75t_L g430 ( .A(n_266), .Y(n_430) );
INVx3_ASAP7_75t_L g473 ( .A(n_266), .Y(n_473) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2x1_ASAP7_75t_L g344 ( .A(n_268), .B(n_269), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_268), .B(n_269), .Y(n_349) );
INVx1_ASAP7_75t_L g358 ( .A(n_268), .Y(n_358) );
INVx2_ASAP7_75t_L g371 ( .A(n_268), .Y(n_371) );
AND2x2_ASAP7_75t_L g375 ( .A(n_268), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g439 ( .A(n_268), .Y(n_439) );
BUFx2_ASAP7_75t_L g353 ( .A(n_269), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_269), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g376 ( .A(n_269), .Y(n_376) );
OR2x2_ASAP7_75t_L g438 ( .A(n_269), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g559 ( .A(n_269), .Y(n_559) );
AND2x2_ASAP7_75t_L g561 ( .A(n_269), .B(n_371), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_270), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_529) );
OR2x6_ASAP7_75t_L g670 ( .A(n_270), .B(n_473), .Y(n_670) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g347 ( .A(n_271), .Y(n_347) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g352 ( .A(n_272), .Y(n_352) );
AND2x4_ASAP7_75t_L g356 ( .A(n_272), .B(n_357), .Y(n_356) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_672), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_515), .B1(n_516), .B2(n_671), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_451), .B(n_514), .Y(n_275) );
OA21x2_ASAP7_75t_L g671 ( .A1(n_276), .A2(n_451), .B(n_514), .Y(n_671) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g514 ( .A(n_277), .B(n_452), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_338), .C(n_381), .Y(n_278) );
OAI31xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_297), .A3(n_320), .B(n_328), .Y(n_279) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g575 ( .A(n_283), .Y(n_575) );
INVx2_ASAP7_75t_SL g680 ( .A(n_283), .Y(n_680) );
OR2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
OR2x4_ASAP7_75t_L g322 ( .A(n_284), .B(n_292), .Y(n_322) );
BUFx3_ASAP7_75t_L g388 ( .A(n_284), .Y(n_388) );
BUFx3_ASAP7_75t_L g481 ( .A(n_284), .Y(n_481) );
BUFx4f_ASAP7_75t_L g603 ( .A(n_284), .Y(n_603) );
INVx2_ASAP7_75t_L g1032 ( .A(n_284), .Y(n_1032) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g296 ( .A(n_285), .Y(n_296) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
AND2x4_ASAP7_75t_L g307 ( .A(n_285), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_285), .B(n_303), .Y(n_327) );
INVx1_ASAP7_75t_L g586 ( .A(n_286), .Y(n_586) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVxp67_ASAP7_75t_L g295 ( .A(n_287), .Y(n_295) );
INVx1_ASAP7_75t_L g292 ( .A(n_288), .Y(n_292) );
AND2x4_ASAP7_75t_L g306 ( .A(n_288), .B(n_307), .Y(n_306) );
OR2x6_ASAP7_75t_L g325 ( .A(n_288), .B(n_326), .Y(n_325) );
NAND3x1_ASAP7_75t_L g410 ( .A(n_288), .B(n_411), .C(n_413), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_288), .B(n_413), .Y(n_622) );
AND2x4_ASAP7_75t_L g1261 ( .A(n_288), .B(n_1262), .Y(n_1261) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
NAND2xp33_ASAP7_75t_SL g385 ( .A(n_289), .B(n_332), .Y(n_385) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g509 ( .A(n_291), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_291), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g791 ( .A(n_291), .Y(n_791) );
INVx1_ASAP7_75t_L g865 ( .A(n_291), .Y(n_865) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g577 ( .A(n_292), .B(n_293), .Y(n_577) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_293), .Y(n_582) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_293), .Y(n_828) );
INVx2_ASAP7_75t_L g830 ( .A(n_293), .Y(n_830) );
INVx2_ASAP7_75t_L g1034 ( .A(n_293), .Y(n_1034) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_294), .Y(n_396) );
INVx2_ASAP7_75t_L g594 ( .A(n_294), .Y(n_594) );
BUFx8_ASAP7_75t_L g613 ( .A(n_294), .Y(n_613) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x4_ASAP7_75t_L g585 ( .A(n_296), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g568 ( .A(n_299), .Y(n_568) );
INVx1_ASAP7_75t_L g688 ( .A(n_299), .Y(n_688) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g391 ( .A(n_300), .Y(n_391) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_300), .Y(n_619) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_300), .Y(n_825) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g418 ( .A(n_301), .Y(n_418) );
BUFx3_ASAP7_75t_L g484 ( .A(n_301), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
BUFx2_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g308 ( .A(n_303), .Y(n_308) );
BUFx2_ASAP7_75t_L g314 ( .A(n_304), .Y(n_314) );
AND2x4_ASAP7_75t_L g590 ( .A(n_304), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g1267 ( .A(n_304), .Y(n_1267) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_305), .B(n_793), .C(n_794), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g950 ( .A(n_305), .B(n_951), .C(n_954), .Y(n_950) );
CKINVDCx8_ASAP7_75t_R g305 ( .A(n_306), .Y(n_305) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_306), .B(n_567), .C(n_573), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_306), .B(n_683), .C(n_685), .Y(n_682) );
CKINVDCx8_ASAP7_75t_R g860 ( .A(n_306), .Y(n_860) );
BUFx2_ASAP7_75t_L g587 ( .A(n_307), .Y(n_587) );
BUFx2_ASAP7_75t_L g645 ( .A(n_307), .Y(n_645) );
INVx2_ASAP7_75t_L g701 ( .A(n_307), .Y(n_701) );
BUFx2_ASAP7_75t_L g795 ( .A(n_307), .Y(n_795) );
BUFx2_ASAP7_75t_L g952 ( .A(n_307), .Y(n_952) );
BUFx3_ASAP7_75t_L g967 ( .A(n_307), .Y(n_967) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_307), .B(n_1293), .Y(n_1295) );
INVx1_ASAP7_75t_L g591 ( .A(n_308), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_315), .B1(n_316), .B2(n_319), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_310), .A2(n_316), .B1(n_500), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_310), .A2(n_316), .B1(n_837), .B2(n_849), .Y(n_848) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g953 ( .A(n_311), .Y(n_953) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
AND2x4_ASAP7_75t_L g317 ( .A(n_312), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g570 ( .A(n_312), .B(n_314), .Y(n_570) );
AND2x2_ASAP7_75t_L g572 ( .A(n_312), .B(n_318), .Y(n_572) );
AND2x4_ASAP7_75t_L g687 ( .A(n_312), .B(n_314), .Y(n_687) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND3x4_ASAP7_75t_L g694 ( .A(n_313), .B(n_332), .C(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_313), .B(n_332), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_315), .A2(n_351), .B1(n_354), .B2(n_359), .Y(n_350) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g689 ( .A(n_317), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_317), .A2(n_687), .B1(n_781), .B2(n_784), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_317), .A2(n_687), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g951 ( .A1(n_317), .A2(n_943), .B1(n_944), .B2(n_945), .C1(n_952), .C2(n_953), .Y(n_951) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g684 ( .A(n_322), .Y(n_684) );
BUFx2_ASAP7_75t_L g843 ( .A(n_322), .Y(n_843) );
INVx2_ASAP7_75t_SL g955 ( .A(n_322), .Y(n_955) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g651 ( .A(n_325), .Y(n_651) );
BUFx3_ASAP7_75t_L g844 ( .A(n_325), .Y(n_844) );
BUFx3_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
INVx1_ASAP7_75t_L g771 ( .A(n_326), .Y(n_771) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g400 ( .A(n_327), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_328), .A2(n_508), .A3(n_510), .B(n_513), .Y(n_507) );
OAI31xp33_ASAP7_75t_L g841 ( .A1(n_328), .A2(n_842), .A3(n_845), .B(n_850), .Y(n_841) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_329), .A2(n_565), .B(n_578), .Y(n_564) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_330), .B(n_333), .Y(n_329) );
AND2x2_ASAP7_75t_L g652 ( .A(n_330), .B(n_333), .Y(n_652) );
AND2x4_ASAP7_75t_L g691 ( .A(n_330), .B(n_333), .Y(n_691) );
AND2x2_ASAP7_75t_L g797 ( .A(n_330), .B(n_333), .Y(n_797) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g1262 ( .A(n_332), .Y(n_1262) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g384 ( .A(n_335), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g449 ( .A(n_335), .Y(n_449) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_335), .B(n_447), .Y(n_640) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI31xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_360), .A3(n_372), .B(n_377), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_343), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_343), .Y(n_468) );
INVx2_ASAP7_75t_SL g740 ( .A(n_343), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_343), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_343), .B(n_1321), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_343), .A2(n_748), .B1(n_1379), .B2(n_1389), .Y(n_1395) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_344), .Y(n_442) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g502 ( .A(n_346), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_346), .B(n_735), .C(n_737), .Y(n_734) );
INVx3_ASAP7_75t_L g779 ( .A(n_346), .Y(n_779) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g528 ( .A(n_347), .B(n_353), .Y(n_528) );
AND2x2_ASAP7_75t_L g656 ( .A(n_347), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g668 ( .A(n_347), .B(n_369), .Y(n_668) );
BUFx3_ASAP7_75t_L g525 ( .A(n_348), .Y(n_525) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_348), .Y(n_1002) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g658 ( .A(n_349), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_351), .A2(n_525), .B1(n_647), .B2(n_648), .C1(n_660), .C2(n_661), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_351), .A2(n_661), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_351), .A2(n_862), .B1(n_869), .B2(n_870), .Y(n_868) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
OR2x2_ASAP7_75t_L g368 ( .A(n_352), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g499 ( .A(n_352), .B(n_353), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_352), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g531 ( .A(n_352), .Y(n_531) );
AND2x2_ASAP7_75t_L g664 ( .A(n_352), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g1339 ( .A(n_353), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_354), .A2(n_498), .B1(n_500), .B2(n_501), .Y(n_497) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g870 ( .A(n_355), .Y(n_870) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g533 ( .A(n_356), .Y(n_533) );
BUFx3_ASAP7_75t_L g661 ( .A(n_356), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_356), .A2(n_528), .B1(n_975), .B2(n_977), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_357), .B(n_1317), .Y(n_1341) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_362), .Y(n_504) );
AND2x4_ASAP7_75t_L g374 ( .A(n_363), .B(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g506 ( .A(n_368), .Y(n_506) );
INVx1_ASAP7_75t_L g535 ( .A(n_368), .Y(n_535) );
INVx8_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g373 ( .A(n_374), .Y(n_373) );
INVx4_ASAP7_75t_L g492 ( .A(n_374), .Y(n_492) );
INVx3_ASAP7_75t_SL g522 ( .A(n_374), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_374), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_981) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_375), .Y(n_552) );
INVx2_ASAP7_75t_L g724 ( .A(n_375), .Y(n_724) );
BUFx3_ASAP7_75t_L g914 ( .A(n_375), .Y(n_914) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_377), .A2(n_491), .A3(n_493), .B(n_503), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g834 ( .A1(n_377), .A2(n_835), .A3(n_839), .B(n_840), .Y(n_834) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_378), .A2(n_654), .B(n_669), .Y(n_653) );
INVx1_ASAP7_75t_L g741 ( .A(n_378), .Y(n_741) );
BUFx2_ASAP7_75t_L g788 ( .A(n_378), .Y(n_788) );
BUFx2_ASAP7_75t_SL g873 ( .A(n_378), .Y(n_873) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g1308 ( .A(n_380), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1340 ( .A(n_380), .B(n_1341), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_420), .Y(n_381) );
OAI33xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .A3(n_392), .B1(n_401), .B2(n_408), .B3(n_414), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_383), .A2(n_408), .B1(n_579), .B2(n_592), .Y(n_578) );
OAI33xp33_ASAP7_75t_L g601 ( .A1(n_383), .A2(n_602), .A3(n_606), .B1(n_611), .B2(n_617), .B3(n_621), .Y(n_601) );
OAI33xp33_ASAP7_75t_L g766 ( .A1(n_383), .A2(n_621), .A3(n_767), .B1(n_769), .B2(n_772), .B3(n_775), .Y(n_766) );
OAI33xp33_ASAP7_75t_L g823 ( .A1(n_383), .A2(n_408), .A3(n_824), .B1(n_826), .B2(n_829), .B3(n_831), .Y(n_823) );
OAI33xp33_ASAP7_75t_L g892 ( .A1(n_383), .A2(n_893), .A3(n_897), .B1(n_898), .B2(n_901), .B3(n_902), .Y(n_892) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx4f_ASAP7_75t_L g477 ( .A(n_384), .Y(n_477) );
BUFx4f_ASAP7_75t_L g1029 ( .A(n_384), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_387), .A2(n_415), .B1(n_427), .B2(n_431), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_388), .A2(n_415), .B1(n_416), .B2(n_419), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g824 ( .A1(n_388), .A2(n_809), .B1(n_817), .B2(n_825), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_388), .A2(n_810), .B1(n_818), .B2(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_388), .A2(n_1287), .B1(n_1288), .B2(n_1289), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_389), .A2(n_419), .B1(n_435), .B2(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g768 ( .A(n_391), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_397), .B2(n_398), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_393), .A2(n_405), .B1(n_435), .B2(n_440), .Y(n_434) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_395), .A2(n_398), .B1(n_460), .B2(n_474), .Y(n_485) );
OAI22xp33_ASAP7_75t_SL g769 ( .A1(n_395), .A2(n_747), .B1(n_759), .B2(n_770), .Y(n_769) );
INVx5_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g404 ( .A(n_396), .Y(n_404) );
INVx2_ASAP7_75t_SL g487 ( .A(n_396), .Y(n_487) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_396), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_397), .A2(n_407), .B1(n_427), .B2(n_431), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_398), .A2(n_541), .B1(n_548), .B2(n_593), .C(n_595), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_398), .A2(n_581), .B1(n_882), .B2(n_890), .Y(n_897) );
CKINVDCx8_ASAP7_75t_R g398 ( .A(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g615 ( .A(n_399), .Y(n_615) );
INVx3_ASAP7_75t_L g1035 ( .A(n_399), .Y(n_1035) );
INVx1_ASAP7_75t_L g1288 ( .A(n_399), .Y(n_1288) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g610 ( .A(n_400), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_406), .B2(n_407), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_406), .A2(n_462), .B1(n_475), .B2(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_406), .A2(n_812), .B1(n_820), .B2(n_827), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_406), .A2(n_813), .B1(n_822), .B2(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_406), .A2(n_883), .B1(n_891), .B2(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g712 ( .A(n_408), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
INVx2_ASAP7_75t_L g901 ( .A(n_409), .Y(n_901) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g935 ( .A(n_410), .Y(n_935) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g1314 ( .A(n_412), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_412), .B(n_1310), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_416), .A2(n_458), .B1(n_469), .B2(n_479), .Y(n_489) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g833 ( .A(n_418), .Y(n_833) );
INVx1_ASAP7_75t_L g847 ( .A(n_418), .Y(n_847) );
OR2x6_ASAP7_75t_L g1271 ( .A(n_418), .B(n_1272), .Y(n_1271) );
OAI33xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_426), .A3(n_434), .B1(n_443), .B2(n_445), .B3(n_450), .Y(n_420) );
OAI33xp33_ASAP7_75t_L g455 ( .A1(n_421), .A2(n_456), .A3(n_459), .B1(n_463), .B2(n_470), .B3(n_471), .Y(n_455) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_421), .A2(n_445), .A3(n_876), .B1(n_881), .B2(n_884), .B3(n_887), .Y(n_875) );
OAI33xp33_ASAP7_75t_L g1342 ( .A1(n_421), .A2(n_761), .A3(n_1343), .B1(n_1346), .B2(n_1348), .B3(n_1350), .Y(n_1342) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g624 ( .A(n_422), .Y(n_624) );
INVx2_ASAP7_75t_L g716 ( .A(n_422), .Y(n_716) );
INVx4_ASAP7_75t_L g757 ( .A(n_422), .Y(n_757) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g563 ( .A(n_423), .Y(n_563) );
OR2x6_ASAP7_75t_L g621 ( .A(n_423), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_423), .B(n_622), .Y(n_1038) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g695 ( .A(n_424), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_424), .B(n_1317), .Y(n_1335) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_429), .A2(n_431), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g752 ( .A(n_430), .Y(n_752) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_430), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_431), .A2(n_472), .B1(n_474), .B2(n_475), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_431), .A2(n_472), .B1(n_809), .B2(n_810), .Y(n_808) );
INVx6_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx5_ASAP7_75t_L g542 ( .A(n_432), .Y(n_542) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx4_ASAP7_75t_L g627 ( .A(n_433), .Y(n_627) );
INVx2_ASAP7_75t_L g638 ( .A(n_433), .Y(n_638) );
INVx1_ASAP7_75t_L g754 ( .A(n_433), .Y(n_754) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_433), .Y(n_1016) );
INVx2_ASAP7_75t_L g1347 ( .A(n_433), .Y(n_1347) );
INVx1_ASAP7_75t_L g1392 ( .A(n_433), .Y(n_1392) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_435), .A2(n_447), .B1(n_544), .B2(n_545), .C(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_435), .A2(n_544), .B1(n_1300), .B2(n_1349), .Y(n_1348) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g461 ( .A(n_437), .Y(n_461) );
INVx2_ASAP7_75t_L g1020 ( .A(n_437), .Y(n_1020) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g466 ( .A(n_438), .Y(n_466) );
BUFx3_ASAP7_75t_L g629 ( .A(n_438), .Y(n_629) );
INVx1_ASAP7_75t_L g633 ( .A(n_438), .Y(n_633) );
AND2x2_ASAP7_75t_L g558 ( .A(n_439), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_441), .Y(n_444) );
INVx1_ASAP7_75t_L g544 ( .A(n_441), .Y(n_544) );
INVx2_ASAP7_75t_L g1394 ( .A(n_441), .Y(n_1394) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx4f_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
BUFx4f_ASAP7_75t_L g549 ( .A(n_442), .Y(n_549) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_442), .Y(n_630) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_442), .Y(n_634) );
BUFx4f_ASAP7_75t_L g764 ( .A(n_442), .Y(n_764) );
OR2x6_ASAP7_75t_L g1332 ( .A(n_442), .B(n_1333), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g470 ( .A(n_446), .Y(n_470) );
AOI33xp33_ASAP7_75t_L g713 ( .A1(n_446), .A2(n_714), .A3(n_717), .B1(n_720), .B2(n_727), .B3(n_728), .Y(n_713) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_490), .C(n_507), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_476), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_457), .A2(n_467), .B1(n_479), .B2(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g816 ( .A(n_461), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_464), .A2(n_739), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g1344 ( .A(n_465), .Y(n_1344) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_468), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_814) );
OAI33xp33_ASAP7_75t_L g807 ( .A1(n_470), .A2(n_715), .A3(n_808), .B1(n_811), .B2(n_814), .B3(n_819), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_472), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_472), .A2(n_1016), .B1(n_1289), .B2(n_1351), .Y(n_1350) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g626 ( .A(n_473), .Y(n_626) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_473), .Y(n_636) );
INVx2_ASAP7_75t_SL g889 ( .A(n_473), .Y(n_889) );
OAI33xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .A3(n_485), .B1(n_486), .B2(n_488), .B3(n_489), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g895 ( .A(n_481), .Y(n_895) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_481), .A2(n_484), .B1(n_1300), .B2(n_1301), .C(n_1302), .Y(n_1299) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_484), .A2(n_603), .B1(n_753), .B2(n_765), .Y(n_775) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_484), .A2(n_1017), .B1(n_1024), .B2(n_1031), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1387 ( .A1(n_484), .A2(n_603), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_487), .A2(n_615), .B1(n_1021), .B2(n_1027), .Y(n_1036) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_496), .A2(n_632), .B1(n_885), .B2(n_886), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_496), .A2(n_1284), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_498), .A2(n_661), .B1(n_837), .B2(n_838), .Y(n_836) );
BUFx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g738 ( .A(n_499), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g942 ( .A1(n_499), .A2(n_525), .B1(n_661), .B2(n_943), .C1(n_944), .C2(n_945), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_499), .A2(n_661), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g787 ( .A(n_506), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_506), .A2(n_664), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
XOR2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_598), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_562), .B(n_564), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_525), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_528), .A2(n_661), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_530), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g736 ( .A(n_535), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_543), .B(n_547), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_542), .A2(n_877), .B1(n_878), .B2(n_880), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_542), .A2(n_888), .B1(n_890), .B2(n_891), .Y(n_887) );
OAI211xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_549), .B(n_550), .C(n_555), .Y(n_547) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_552), .B(n_1310), .Y(n_1329) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g718 ( .A(n_557), .Y(n_718) );
INVx2_ASAP7_75t_SL g729 ( .A(n_557), .Y(n_729) );
INVx2_ASAP7_75t_L g1000 ( .A(n_557), .Y(n_1000) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_558), .B(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_558), .B(n_1317), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_560), .Y(n_719) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g731 ( .A(n_561), .Y(n_731) );
INVx2_ASAP7_75t_L g1304 ( .A(n_562), .Y(n_1304) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_566), .B(n_574), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_568), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_570), .A2(n_572), .B1(n_645), .B2(n_646), .C1(n_647), .C2(n_648), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_570), .A2(n_572), .B1(n_977), .B2(n_978), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_570), .A2(n_572), .B1(n_1042), .B2(n_1050), .Y(n_1049) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_572), .A2(n_687), .B1(n_1363), .B2(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g851 ( .A(n_575), .Y(n_851) );
INVx2_ASAP7_75t_L g643 ( .A(n_577), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_583), .C(n_588), .Y(n_579) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g699 ( .A(n_584), .Y(n_699) );
BUFx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx8_ASAP7_75t_L g597 ( .A(n_585), .Y(n_597) );
BUFx3_ASAP7_75t_L g929 ( .A(n_585), .Y(n_929) );
NAND2x1p5_ASAP7_75t_L g1260 ( .A(n_585), .B(n_1261), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_585), .B(n_1293), .Y(n_1292) );
BUFx2_ASAP7_75t_L g708 ( .A(n_587), .Y(n_708) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx5_ASAP7_75t_L g706 ( .A(n_590), .Y(n_706) );
BUFx3_ASAP7_75t_L g925 ( .A(n_590), .Y(n_925) );
BUFx12f_ASAP7_75t_L g933 ( .A(n_590), .Y(n_933) );
AND2x4_ASAP7_75t_L g1279 ( .A(n_590), .B(n_1276), .Y(n_1279) );
BUFx3_ASAP7_75t_L g1298 ( .A(n_590), .Y(n_1298) );
INVx1_ASAP7_75t_L g1270 ( .A(n_591), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_593), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g704 ( .A(n_594), .Y(n_704) );
INVx1_ASAP7_75t_L g710 ( .A(n_594), .Y(n_710) );
INVx3_ASAP7_75t_L g900 ( .A(n_594), .Y(n_900) );
OR2x6_ASAP7_75t_SL g1274 ( .A(n_594), .B(n_1275), .Y(n_1274) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_641), .C(n_653), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_623), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_603), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_603), .A2(n_751), .B1(n_763), .B2(n_768), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g1377 ( .A1(n_603), .A2(n_619), .B1(n_1378), .B2(n_1379), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_604), .A2(n_618), .B1(n_626), .B2(n_627), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_605), .A2(n_620), .B1(n_632), .B2(n_634), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_607), .A2(n_614), .B1(n_629), .B2(n_630), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_608), .A2(n_616), .B1(n_636), .B2(n_637), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_609), .A2(n_1384), .B1(n_1385), .B2(n_1386), .Y(n_1383) );
BUFx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g774 ( .A(n_610), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_612), .A2(n_749), .B1(n_760), .B2(n_773), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_612), .A2(n_770), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g1283 ( .A(n_613), .Y(n_1283) );
INVx2_ASAP7_75t_SL g1384 ( .A(n_613), .Y(n_1384) );
INVx1_ASAP7_75t_L g859 ( .A(n_619), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_619), .A2(n_880), .B1(n_886), .B2(n_894), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_619), .A2(n_1015), .B1(n_1023), .B2(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g970 ( .A(n_621), .Y(n_970) );
INVx3_ASAP7_75t_L g1302 ( .A(n_622), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .A3(n_628), .B1(n_631), .B2(n_635), .B3(n_639), .Y(n_623) );
OAI33xp33_ASAP7_75t_L g1390 ( .A1(n_624), .A2(n_639), .A3(n_1391), .B1(n_1393), .B2(n_1395), .B3(n_1396), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_626), .A2(n_637), .B1(n_759), .B2(n_760), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_627), .A2(n_1382), .B1(n_1386), .B2(n_1397), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_629), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_632), .A2(n_739), .B1(n_882), .B2(n_883), .Y(n_881) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g748 ( .A(n_633), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_634), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_634), .A2(n_1020), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1361 ( .A(n_634), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_637), .A2(n_752), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g761 ( .A(n_640), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_640), .B(n_919), .C(n_921), .Y(n_918) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_640), .A2(n_998), .A3(n_999), .B1(n_1001), .B2(n_1003), .B3(n_1004), .Y(n_997) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_649), .B(n_652), .Y(n_641) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_651), .A2(n_940), .B1(n_941), .B2(n_955), .Y(n_954) );
OAI21xp5_ASAP7_75t_L g947 ( .A1(n_652), .A2(n_948), .B(n_950), .Y(n_947) );
OAI31xp33_ASAP7_75t_SL g1046 ( .A1(n_652), .A2(n_1047), .A3(n_1048), .B(n_1051), .Y(n_1046) );
OAI31xp33_ASAP7_75t_L g1367 ( .A1(n_652), .A2(n_1368), .A3(n_1369), .B(n_1374), .Y(n_1367) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_659), .C(n_662), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_655), .B(n_939), .C(n_942), .Y(n_938) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g992 ( .A(n_656), .Y(n_992) );
INVx1_ASAP7_75t_L g991 ( .A(n_657), .Y(n_991) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g726 ( .A(n_658), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_667), .Y(n_662) );
INVx3_ASAP7_75t_L g917 ( .A(n_665), .Y(n_917) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_665), .Y(n_920) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g983 ( .A(n_670), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_905), .B1(n_1054), .B2(n_1055), .Y(n_672) );
INVx1_ASAP7_75t_L g1055 ( .A(n_673), .Y(n_1055) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_802), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_742), .B1(n_800), .B2(n_801), .Y(n_674) );
INVx1_ASAP7_75t_L g801 ( .A(n_675), .Y(n_801) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_677), .B(n_692), .C(n_713), .D(n_732), .Y(n_676) );
AO21x1_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B(n_690), .Y(n_677) );
INVx2_ASAP7_75t_SL g949 ( .A(n_680), .Y(n_949) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx14_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
OAI31xp33_ASAP7_75t_L g855 ( .A1(n_691), .A2(n_856), .A3(n_857), .B(n_864), .Y(n_855) );
AOI33xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .A3(n_702), .B1(n_707), .B2(n_709), .B3(n_712), .Y(n_692) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_694), .B(n_923), .C(n_926), .Y(n_922) );
INVx1_ASAP7_75t_L g963 ( .A(n_694), .Y(n_963) );
BUFx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_699), .A2(n_966), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_700), .B(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g930 ( .A(n_701), .Y(n_930) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g711 ( .A(n_706), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI33xp33_ASAP7_75t_L g1013 ( .A1(n_716), .A2(n_761), .A3(n_1014), .B1(n_1018), .B2(n_1022), .B3(n_1025), .Y(n_1013) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_L g1322 ( .A(n_731), .Y(n_1322) );
AO21x1_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_741), .Y(n_732) );
INVx5_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AO21x1_ASAP7_75t_L g980 ( .A1(n_741), .A2(n_981), .B(n_985), .Y(n_980) );
INVx3_ASAP7_75t_SL g800 ( .A(n_742), .Y(n_800) );
INVx1_ASAP7_75t_L g799 ( .A(n_743), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_776), .C(n_789), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_766), .Y(n_744) );
OAI33xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_750), .A3(n_755), .B1(n_758), .B2(n_761), .B3(n_762), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_748), .A2(n_1381), .B1(n_1385), .B2(n_1394), .Y(n_1393) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_752), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_752), .A2(n_1378), .B1(n_1388), .B2(n_1392), .Y(n_1391) );
BUFx3_ASAP7_75t_L g821 ( .A(n_754), .Y(n_821) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_756), .B(n_911), .C(n_915), .Y(n_910) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_SL g998 ( .A(n_757), .Y(n_998) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI31xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .A3(n_785), .B(n_788), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .C(n_783), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_782), .B(n_795), .Y(n_794) );
OAI31xp33_ASAP7_75t_L g1039 ( .A1(n_788), .A2(n_1040), .A3(n_1044), .B(n_1045), .Y(n_1039) );
OAI31xp33_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_792), .A3(n_796), .B(n_797), .Y(n_789) );
OAI31xp33_ASAP7_75t_SL g971 ( .A1(n_797), .A2(n_972), .A3(n_973), .B(n_979), .Y(n_971) );
OA22x2_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .B1(n_852), .B2(n_853), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_834), .C(n_841), .Y(n_805) );
NOR2xp33_ASAP7_75t_SL g806 ( .A(n_807), .B(n_823), .Y(n_806) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVxp67_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
INVxp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g896 ( .A(n_847), .Y(n_896) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g903 ( .A(n_854), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_866), .C(n_874), .Y(n_854) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
NAND3xp33_ASAP7_75t_SL g973 ( .A(n_860), .B(n_974), .C(n_976), .Y(n_973) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_860), .B(n_1370), .C(n_1372), .Y(n_1369) );
OAI31xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_871), .A3(n_872), .B(n_873), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_873), .A2(n_938), .B(n_946), .Y(n_937) );
OAI31xp33_ASAP7_75t_SL g1359 ( .A1(n_873), .A2(n_1360), .A3(n_1365), .B(n_1366), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_892), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_877), .A2(n_885), .B1(n_894), .B2(n_896), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_878), .A2(n_1287), .B1(n_1301), .B2(n_1347), .Y(n_1346) );
INVx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g1054 ( .A(n_905), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_956), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_937), .C(n_947), .Y(n_908) );
AND4x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_918), .C(n_922), .D(n_931), .Y(n_909) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1005 ( .A(n_917), .Y(n_1005) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_932), .B(n_934), .C(n_936), .Y(n_931) );
BUFx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_1009), .B1(n_1052), .B2(n_1053), .Y(n_956) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_957), .Y(n_1053) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_993), .Y(n_958) );
INVx1_ASAP7_75t_L g995 ( .A(n_960), .Y(n_995) );
AOI21xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_962), .B(n_964), .Y(n_960) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
HB1xp67_ASAP7_75t_L g1373 ( .A(n_967), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_971), .B(n_980), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_978), .B(n_990), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .C(n_992), .Y(n_987) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI31xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .A3(n_996), .B(n_1006), .Y(n_993) );
INVx1_ASAP7_75t_L g1008 ( .A(n_997), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_1009), .Y(n_1052) );
HB1xp67_ASAP7_75t_SL g1009 ( .A(n_1010), .Y(n_1009) );
AND3x1_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1039), .C(n_1046), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1028), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_1019), .A2(n_1026), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
OAI33xp33_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1030), .A3(n_1033), .B1(n_1036), .B2(n_1037), .B3(n_1038), .Y(n_1028) );
OAI33xp33_ASAP7_75t_L g1376 ( .A1(n_1029), .A2(n_1038), .A3(n_1377), .B1(n_1380), .B2(n_1383), .B3(n_1387), .Y(n_1376) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1034), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1064), .B(n_1253), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_1058), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_1059), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_1059), .A2(n_1161), .B1(n_1162), .B2(n_1163), .C(n_1164), .Y(n_1160) );
INVx2_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
AND2x6_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1062), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_1061), .B(n_1073), .Y(n_1072) );
AND2x6_ASAP7_75t_L g1076 ( .A(n_1061), .B(n_1077), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1061), .B(n_1079), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1061), .B(n_1079), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1061), .B(n_1079), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1061), .B(n_1073), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_1062), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1063), .B(n_1074), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1195), .Y(n_1064) );
OAI32xp33_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1125), .A3(n_1157), .B1(n_1170), .B2(n_1185), .Y(n_1065) );
OAI311xp33_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1090), .A3(n_1095), .B1(n_1099), .C1(n_1118), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1080), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1068), .B(n_1180), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_1069), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1069), .B(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1069), .B(n_1117), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1069), .B(n_1152), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1069), .B(n_1134), .Y(n_1207) );
NOR2xp33_ASAP7_75t_L g1236 ( .A(n_1069), .B(n_1148), .Y(n_1236) );
INVx4_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1070), .B(n_1103), .Y(n_1102) );
INVx4_ASAP7_75t_L g1122 ( .A(n_1070), .Y(n_1122) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1070), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1070), .B(n_1136), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1070), .B(n_1128), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1070), .B(n_1124), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1070), .A2(n_1122), .B1(n_1190), .B2(n_1191), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1212 ( .A(n_1070), .B(n_1129), .Y(n_1212) );
NAND2xp5_ASAP7_75t_SL g1221 ( .A(n_1070), .B(n_1124), .Y(n_1221) );
AND2x4_ASAP7_75t_SL g1070 ( .A(n_1071), .B(n_1075), .Y(n_1070) );
AOI222xp33_ASAP7_75t_L g1176 ( .A1(n_1080), .A2(n_1177), .B1(n_1178), .B2(n_1181), .C1(n_1182), .C2(n_1183), .Y(n_1176) );
O2A1O1Ixp33_ASAP7_75t_SL g1215 ( .A1(n_1080), .A2(n_1212), .B(n_1216), .C(n_1222), .Y(n_1215) );
O2A1O1Ixp33_ASAP7_75t_L g1237 ( .A1(n_1080), .A2(n_1238), .B(n_1239), .C(n_1240), .Y(n_1237) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_1081), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1081), .B(n_1116), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1086), .Y(n_1081) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1082), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1085), .Y(n_1082) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1086), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1086), .B(n_1130), .Y(n_1142) );
NOR2xp33_ASAP7_75t_L g1242 ( .A(n_1086), .B(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_1087), .B(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1087), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1090), .B(n_1146), .Y(n_1145) );
OAI211xp5_ASAP7_75t_L g1196 ( .A1(n_1090), .A2(n_1197), .B(n_1205), .C(n_1215), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1090), .B(n_1129), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1090), .B(n_1203), .Y(n_1247) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx3_ASAP7_75t_L g1116 ( .A(n_1091), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1091), .B(n_1130), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1091), .B(n_1177), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1091), .B(n_1130), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1095), .B(n_1104), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1134 ( .A(n_1095), .B(n_1123), .Y(n_1134) );
OAI21xp33_ASAP7_75t_L g1150 ( .A1(n_1095), .A2(n_1151), .B(n_1152), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1095), .B(n_1124), .Y(n_1171) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_1096), .B(n_1104), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1096), .B(n_1104), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1096), .B(n_1154), .Y(n_1153) );
NAND2x1p5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1098), .Y(n_1096) );
OAI21xp5_ASAP7_75t_SL g1099 ( .A1(n_1100), .A2(n_1107), .B(n_1114), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
NAND3xp33_ASAP7_75t_SL g1234 ( .A(n_1101), .B(n_1230), .C(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1102), .B(n_1109), .Y(n_1229) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1103), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1103), .B(n_1188), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1103), .B(n_1123), .Y(n_1217) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1104), .Y(n_1149) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1104), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1104), .B(n_1124), .Y(n_1180) );
OAI32xp33_ASAP7_75t_L g1245 ( .A1(n_1104), .A2(n_1133), .A3(n_1179), .B1(n_1184), .B2(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1106), .Y(n_1104) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1108), .B(n_1172), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1112), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1109), .B(n_1153), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1109), .B(n_1128), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1110), .B(n_1111), .Y(n_1124) );
NOR2x1_ASAP7_75t_L g1121 ( .A(n_1112), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1113), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1113), .B(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
CKINVDCx14_ASAP7_75t_R g1138 ( .A(n_1116), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1116), .B(n_1141), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1116), .B(n_1130), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1116), .B(n_1142), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1116), .B(n_1137), .Y(n_1250) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1117), .Y(n_1119) );
O2A1O1Ixp33_ASAP7_75t_L g1185 ( .A1(n_1117), .A2(n_1186), .B(n_1189), .C(n_1193), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1120), .Y(n_1118) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_1120), .A2(n_1138), .B(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1123), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1122), .B(n_1177), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_1122), .Y(n_1203) );
O2A1O1Ixp33_ASAP7_75t_SL g1228 ( .A1(n_1122), .A2(n_1171), .B(n_1229), .C(n_1230), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1122), .B(n_1160), .Y(n_1252) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_1123), .A2(n_1126), .B1(n_1138), .B2(n_1139), .C(n_1143), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1123), .B(n_1128), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1123), .B(n_1153), .Y(n_1192) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1124), .B(n_1149), .Y(n_1148) );
AOI22xp5_ASAP7_75t_SL g1126 ( .A1(n_1127), .A2(n_1129), .B1(n_1131), .B2(n_1135), .Y(n_1126) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1127), .Y(n_1214) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1128), .Y(n_1200) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1129), .Y(n_1155) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1130), .Y(n_1169) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1130), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1130), .B(n_1137), .Y(n_1204) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND2xp5_ASAP7_75t_SL g1173 ( .A(n_1136), .B(n_1174), .Y(n_1173) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g1208 ( .A(n_1137), .B(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_1140), .A2(n_1182), .B1(n_1190), .B2(n_1249), .Y(n_1248) );
O2A1O1Ixp33_ASAP7_75t_L g1244 ( .A1(n_1141), .A2(n_1190), .B(n_1207), .C(n_1245), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_1142), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1147), .B1(n_1150), .B2(n_1155), .C(n_1156), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1146), .Y(n_1224) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
AOI22xp5_ASAP7_75t_L g1197 ( .A1(n_1149), .A2(n_1198), .B1(n_1201), .B2(n_1202), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1153), .B(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1155), .B(n_1247), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1165), .Y(n_1156) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1157), .Y(n_1225) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1168), .C(n_1169), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1168), .B(n_1220), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B(n_1173), .C(n_1176), .Y(n_1170) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1180), .Y(n_1182) );
CKINVDCx14_ASAP7_75t_R g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AOI21xp5_ASAP7_75t_L g1222 ( .A1(n_1192), .A2(n_1223), .B(n_1224), .Y(n_1222) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AOI21xp5_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1225), .B(n_1226), .Y(n_1195) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1204), .Y(n_1251) );
AOI211xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .B(n_1208), .C(n_1210), .Y(n_1205) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1206), .Y(n_1213) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1209), .Y(n_1238) );
AOI21xp33_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1213), .B(n_1214), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
NAND5xp2_ASAP7_75t_SL g1226 ( .A(n_1227), .B(n_1237), .C(n_1241), .D(n_1244), .E(n_1248), .Y(n_1226) );
OAI21xp5_ASAP7_75t_SL g1227 ( .A1(n_1228), .A2(n_1232), .B(n_1234), .Y(n_1227) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVxp67_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1239), .Y(n_1243) );
AOI21xp33_ASAP7_75t_L g1249 ( .A1(n_1250), .A2(n_1251), .B(n_1252), .Y(n_1249) );
AOI211x1_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1303), .B(n_1305), .C(n_1330), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1280), .Y(n_1256) );
AOI211xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1259), .B(n_1263), .C(n_1273), .Y(n_1257) );
AOI222xp33_ASAP7_75t_L g1311 ( .A1(n_1258), .A2(n_1312), .B1(n_1318), .B2(n_1319), .C1(n_1323), .C2(n_1325), .Y(n_1311) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AND2x6_ASAP7_75t_L g1265 ( .A(n_1261), .B(n_1266), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1261), .B(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1261), .Y(n_1272) );
INVx4_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx3_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1277), .Y(n_1293) );
INVx3_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NOR3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1290), .C(n_1296), .Y(n_1280) );
OAI21xp33_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1284), .B(n_1285), .Y(n_1282) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx3_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
AND2x4_ASAP7_75t_L g1328 ( .A(n_1308), .B(n_1329), .Y(n_1328) );
AND2x4_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
AND2x4_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1322), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
OR3x1_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1336), .C(n_1342), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
NAND2x2_ASAP7_75t_L g1337 ( .A(n_1334), .B(n_1338), .Y(n_1337) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx2_ASAP7_75t_SL g1338 ( .A(n_1339), .Y(n_1338) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g1355 ( .A(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
NAND3xp33_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1367), .C(n_1375), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1364), .B(n_1373), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1390), .Y(n_1375) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
HB1xp67_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
OAI21xp5_ASAP7_75t_L g1403 ( .A1(n_1404), .A2(n_1405), .B(n_1406), .Y(n_1403) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
endmodule