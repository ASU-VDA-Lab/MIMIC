module fake_netlist_6_1356_n_1803 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1803);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1803;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_86),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_61),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_19),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_96),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_139),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_10),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_31),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g193 ( 
.A(n_126),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_25),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_14),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_36),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_92),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_45),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_69),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_19),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_70),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_46),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_57),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_33),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_31),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_34),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_78),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_50),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_66),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_60),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_122),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_167),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_102),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_55),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_27),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_110),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_174),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_145),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_83),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_25),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_95),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_87),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_28),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_142),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_154),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_3),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_119),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_108),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_114),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_54),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_81),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_125),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_109),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_85),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_164),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_62),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_150),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_1),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_162),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_79),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_115),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_88),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_84),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_91),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_16),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_77),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_56),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_73),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_141),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_107),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_9),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_48),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_44),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_40),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_40),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_11),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_130),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_67),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_166),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_64),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_93),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_161),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_105),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_123),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_39),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_89),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_15),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_16),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_100),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_144),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_137),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_101),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_33),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_99),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_152),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_42),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_169),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_75),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_20),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_7),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_120),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_165),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_53),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_37),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_5),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_37),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_47),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_103),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_211),
.B(n_0),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_178),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_229),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_178),
.Y(n_353)
);

BUFx6f_ASAP7_75t_SL g354 ( 
.A(n_342),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_270),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_217),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_190),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_195),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_190),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_195),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_188),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_197),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_189),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_191),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_245),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_198),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_264),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_272),
.B(n_4),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_209),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_197),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_184),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_286),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_212),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_225),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_198),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_199),
.B(n_5),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_203),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_212),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_197),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_226),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_220),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_204),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_236),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_255),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_208),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_271),
.Y(n_398)
);

BUFx6f_ASAP7_75t_SL g399 ( 
.A(n_342),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_283),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_210),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_235),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_215),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_220),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_305),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_310),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_286),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_242),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_298),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_272),
.B(n_8),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_219),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_199),
.B(n_10),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_242),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_227),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_235),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_247),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_248),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_249),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_272),
.B(n_12),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_179),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_248),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_254),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_257),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_181),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_260),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_183),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_265),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_282),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_360),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_292),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_362),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_360),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_292),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_349),
.B(n_192),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_366),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_402),
.B(n_287),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_349),
.A2(n_296),
.B(n_244),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_194),
.Y(n_459)
);

BUFx2_ASAP7_75t_SL g460 ( 
.A(n_375),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_391),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_418),
.B(n_192),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_368),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_244),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_281),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_281),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_321),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_352),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_352),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_361),
.B(n_321),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_369),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_369),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_364),
.B(n_296),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_L g477 ( 
.A(n_350),
.B(n_223),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_351),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_373),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_415),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_416),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_387),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_353),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_355),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_379),
.B(n_194),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_423),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_396),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_356),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_394),
.B(n_372),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_370),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_401),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_357),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_466),
.B(n_273),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_462),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_463),
.B(n_273),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_403),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_463),
.B(n_273),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_223),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_371),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_463),
.B(n_273),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_463),
.B(n_291),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_489),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_378),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_490),
.B(n_414),
.Y(n_532)
);

BUFx8_ASAP7_75t_SL g533 ( 
.A(n_478),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_498),
.A2(n_196),
.B1(n_206),
.B2(n_213),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_512),
.A2(n_425),
.B1(n_435),
.B2(n_432),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_498),
.A2(n_291),
.B1(n_318),
.B2(n_239),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_414),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_460),
.B(n_421),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_441),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_509),
.B(n_421),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_509),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_512),
.A2(n_436),
.B1(n_435),
.B2(n_432),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_466),
.B(n_291),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_509),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_466),
.A2(n_291),
.B1(n_318),
.B2(n_224),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_500),
.B(n_371),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_201),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_443),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g560 ( 
.A(n_466),
.B(n_291),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_500),
.B(n_385),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_501),
.B(n_500),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_453),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_425),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_456),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_501),
.B(n_318),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_470),
.B(n_409),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_461),
.B(n_258),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_385),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_503),
.B(n_430),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_506),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_466),
.A2(n_318),
.B1(n_230),
.B2(n_237),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_438),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_460),
.B(n_430),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_469),
.B(n_318),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_470),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_501),
.B(n_436),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_454),
.B(n_221),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_438),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_471),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_504),
.B(n_433),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_504),
.B(n_411),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_506),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_454),
.B(n_243),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_438),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_469),
.B(n_302),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_444),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_438),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_354),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_464),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_496),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_482),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_506),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_478),
.A2(n_196),
.B1(n_206),
.B2(n_213),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_469),
.B(n_202),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_438),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_469),
.A2(n_323),
.B1(n_205),
.B2(n_276),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_513),
.B(n_354),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_444),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_511),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_354),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_399),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_458),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_457),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_470),
.B(n_193),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_469),
.A2(n_455),
.B1(n_448),
.B2(n_477),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_501),
.B(n_269),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_R g625 ( 
.A(n_437),
.B(n_284),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_488),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_501),
.B(n_289),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_506),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_452),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_458),
.A2(n_258),
.B1(n_263),
.B2(n_275),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_496),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_259),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_501),
.B(n_297),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_455),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_442),
.B(n_175),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_488),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_497),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_501),
.A2(n_324),
.B1(n_267),
.B2(n_345),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_508),
.B(n_285),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_448),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_452),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_488),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_465),
.B(n_473),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_444),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_499),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_445),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_485),
.A2(n_278),
.B1(n_275),
.B2(n_263),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_485),
.B(n_298),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_499),
.B(n_399),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_496),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_444),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_442),
.B(n_176),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_465),
.B(n_473),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

INVx4_ASAP7_75t_SL g660 ( 
.A(n_496),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_496),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_499),
.B(n_300),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_486),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_508),
.B(n_307),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_562),
.B(n_499),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_562),
.B(n_499),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_525),
.B(n_502),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_520),
.A2(n_477),
.B1(n_448),
.B2(n_465),
.Y(n_669)
);

AO22x1_ASAP7_75t_L g670 ( 
.A1(n_592),
.A2(n_502),
.B1(n_507),
.B2(n_445),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_502),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_643),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_665),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_593),
.A2(n_555),
.B1(n_561),
.B2(n_547),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_555),
.B(n_502),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_561),
.B(n_502),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_643),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_520),
.A2(n_448),
.B1(n_468),
.B2(n_473),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_642),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_560),
.B(n_447),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_523),
.A2(n_447),
.B(n_448),
.C(n_468),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_544),
.B(n_450),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_523),
.A2(n_468),
.B(n_510),
.C(n_508),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_535),
.B(n_507),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_515),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_524),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_519),
.B(n_450),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_551),
.B(n_474),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_518),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_521),
.B(n_508),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_587),
.B(n_595),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_519),
.B(n_474),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_648),
.B(n_476),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_579),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_560),
.B(n_475),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_529),
.Y(n_698)
);

O2A1O1Ixp5_ASAP7_75t_L g699 ( 
.A1(n_527),
.A2(n_452),
.B(n_446),
.C(n_449),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_537),
.B(n_510),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_524),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_648),
.A2(n_475),
.B1(n_320),
.B2(n_278),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_623),
.A2(n_320),
.B1(n_182),
.B2(n_315),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_575),
.B(n_472),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_486),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_527),
.A2(n_510),
.B(n_476),
.C(n_493),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_575),
.B(n_472),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_594),
.B(n_486),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_528),
.A2(n_476),
.B1(n_324),
.B2(n_267),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_579),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_604),
.B(n_658),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_658),
.B(n_486),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_543),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_574),
.B(n_510),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_532),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_556),
.B(n_486),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_486),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_638),
.B(n_486),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_574),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_657),
.B(n_654),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_573),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_550),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_650),
.B(n_467),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_528),
.A2(n_338),
.B1(n_341),
.B2(n_348),
.Y(n_726)
);

BUFx8_ASAP7_75t_L g727 ( 
.A(n_585),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_554),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_650),
.B(n_467),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_654),
.B(n_486),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_597),
.B(n_487),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_631),
.B(n_262),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_577),
.A2(n_327),
.B1(n_424),
.B2(n_388),
.Y(n_734)
);

AO22x1_ASAP7_75t_L g735 ( 
.A1(n_542),
.A2(n_319),
.B1(n_309),
.B2(n_308),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_631),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_564),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_539),
.B(n_262),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_605),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_605),
.B(n_467),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_612),
.B(n_467),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_567),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_SL g743 ( 
.A1(n_606),
.A2(n_404),
.B1(n_363),
.B2(n_428),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_653),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_540),
.B(n_487),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_552),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_612),
.B(n_467),
.Y(n_747)
);

AO22x1_ASAP7_75t_L g748 ( 
.A1(n_600),
.A2(n_294),
.B1(n_336),
.B2(n_290),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_565),
.B(n_280),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_SL g750 ( 
.A(n_566),
.B(n_365),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_583),
.B(n_280),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_586),
.B(n_177),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_540),
.B(n_487),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_620),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_626),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_530),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_626),
.B(n_487),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_536),
.A2(n_253),
.B1(n_307),
.B2(n_299),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_545),
.B(n_487),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_637),
.B(n_663),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_637),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_530),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_625),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_610),
.A2(n_481),
.B1(n_493),
.B2(n_492),
.C(n_480),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_663),
.B(n_487),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_598),
.B(n_487),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_586),
.A2(n_376),
.B1(n_382),
.B2(n_392),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_619),
.B(n_399),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_621),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_617),
.B(n_618),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_551),
.B(n_467),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_536),
.B(n_467),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_641),
.B(n_304),
.C(n_331),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_617),
.B(n_467),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_559),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_628),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_SL g778 ( 
.A(n_616),
.B(n_410),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_618),
.B(n_480),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_577),
.B(n_480),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_610),
.A2(n_420),
.B1(n_293),
.B2(n_288),
.Y(n_781)
);

NAND2x1_ASAP7_75t_L g782 ( 
.A(n_569),
.B(n_452),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_628),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_629),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_624),
.A2(n_228),
.B1(n_233),
.B2(n_232),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_635),
.B(n_600),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_625),
.B(n_641),
.C(n_613),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_578),
.B(n_580),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_582),
.B(n_480),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_629),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_603),
.B(n_481),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_481),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_R g793 ( 
.A(n_651),
.B(n_514),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_635),
.B(n_322),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_614),
.Y(n_795)
);

INVxp33_ASAP7_75t_SL g796 ( 
.A(n_640),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_571),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_533),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_624),
.A2(n_253),
.B1(n_307),
.B2(n_325),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_613),
.B(n_185),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_627),
.B(n_481),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_630),
.A2(n_253),
.B1(n_332),
.B2(n_492),
.Y(n_802)
);

NOR3x1_ASAP7_75t_L g803 ( 
.A(n_534),
.B(n_514),
.C(n_497),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_639),
.B(n_644),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_516),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_548),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_630),
.A2(n_207),
.B1(n_343),
.B2(n_337),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_516),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_646),
.B(n_253),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_538),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_647),
.B(n_636),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_635),
.B(n_622),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_636),
.A2(n_253),
.B1(n_492),
.B2(n_483),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_530),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_541),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_570),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_570),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_558),
.B(n_483),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_541),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_608),
.A2(n_253),
.B1(n_492),
.B2(n_483),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_622),
.A2(n_187),
.B1(n_334),
.B2(n_333),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_549),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_568),
.B(n_493),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_534),
.B(n_493),
.C(n_274),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_186),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_568),
.B(n_253),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_656),
.B(n_452),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_718),
.A2(n_655),
.B(n_662),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_692),
.A2(n_676),
.B1(n_771),
.B2(n_673),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_695),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_739),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_692),
.B(n_608),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_715),
.A2(n_710),
.B(n_720),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_757),
.A2(n_655),
.B(n_662),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_695),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_674),
.B(n_563),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_739),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_760),
.A2(n_664),
.B(n_645),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_808),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_732),
.A2(n_741),
.B(n_740),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_805),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_739),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_691),
.B(n_651),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_676),
.A2(n_608),
.B1(n_652),
.B2(n_633),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_810),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_774),
.A2(n_608),
.B1(n_607),
.B2(n_588),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_740),
.A2(n_661),
.B(n_602),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_741),
.A2(n_661),
.B(n_602),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_739),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_668),
.A2(n_675),
.B1(n_671),
.B2(n_696),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_683),
.A2(n_632),
.B(n_645),
.C(n_572),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_715),
.A2(n_632),
.B(n_572),
.C(n_588),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_704),
.A2(n_607),
.B(n_591),
.C(n_570),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_699),
.A2(n_747),
.B(n_681),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_711),
.A2(n_591),
.B1(n_649),
.B2(n_590),
.Y(n_856)
);

INVx11_ASAP7_75t_L g857 ( 
.A(n_727),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_771),
.B(n_608),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_761),
.A2(n_569),
.B1(n_590),
.B2(n_599),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_755),
.A2(n_609),
.B(n_599),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_716),
.B(n_563),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_763),
.B(n_601),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_719),
.A2(n_589),
.B(n_596),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_727),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_701),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_796),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_713),
.A2(n_581),
.B(n_596),
.Y(n_867)
);

BUFx4f_ASAP7_75t_L g868 ( 
.A(n_756),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_744),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_755),
.A2(n_581),
.B(n_596),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_731),
.A2(n_581),
.B(n_596),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_733),
.B(n_609),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_679),
.B(n_601),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_705),
.B(n_708),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_787),
.A2(n_214),
.B(n_216),
.C(n_200),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_806),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_722),
.B(n_611),
.Y(n_878)
);

AO22x1_ASAP7_75t_L g879 ( 
.A1(n_803),
.A2(n_517),
.B1(n_546),
.B2(n_584),
.Y(n_879)
);

BUFx4f_ASAP7_75t_L g880 ( 
.A(n_825),
.Y(n_880)
);

BUFx12f_ASAP7_75t_L g881 ( 
.A(n_798),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_806),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_680),
.A2(n_584),
.B(n_546),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_762),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_733),
.B(n_517),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_815),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_666),
.A2(n_548),
.B(n_659),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_738),
.B(n_517),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_819),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_738),
.B(n_517),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_667),
.A2(n_548),
.B(n_659),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_517),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_749),
.B(n_546),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_795),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_751),
.B(n_611),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_759),
.A2(n_546),
.B1(n_584),
.B2(n_218),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_725),
.A2(n_548),
.B(n_659),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_751),
.B(n_546),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_725),
.A2(n_659),
.B(n_634),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_822),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_730),
.A2(n_634),
.B(n_557),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_712),
.B(n_697),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_686),
.B(n_660),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_730),
.A2(n_634),
.B(n_557),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_746),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_806),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_678),
.B(n_584),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_759),
.A2(n_584),
.B1(n_222),
.B2(n_301),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_678),
.B(n_634),
.Y(n_909)
);

O2A1O1Ixp5_ASAP7_75t_L g910 ( 
.A1(n_779),
.A2(n_449),
.B(n_446),
.C(n_440),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_707),
.B(n_295),
.C(n_234),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_814),
.Y(n_912)
);

BUFx2_ASAP7_75t_SL g913 ( 
.A(n_684),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_682),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_745),
.A2(n_753),
.B(n_766),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_726),
.A2(n_721),
.B1(n_669),
.B2(n_697),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_688),
.A2(n_726),
.B(n_786),
.C(n_689),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_786),
.A2(n_329),
.B(n_238),
.C(n_231),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_781),
.B(n_316),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_685),
.A2(n_240),
.B(n_241),
.C(n_246),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_702),
.B(n_690),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_669),
.A2(n_311),
.B1(n_251),
.B2(n_252),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_818),
.A2(n_557),
.B(n_449),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_687),
.A2(n_446),
.B(n_440),
.C(n_261),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_793),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_734),
.B(n_250),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_780),
.A2(n_440),
.B(n_312),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_775),
.A2(n_660),
.B(n_326),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_824),
.A2(n_342),
.B1(n_303),
.B2(n_314),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_776),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_693),
.B(n_313),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_703),
.B(n_670),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_767),
.B(n_256),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_698),
.B(n_279),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_710),
.A2(n_277),
.B1(n_268),
.B2(n_660),
.Y(n_935)
);

AOI33xp33_ASAP7_75t_L g936 ( 
.A1(n_743),
.A2(n_12),
.A3(n_13),
.B1(n_20),
.B2(n_21),
.B3(n_23),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_706),
.A2(n_68),
.B(n_171),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_SL g938 ( 
.A(n_778),
.B(n_21),
.Y(n_938)
);

NOR2x1_ASAP7_75t_L g939 ( 
.A(n_687),
.B(n_65),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_709),
.A2(n_74),
.B(n_157),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_700),
.B(n_23),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_714),
.B(n_26),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_811),
.A2(n_80),
.B(n_156),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_672),
.A2(n_63),
.B1(n_149),
.B2(n_140),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_788),
.A2(n_52),
.B(n_134),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_723),
.B(n_49),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_804),
.B(n_772),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_728),
.A2(n_27),
.B(n_30),
.C(n_34),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_717),
.A2(n_765),
.B(n_827),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_729),
.B(n_742),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_694),
.B(n_90),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_817),
.B(n_30),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_677),
.A2(n_694),
.B1(n_737),
.B2(n_820),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_750),
.B(n_35),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_797),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_752),
.A2(n_809),
.B(n_758),
.C(n_826),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_782),
.A2(n_98),
.B(n_132),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_825),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_816),
.B(n_58),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_724),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_772),
.A2(n_172),
.B(n_127),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_754),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_768),
.B(n_35),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_769),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_820),
.A2(n_121),
.B1(n_116),
.B2(n_113),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_789),
.A2(n_112),
.B(n_41),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_791),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_770),
.B(n_38),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_794),
.B(n_41),
.Y(n_969)
);

NOR2x1p5_ASAP7_75t_SL g970 ( 
.A(n_777),
.B(n_42),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_823),
.A2(n_44),
.B(n_47),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_792),
.A2(n_48),
.B(n_801),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_758),
.A2(n_799),
.B1(n_812),
.B2(n_802),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_768),
.B(n_794),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_809),
.A2(n_783),
.B(n_784),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_812),
.A2(n_799),
.B(n_790),
.C(n_802),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_826),
.A2(n_764),
.B(n_800),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_821),
.A2(n_785),
.B(n_807),
.C(n_748),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_813),
.A2(n_735),
.B(n_793),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_813),
.B(n_674),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_676),
.A2(n_668),
.B1(n_675),
.B2(n_671),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_695),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_736),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_SL g987 ( 
.A(n_739),
.B(n_755),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_736),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_692),
.A2(n_676),
.B1(n_771),
.B2(n_673),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_676),
.A2(n_668),
.B1(n_675),
.B2(n_671),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_718),
.A2(n_760),
.B(n_699),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_691),
.B(n_544),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_704),
.A2(n_720),
.B(n_676),
.C(n_688),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_740),
.A2(n_747),
.B(n_741),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_740),
.A2(n_747),
.B(n_741),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_720),
.B(n_692),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_999)
);

AOI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_692),
.A2(n_676),
.B(n_715),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_692),
.A2(n_676),
.B(n_683),
.C(n_715),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_692),
.B(n_676),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_692),
.A2(n_676),
.B(n_683),
.C(n_715),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_692),
.B(n_676),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_718),
.A2(n_519),
.B(n_757),
.Y(n_1006)
);

AO31x2_ASAP7_75t_L g1007 ( 
.A1(n_982),
.A2(n_990),
.A3(n_1004),
.B(n_1001),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_864),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_981),
.A2(n_985),
.B(n_984),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_887),
.A2(n_863),
.B(n_834),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_866),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_876),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_828),
.A2(n_910),
.B(n_949),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_962),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_899),
.A2(n_897),
.B(n_867),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_991),
.A2(n_999),
.B(n_995),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_964),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_993),
.B(n_865),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_SL g1021 ( 
.A1(n_971),
.A2(n_997),
.B(n_996),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_865),
.B(n_998),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_1003),
.A2(n_1006),
.B(n_882),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_841),
.A2(n_992),
.B(n_855),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_1000),
.A2(n_994),
.B(n_833),
.C(n_926),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_902),
.A2(n_872),
.B(n_851),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_882),
.A2(n_832),
.B(n_977),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_831),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_947),
.A2(n_916),
.B(n_980),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_976),
.A2(n_973),
.B(n_853),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_882),
.A2(n_858),
.B(n_860),
.Y(n_1031)
);

BUFx2_ASAP7_75t_SL g1032 ( 
.A(n_866),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_848),
.A2(n_849),
.B(n_975),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_928),
.A2(n_890),
.B(n_888),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_889),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_869),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_874),
.A2(n_969),
.B(n_845),
.C(n_854),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_852),
.A2(n_927),
.B(n_989),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_829),
.B(n_967),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_860),
.A2(n_909),
.B(n_870),
.Y(n_1040)
);

AOI221x1_ASAP7_75t_L g1041 ( 
.A1(n_971),
.A2(n_932),
.B1(n_911),
.B2(n_972),
.C(n_917),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_892),
.A2(n_898),
.B(n_893),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_831),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_839),
.A2(n_907),
.B(n_885),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_927),
.A2(n_951),
.B(n_979),
.C(n_918),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_956),
.A2(n_933),
.B(n_919),
.C(n_954),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_911),
.A2(n_953),
.B(n_883),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_SL g1048 ( 
.A1(n_974),
.A2(n_963),
.B(n_844),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_873),
.B(n_836),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_876),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_950),
.B(n_840),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_846),
.B(n_886),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_986),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_883),
.A2(n_847),
.B(n_859),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_938),
.A2(n_914),
.B1(n_929),
.B2(n_978),
.C(n_837),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_923),
.A2(n_904),
.B(n_901),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_856),
.A2(n_957),
.B(n_961),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_843),
.A2(n_924),
.B(n_894),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_881),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_941),
.A2(n_942),
.B(n_946),
.C(n_983),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_900),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_905),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_875),
.A2(n_896),
.B(n_939),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_838),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_968),
.A2(n_948),
.A3(n_920),
.B(n_966),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_838),
.Y(n_1066)
);

OA22x2_ASAP7_75t_L g1067 ( 
.A1(n_914),
.A2(n_952),
.B1(n_884),
.B2(n_912),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_930),
.A2(n_955),
.B(n_943),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_843),
.A2(n_850),
.B(n_876),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_842),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_895),
.B(n_938),
.C(n_931),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_877),
.Y(n_1072)
);

OA22x2_ASAP7_75t_L g1073 ( 
.A1(n_952),
.A2(n_988),
.B1(n_913),
.B2(n_921),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_861),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_945),
.A2(n_940),
.B(n_937),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_878),
.B(n_925),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_830),
.B(n_835),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_921),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_946),
.A2(n_880),
.B1(n_850),
.B2(n_965),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_959),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_850),
.A2(n_877),
.B(n_906),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_934),
.A2(n_944),
.B(n_908),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_935),
.A2(n_922),
.B1(n_959),
.B2(n_960),
.C(n_970),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_987),
.B(n_958),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_960),
.B(n_903),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_862),
.B(n_903),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_880),
.A2(n_936),
.B(n_878),
.C(n_868),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_877),
.A2(n_906),
.B(n_879),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_906),
.A2(n_868),
.B(n_958),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_958),
.B(n_952),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_857),
.A2(n_519),
.B(n_755),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_969),
.B(n_573),
.C(n_445),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_981),
.A2(n_519),
.B(n_755),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_981),
.A2(n_1003),
.B(n_999),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_974),
.A2(n_692),
.B1(n_998),
.B2(n_874),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_829),
.B(n_989),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_982),
.A2(n_990),
.A3(n_1004),
.B(n_1001),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_840),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_1000),
.A2(n_771),
.B(n_676),
.C(n_650),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_881),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_981),
.A2(n_519),
.B(n_755),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_927),
.A2(n_855),
.B(n_839),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_866),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_1000),
.A2(n_771),
.B(n_676),
.C(n_650),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_840),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_981),
.A2(n_985),
.B(n_984),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_962),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_881),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_1000),
.A2(n_771),
.B(n_676),
.C(n_650),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_981),
.A2(n_985),
.B(n_984),
.Y(n_1118)
);

AOI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_994),
.A2(n_833),
.B(n_926),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_L g1120 ( 
.A1(n_981),
.A2(n_1003),
.B(n_999),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1000),
.A2(n_994),
.B(n_833),
.C(n_1002),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1000),
.A2(n_994),
.B(n_833),
.C(n_1002),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_998),
.B(n_720),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_962),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_829),
.B(n_989),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_981),
.A2(n_985),
.B(n_984),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_1000),
.A2(n_771),
.B(n_676),
.C(n_650),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_866),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_981),
.A2(n_519),
.B(n_755),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_865),
.B(n_544),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1002),
.A2(n_1005),
.B1(n_1001),
.B2(n_1004),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_993),
.B(n_691),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_969),
.B(n_998),
.C(n_787),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1000),
.A2(n_994),
.B(n_833),
.C(n_1002),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_876),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_881),
.B(n_744),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_831),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1000),
.A2(n_994),
.B(n_833),
.C(n_1002),
.Y(n_1140)
);

OA22x2_ASAP7_75t_L g1141 ( 
.A1(n_845),
.A2(n_633),
.B1(n_652),
.B2(n_606),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_981),
.A2(n_519),
.B(n_755),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_SL g1143 ( 
.A1(n_971),
.A2(n_997),
.B(n_996),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_981),
.A2(n_985),
.B(n_984),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_881),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_SL g1146 ( 
.A1(n_858),
.A2(n_832),
.B(n_885),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_833),
.A2(n_641),
.B1(n_534),
.B2(n_710),
.C(n_734),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_913),
.B(n_881),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_SL g1150 ( 
.A1(n_971),
.A2(n_997),
.B(n_996),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_974),
.A2(n_692),
.B1(n_998),
.B2(n_874),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_998),
.B(n_720),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_871),
.A2(n_915),
.B(n_891),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_939),
.B(n_739),
.Y(n_1154)
);

BUFx5_ASAP7_75t_L g1155 ( 
.A(n_903),
.Y(n_1155)
);

AO21x1_ASAP7_75t_L g1156 ( 
.A1(n_1000),
.A2(n_916),
.B(n_994),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1002),
.B(n_1005),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_981),
.A2(n_519),
.B(n_755),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_SL g1159 ( 
.A1(n_971),
.A2(n_997),
.B(n_996),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1061),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1092),
.A2(n_1106),
.B1(n_1157),
.B2(n_1095),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1130),
.B(n_1020),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1030),
.A2(n_1047),
.B(n_1038),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1022),
.B(n_1132),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1080),
.B(n_1078),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1062),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_L g1167 ( 
.A(n_1046),
.B(n_1155),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1009),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1102),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1028),
.Y(n_1170)
);

AOI222xp33_ASAP7_75t_L g1171 ( 
.A1(n_1147),
.A2(n_1125),
.B1(n_1099),
.B2(n_1133),
.C1(n_1093),
.C2(n_1152),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1112),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1098),
.B(n_1151),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1123),
.B(n_1076),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1012),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1053),
.Y(n_1176)
);

AO22x1_ASAP7_75t_L g1177 ( 
.A1(n_1086),
.A2(n_1049),
.B1(n_1039),
.B2(n_1128),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1131),
.A2(n_1024),
.B(n_1018),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1131),
.A2(n_1024),
.B(n_1018),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1052),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1106),
.B(n_1157),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1090),
.B(n_1138),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1066),
.B(n_1028),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1017),
.A2(n_1096),
.B1(n_1149),
.B2(n_1103),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1090),
.B(n_1035),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1109),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1036),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1032),
.B(n_1148),
.Y(n_1190)
);

INVx2_ASAP7_75t_R g1191 ( 
.A(n_1066),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1074),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1105),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1066),
.B(n_1043),
.Y(n_1194)
);

AND2x2_ASAP7_75t_SL g1195 ( 
.A(n_1055),
.B(n_1108),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1010),
.A2(n_1126),
.B(n_1113),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1141),
.B(n_1048),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1048),
.B(n_1073),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1067),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1043),
.B(n_1139),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1051),
.B(n_1015),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1135),
.B(n_1140),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1025),
.B(n_1133),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1010),
.A2(n_1126),
.B(n_1144),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1037),
.B(n_1119),
.Y(n_1206)
);

AO21x1_ASAP7_75t_L g1207 ( 
.A1(n_1119),
.A2(n_1038),
.B(n_1029),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1064),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1077),
.B(n_1071),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1059),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1148),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1148),
.B(n_1089),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1013),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1013),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_1013),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1115),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1071),
.A2(n_1079),
.B1(n_1156),
.B2(n_1084),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1019),
.B(n_1114),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1139),
.B(n_1050),
.Y(n_1219)
);

AND2x6_ASAP7_75t_L g1220 ( 
.A(n_1050),
.B(n_1072),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1050),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1124),
.B(n_1087),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1060),
.A2(n_1029),
.B(n_1045),
.C(n_1079),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1104),
.A2(n_1116),
.B(n_1110),
.C(n_1127),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1145),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1072),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1137),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_1064),
.B(n_1137),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1085),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1007),
.B(n_1101),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1091),
.B(n_1083),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1155),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1155),
.B(n_1007),
.Y(n_1233)
);

INVx3_ASAP7_75t_SL g1234 ( 
.A(n_1155),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1155),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1007),
.B(n_1101),
.Y(n_1236)
);

INVx3_ASAP7_75t_SL g1237 ( 
.A(n_1154),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1069),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1113),
.A2(n_1144),
.B(n_1118),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1063),
.A2(n_1047),
.B(n_1030),
.C(n_1082),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1101),
.B(n_1065),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1118),
.A2(n_1027),
.B(n_1158),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1081),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1094),
.A2(n_1129),
.B(n_1107),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1068),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1088),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1021),
.Y(n_1247)
);

CKINVDCx8_ASAP7_75t_R g1248 ( 
.A(n_1154),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1041),
.B(n_1044),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1063),
.A2(n_1054),
.B(n_1159),
.C(n_1150),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1143),
.Y(n_1251)
);

AOI222xp33_ASAP7_75t_L g1252 ( 
.A1(n_1054),
.A2(n_1154),
.B1(n_1075),
.B2(n_1057),
.C1(n_1014),
.C2(n_1108),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1065),
.B(n_1040),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1031),
.A2(n_1026),
.B1(n_1142),
.B2(n_1023),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1008),
.A2(n_1100),
.B(n_1153),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1058),
.A2(n_1111),
.B1(n_1117),
.B2(n_1134),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1056),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1136),
.B(n_1016),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1097),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1033),
.A2(n_1011),
.B1(n_1146),
.B2(n_1034),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1053),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1030),
.A2(n_771),
.B(n_969),
.C(n_786),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1009),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1012),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1046),
.A2(n_778),
.B1(n_750),
.B2(n_919),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1053),
.Y(n_1269)
);

AND2x2_ASAP7_75t_SL g1270 ( 
.A(n_1147),
.B(n_938),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1061),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1012),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1009),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1053),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1130),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1061),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1061),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1053),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1053),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1131),
.A2(n_519),
.B(n_1024),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1080),
.B(n_1020),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1080),
.B(n_1020),
.Y(n_1282)
);

AOI21xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1141),
.A2(n_566),
.B(n_606),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_L g1284 ( 
.A(n_1032),
.B(n_866),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1141),
.A2(n_1147),
.B1(n_926),
.B2(n_969),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1020),
.B(n_1022),
.Y(n_1286)
);

AND3x2_ASAP7_75t_L g1287 ( 
.A(n_1147),
.B(n_938),
.C(n_490),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1046),
.B(n_969),
.C(n_1147),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1013),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1092),
.A2(n_1002),
.B1(n_1005),
.B2(n_1095),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1028),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1292)
);

BUFx8_ASAP7_75t_SL g1293 ( 
.A(n_1105),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1032),
.B(n_1148),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1027),
.A2(n_519),
.B(n_650),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1141),
.A2(n_1147),
.B1(n_926),
.B2(n_969),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1066),
.B(n_987),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1079),
.A2(n_971),
.B(n_1021),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1009),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1032),
.B(n_1148),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1023),
.A2(n_1120),
.B(n_1097),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1061),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1242),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1168),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1270),
.A2(n_1296),
.B1(n_1285),
.B2(n_1288),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1172),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1217),
.B(n_1251),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1293),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1193),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1288),
.A2(n_1171),
.B1(n_1173),
.B2(n_1197),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1174),
.A2(n_1198),
.B1(n_1199),
.B2(n_1167),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1171),
.B(n_1181),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1233),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1185),
.B(n_1181),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1268),
.A2(n_1263),
.B1(n_1302),
.B2(n_1301),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1192),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1287),
.A2(n_1206),
.B1(n_1207),
.B2(n_1204),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1176),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1175),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1248),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1264),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1274),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1182),
.B(n_1262),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1166),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1206),
.A2(n_1204),
.B1(n_1163),
.B2(n_1209),
.Y(n_1328)
);

AO21x1_ASAP7_75t_SL g1329 ( 
.A1(n_1202),
.A2(n_1203),
.B(n_1230),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1163),
.A2(n_1164),
.B1(n_1281),
.B2(n_1282),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1188),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1185),
.B(n_1182),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1169),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1299),
.A2(n_1202),
.B1(n_1203),
.B2(n_1275),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1281),
.A2(n_1282),
.B1(n_1290),
.B2(n_1286),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1266),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1236),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1212),
.B(n_1186),
.Y(n_1339)
);

BUFx2_ASAP7_75t_R g1340 ( 
.A(n_1273),
.Y(n_1340)
);

AOI21xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1190),
.A2(n_1294),
.B(n_1303),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1300),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1262),
.B(n_1263),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1161),
.A2(n_1183),
.B1(n_1290),
.B2(n_1292),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1267),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1272),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1189),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1216),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1225),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1276),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1212),
.B(n_1186),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1277),
.Y(n_1352)
);

BUFx4f_ASAP7_75t_SL g1353 ( 
.A(n_1269),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1247),
.B(n_1231),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1278),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1161),
.A2(n_1183),
.B1(n_1297),
.B2(n_1292),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1279),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1222),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1195),
.A2(n_1222),
.B1(n_1178),
.B2(n_1179),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1255),
.A2(n_1242),
.B(n_1280),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1162),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1226),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1305),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1187),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1180),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1297),
.B(n_1301),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1235),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1302),
.B(n_1201),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1218),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1232),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1241),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1211),
.A2(n_1231),
.B1(n_1294),
.B2(n_1303),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1283),
.B(n_1229),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1258),
.Y(n_1374)
);

AO21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1256),
.A2(n_1246),
.B(n_1249),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1208),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1165),
.A2(n_1238),
.B1(n_1280),
.B2(n_1239),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1190),
.A2(n_1303),
.B1(n_1294),
.B2(n_1210),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1190),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1221),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1240),
.B(n_1243),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1284),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1227),
.Y(n_1384)
);

BUFx2_ASAP7_75t_R g1385 ( 
.A(n_1237),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1215),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1177),
.B(n_1265),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1243),
.A2(n_1256),
.B1(n_1196),
.B2(n_1205),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1260),
.A2(n_1249),
.B1(n_1254),
.B2(n_1252),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1228),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1260),
.A2(n_1254),
.B1(n_1252),
.B2(n_1245),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1289),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1220),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1255),
.A2(n_1261),
.B(n_1257),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1298),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1213),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1223),
.B(n_1214),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1298),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1219),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1295),
.A2(n_1259),
.B(n_1224),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1213),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1291),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1291),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1170),
.Y(n_1404)
);

AOI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1250),
.A2(n_1147),
.B1(n_1270),
.B2(n_606),
.C1(n_641),
.C2(n_534),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1191),
.A2(n_1184),
.B(n_1194),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1200),
.B(n_998),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1160),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1248),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1174),
.A2(n_1141),
.B1(n_954),
.B2(n_969),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1196),
.A2(n_1018),
.B(n_1010),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1234),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1160),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1234),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1193),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1160),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1270),
.A2(n_1296),
.B1(n_1285),
.B2(n_1288),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1316),
.B(n_1337),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1306),
.A2(n_1388),
.B(n_1360),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1306),
.A2(n_1387),
.B(n_1360),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1410),
.A2(n_1313),
.B(n_1308),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1375),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1317),
.A2(n_1332),
.B(n_1318),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1358),
.B(n_1339),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1371),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1400),
.A2(n_1389),
.B(n_1391),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1319),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1319),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1354),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1370),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1383),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1354),
.B(n_1310),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1316),
.B(n_1337),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1370),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1381),
.A2(n_1344),
.B(n_1397),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1381),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1315),
.B(n_1356),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1310),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1310),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1341),
.A2(n_1315),
.B(n_1350),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1326),
.B(n_1343),
.Y(n_1441)
);

OR2x6_ASAP7_75t_L g1442 ( 
.A(n_1411),
.B(n_1374),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1411),
.Y(n_1443)
);

AO21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1359),
.A2(n_1320),
.B(n_1377),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1307),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1321),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1326),
.B(n_1343),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1327),
.A2(n_1352),
.B(n_1363),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1333),
.Y(n_1449)
);

INVxp67_ASAP7_75t_R g1450 ( 
.A(n_1368),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1338),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1394),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1361),
.B(n_1312),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1364),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1394),
.Y(n_1455)
);

INVx4_ASAP7_75t_SL g1456 ( 
.A(n_1386),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1368),
.B(n_1366),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1366),
.B(n_1417),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1329),
.B(n_1328),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1324),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1365),
.B(n_1347),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1367),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1329),
.B(n_1339),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1325),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1367),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1330),
.A2(n_1416),
.B(n_1309),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1339),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1405),
.B(n_1335),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1351),
.B(n_1375),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1351),
.B(n_1334),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1408),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1413),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1351),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1406),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1406),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1369),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1406),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1314),
.B(n_1372),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1407),
.A2(n_1403),
.B(n_1402),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1404),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1412),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1380),
.B(n_1384),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1346),
.B(n_1373),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1322),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1322),
.A2(n_1345),
.B1(n_1378),
.B2(n_1409),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1435),
.B(n_1376),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1435),
.B(n_1423),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1479),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1462),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1421),
.A2(n_1379),
.B1(n_1382),
.B2(n_1331),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1435),
.B(n_1345),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1468),
.A2(n_1437),
.B1(n_1458),
.B2(n_1483),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1443),
.B(n_1392),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1422),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1479),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1442),
.B(n_1379),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1475),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1442),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1462),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1442),
.B(n_1398),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1432),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1459),
.B(n_1398),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1440),
.B(n_1355),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1440),
.B(n_1362),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1423),
.B(n_1412),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1459),
.B(n_1398),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1414),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1425),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1440),
.B(n_1357),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1425),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1412),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1453),
.B(n_1312),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1448),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1448),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1431),
.B(n_1395),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1448),
.Y(n_1522)
);

INVx3_ASAP7_75t_SL g1523 ( 
.A(n_1456),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1418),
.B(n_1357),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1432),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1477),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1447),
.B(n_1399),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1494),
.A2(n_1444),
.B1(n_1478),
.B2(n_1426),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1491),
.B(n_1446),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1491),
.B(n_1460),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1486),
.C(n_1438),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1506),
.B(n_1450),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1492),
.A2(n_1478),
.B1(n_1323),
.B2(n_1409),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1488),
.A2(n_1432),
.B(n_1419),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1501),
.B(n_1457),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1506),
.B(n_1450),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1488),
.A2(n_1510),
.B1(n_1509),
.B2(n_1493),
.C(n_1502),
.Y(n_1537)
);

OAI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1510),
.A2(n_1464),
.B1(n_1409),
.B2(n_1323),
.C(n_1485),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1501),
.B(n_1436),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1509),
.A2(n_1470),
.B1(n_1428),
.B2(n_1427),
.C(n_1461),
.Y(n_1540)
);

OA211x2_ASAP7_75t_L g1541 ( 
.A1(n_1502),
.A2(n_1456),
.B(n_1444),
.C(n_1420),
.Y(n_1541)
);

NAND4xp25_ASAP7_75t_L g1542 ( 
.A(n_1487),
.B(n_1493),
.C(n_1507),
.D(n_1515),
.Y(n_1542)
);

NAND4xp25_ASAP7_75t_L g1543 ( 
.A(n_1487),
.B(n_1507),
.C(n_1515),
.D(n_1482),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1505),
.B(n_1430),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1498),
.A2(n_1438),
.B(n_1439),
.C(n_1429),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1518),
.A2(n_1426),
.B1(n_1470),
.B2(n_1323),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1482),
.C(n_1476),
.D(n_1451),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1527),
.A2(n_1476),
.B1(n_1434),
.B2(n_1484),
.C(n_1465),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_SL g1549 ( 
.A(n_1523),
.B(n_1311),
.Y(n_1549)
);

OR2x6_ASAP7_75t_SL g1550 ( 
.A(n_1524),
.B(n_1311),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1489),
.B(n_1439),
.C(n_1484),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1508),
.B(n_1465),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1504),
.B(n_1426),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_L g1554 ( 
.A(n_1489),
.B(n_1466),
.C(n_1431),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1524),
.A2(n_1432),
.B1(n_1385),
.B2(n_1348),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1433),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1498),
.B(n_1424),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1490),
.A2(n_1432),
.B1(n_1463),
.B2(n_1390),
.C(n_1469),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1498),
.B(n_1424),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1497),
.B(n_1466),
.C(n_1426),
.Y(n_1560)
);

OAI221xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1490),
.A2(n_1463),
.B1(n_1473),
.B2(n_1472),
.C(n_1471),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1504),
.A2(n_1424),
.B(n_1422),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1525),
.A2(n_1424),
.B(n_1422),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1521),
.B(n_1449),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1451),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1519),
.A2(n_1455),
.B(n_1452),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1523),
.A2(n_1422),
.B1(n_1467),
.B2(n_1481),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1516),
.B(n_1454),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_1466),
.C(n_1480),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1511),
.B(n_1466),
.C(n_1480),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1566),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1568),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1565),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1500),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1500),
.Y(n_1576)
);

NAND2x1_ASAP7_75t_L g1577 ( 
.A(n_1551),
.B(n_1496),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1569),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1564),
.Y(n_1580)
);

AND2x4_ASAP7_75t_SL g1581 ( 
.A(n_1532),
.B(n_1496),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1557),
.B(n_1499),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1499),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1535),
.B(n_1511),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1539),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1529),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1570),
.B(n_1519),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1537),
.B(n_1526),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1536),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.Y(n_1591)
);

NOR2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1531),
.B(n_1467),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1530),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1571),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1547),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1495),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1559),
.B(n_1517),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1544),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1587),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1596),
.B(n_1546),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1587),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1594),
.B(n_1558),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1573),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1574),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1590),
.B(n_1545),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1520),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1546),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1586),
.B(n_1528),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1572),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1575),
.B(n_1576),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

AOI32xp33_ASAP7_75t_L g1618 ( 
.A1(n_1578),
.A2(n_1528),
.A3(n_1533),
.B1(n_1549),
.B2(n_1555),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1578),
.A2(n_1540),
.B(n_1538),
.C(n_1561),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1580),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1520),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1522),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1626)
);

NAND4xp25_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1541),
.C(n_1563),
.D(n_1517),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1595),
.B(n_1522),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1590),
.B(n_1550),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1550),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1503),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1575),
.B(n_1503),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1603),
.B(n_1445),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1608),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1597),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1629),
.B(n_1595),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1609),
.B(n_1620),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1626),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1606),
.B(n_1575),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1611),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1616),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1630),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1597),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1613),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1630),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1632),
.B(n_1576),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1618),
.B(n_1594),
.C(n_1591),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1632),
.A2(n_1592),
.B1(n_1591),
.B2(n_1588),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1634),
.B(n_1588),
.Y(n_1655)
);

AOI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1628),
.A2(n_1591),
.B(n_1577),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1634),
.B(n_1576),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1627),
.A2(n_1598),
.B(n_1593),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1629),
.A2(n_1598),
.B1(n_1601),
.B2(n_1600),
.C(n_1585),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1615),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1631),
.B(n_1577),
.C(n_1415),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1610),
.B(n_1592),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1615),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1610),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1617),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1660),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1602),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1622),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1649),
.B(n_1624),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1653),
.B(n_1625),
.C(n_1415),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1646),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1639),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1644),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1639),
.B(n_1604),
.Y(n_1680)
);

INVx5_ASAP7_75t_L g1681 ( 
.A(n_1655),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1655),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1645),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1641),
.B(n_1640),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1635),
.B(n_1307),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1662),
.B(n_1582),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1660),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1650),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1642),
.A2(n_1601),
.B1(n_1600),
.B2(n_1621),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1650),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1658),
.B(n_1340),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1654),
.A2(n_1583),
.B1(n_1582),
.B2(n_1581),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1652),
.B(n_1617),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1646),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1599),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1660),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1651),
.A2(n_1605),
.B1(n_1607),
.B2(n_1467),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1661),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1664),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1697),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1677),
.B(n_1637),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1685),
.B(n_1637),
.Y(n_1706)
);

AO221x1_ASAP7_75t_L g1707 ( 
.A1(n_1683),
.A2(n_1664),
.B1(n_1666),
.B2(n_1567),
.C(n_1654),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1673),
.B(n_1659),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1699),
.B(n_1643),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1674),
.B(n_1638),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1674),
.A2(n_1656),
.B(n_1655),
.C(n_1643),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1672),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1672),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1693),
.B(n_1691),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1675),
.B(n_1657),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1681),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_SL g1717 ( 
.A(n_1688),
.B(n_1663),
.C(n_1665),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1697),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1676),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1676),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1698),
.B(n_1648),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1678),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1680),
.B(n_1657),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1680),
.B(n_1648),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1678),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1695),
.A2(n_1656),
.B1(n_1702),
.B2(n_1703),
.C(n_1682),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1679),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1679),
.Y(n_1729)
);

AOI21xp33_ASAP7_75t_L g1730 ( 
.A1(n_1710),
.A2(n_1697),
.B(n_1681),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1696),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1708),
.B(n_1686),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1704),
.B(n_1696),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1698),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1713),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1718),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1718),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1711),
.B(n_1681),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1719),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1721),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1725),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1716),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1722),
.B(n_1669),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1726),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1720),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1707),
.B(n_1669),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1715),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1728),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1739),
.A2(n_1717),
.B1(n_1714),
.B2(n_1711),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1739),
.A2(n_1727),
.B(n_1720),
.C(n_1723),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1733),
.B(n_1724),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1733),
.B(n_1342),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1747),
.A2(n_1681),
.B(n_1723),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_SL g1755 ( 
.A(n_1748),
.B(n_1743),
.C(n_1746),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1730),
.A2(n_1681),
.B(n_1729),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1742),
.A2(n_1697),
.B1(n_1663),
.B2(n_1683),
.C(n_1701),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1735),
.A2(n_1655),
.B1(n_1683),
.B2(n_1667),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1670),
.Y(n_1759)
);

OAI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1744),
.A2(n_1670),
.B(n_1683),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1759),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1753),
.Y(n_1762)
);

NOR3x1_ASAP7_75t_L g1763 ( 
.A(n_1755),
.B(n_1738),
.C(n_1737),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1760),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_1746),
.C(n_1745),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1752),
.B(n_1734),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1750),
.B(n_1745),
.C(n_1736),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1754),
.B(n_1731),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1756),
.B(n_1740),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1758),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1767),
.B(n_1336),
.Y(n_1771)
);

AO21x1_ASAP7_75t_L g1772 ( 
.A1(n_1765),
.A2(n_1749),
.B(n_1741),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1768),
.A2(n_1757),
.B(n_1703),
.C(n_1702),
.Y(n_1773)
);

AOI322xp5_ASAP7_75t_L g1774 ( 
.A1(n_1764),
.A2(n_1665),
.A3(n_1694),
.B1(n_1692),
.B2(n_1690),
.C1(n_1682),
.C2(n_1684),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1770),
.B(n_1684),
.Y(n_1775)
);

INVxp33_ASAP7_75t_SL g1776 ( 
.A(n_1763),
.Y(n_1776)
);

NOR2xp67_ASAP7_75t_L g1777 ( 
.A(n_1775),
.B(n_1761),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1776),
.A2(n_1762),
.B1(n_1766),
.B2(n_1769),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1771),
.Y(n_1779)
);

NOR2xp67_ASAP7_75t_SL g1780 ( 
.A(n_1772),
.B(n_1342),
.Y(n_1780)
);

XNOR2xp5_ASAP7_75t_L g1781 ( 
.A(n_1773),
.B(n_1336),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1774),
.B(n_1671),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1775),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1780),
.B(n_1401),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1782),
.B(n_1671),
.Y(n_1785)
);

NOR2xp67_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1690),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1778),
.A2(n_1692),
.B1(n_1694),
.B2(n_1700),
.Y(n_1787)
);

NOR3xp33_ASAP7_75t_SL g1788 ( 
.A(n_1781),
.B(n_1777),
.C(n_1782),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1784),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1785),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1786),
.B(n_1783),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1788),
.B1(n_1787),
.B2(n_1789),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1793),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1793),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1794),
.A2(n_1790),
.B(n_1791),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1791),
.B(n_1789),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1791),
.B1(n_1700),
.B2(n_1687),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1796),
.Y(n_1799)
);

XNOR2xp5_ASAP7_75t_L g1800 ( 
.A(n_1799),
.B(n_1798),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1800),
.A2(n_1353),
.B1(n_1349),
.B2(n_1348),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_R g1802 ( 
.A1(n_1801),
.A2(n_1689),
.B1(n_1668),
.B2(n_1687),
.C(n_1349),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1689),
.B(n_1668),
.C(n_1396),
.Y(n_1803)
);


endmodule