module real_jpeg_5773_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_52),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_1),
.A2(n_52),
.B1(n_178),
.B2(n_188),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_1),
.A2(n_52),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_2),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_93),
.B(n_94),
.C(n_102),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_80),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_209),
.C(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_28),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_167),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_2),
.B(n_118),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_2),
.A2(n_80),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_24),
.B1(n_87),
.B2(n_90),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_6),
.A2(n_24),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_9),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_201),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_199),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_139),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_15),
.B(n_139),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.C(n_106),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_16),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_56),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_17),
.B(n_57),
.C(n_68),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_19),
.Y(n_193)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_27),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_28),
.B(n_48),
.Y(n_194)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_36),
.Y(n_133)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_42),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_43),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_59),
.B(n_187),
.Y(n_186)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_59)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_65),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_84),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_69),
.B(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_76),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_70),
.B(n_86),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_70),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_76),
.Y(n_218)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_95),
.B(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_80),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_80),
.A2(n_153),
.B(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_84),
.B(n_220),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_87),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_88),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_91),
.A2(n_106),
.B1(n_107),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_91),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_92),
.A2(n_103),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_92),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_101),
.Y(n_231)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_103),
.Y(n_275)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_125),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_117),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_110),
.A2(n_117),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_111),
.B(n_130),
.Y(n_214)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_116),
.B(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_116),
.Y(n_229)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_118),
.B(n_126),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_118),
.B(n_228),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_130),
.B(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_169),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_160),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.A3(n_149),
.B1(n_152),
.B2(n_156),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_168),
.Y(n_160)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_189),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_186),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_194),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_278),
.B(n_283),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_261),
.B(n_277),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_235),
.B(n_260),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_205),
.B(n_215),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_207),
.B1(n_212),
.B2(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_225),
.Y(n_215)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_225)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_233),
.C(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_247),
.B(n_259),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_258),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_268),
.C(n_274),
.Y(n_282)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_282),
.Y(n_283)
);


endmodule