module fake_jpeg_17585_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_17),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_13),
.B1(n_24),
.B2(n_15),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.C(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_20),
.C(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_12),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_33),
.B(n_26),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_18),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_15),
.C(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_29),
.C(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_25),
.B1(n_19),
.B2(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_30),
.C(n_23),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_39),
.C(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_25),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_40),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_45),
.C(n_46),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_48),
.B(n_19),
.Y(n_51)
);


endmodule