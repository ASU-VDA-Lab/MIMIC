module fake_aes_6659_n_636 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_636);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_636;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g71 ( .A(n_70), .Y(n_71) );
INVx1_ASAP7_75t_SL g72 ( .A(n_10), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_62), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_3), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_35), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_16), .Y(n_76) );
HB1xp67_ASAP7_75t_L g77 ( .A(n_55), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_24), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_16), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_3), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_68), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_36), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_52), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_40), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_23), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_14), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_56), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_54), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_34), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_15), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_27), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_19), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_61), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_59), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_67), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_19), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
AND2x6_ASAP7_75t_L g119 ( .A(n_71), .B(n_31), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_88), .B(n_0), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_110), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_115), .B(n_0), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_77), .B(n_1), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_84), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_73), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_90), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_75), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_85), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_90), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_75), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_80), .B(n_2), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_72), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_74), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_114), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_78), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_78), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_89), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
NAND2xp33_ASAP7_75t_R g145 ( .A(n_108), .B(n_33), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_79), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_94), .B(n_2), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_96), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_79), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_82), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_82), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_74), .B(n_4), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_76), .B(n_4), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_116), .Y(n_159) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_116), .B(n_69), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_150), .A2(n_76), .B1(n_92), .B2(n_91), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_154), .B(n_87), .Y(n_163) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_129), .B(n_103), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_149), .B(n_102), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_150), .B(n_97), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_141), .B(n_118), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_122), .B(n_99), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_136), .B(n_91), .Y(n_179) );
AO22x2_ASAP7_75t_L g180 ( .A1(n_123), .A2(n_117), .B1(n_113), .B2(n_104), .Y(n_180) );
CKINVDCx11_ASAP7_75t_R g181 ( .A(n_121), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_135), .Y(n_186) );
CKINVDCx11_ASAP7_75t_R g187 ( .A(n_121), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_122), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_123), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_127), .B(n_117), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_131), .B(n_100), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_127), .B(n_92), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_128), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_130), .B(n_101), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_125), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_133), .B(n_113), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_133), .B(n_105), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_138), .B(n_105), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_139), .B(n_112), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_140), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_146), .B(n_104), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g216 ( .A1(n_120), .A2(n_112), .B1(n_101), .B2(n_103), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_146), .B(n_111), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_147), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_151), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_124), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_152), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
NAND2xp33_ASAP7_75t_SL g227 ( .A(n_172), .B(n_145), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_169), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_212), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_193), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_164), .A2(n_160), .B(n_161), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_212), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_214), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_181), .Y(n_234) );
AOI22xp5_ASAP7_75t_SL g235 ( .A1(n_203), .A2(n_134), .B1(n_95), .B2(n_107), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_180), .B(n_179), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_214), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_163), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_188), .B(n_161), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_179), .B(n_158), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_186), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
BUFx12f_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
AND2x6_ASAP7_75t_SL g248 ( .A(n_203), .B(n_106), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_172), .A2(n_158), .B(n_156), .C(n_153), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_220), .B(n_156), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_164), .B(n_148), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_179), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_204), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
NOR3xp33_ASAP7_75t_SL g259 ( .A(n_216), .B(n_106), .C(n_153), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_163), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_163), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_205), .B(n_111), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_165), .B(n_119), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
BUFx4f_ASAP7_75t_L g266 ( .A(n_163), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_173), .A2(n_93), .B(n_109), .C(n_119), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_177), .Y(n_268) );
NOR3xp33_ASAP7_75t_SL g269 ( .A(n_170), .B(n_93), .C(n_6), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_163), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_201), .Y(n_271) );
AND2x6_ASAP7_75t_L g272 ( .A(n_173), .B(n_119), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_163), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_201), .Y(n_275) );
NOR3xp33_ASAP7_75t_SL g276 ( .A(n_166), .B(n_5), .C(n_6), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_180), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_221), .B(n_119), .Y(n_278) );
OR2x6_ASAP7_75t_L g279 ( .A(n_180), .B(n_119), .Y(n_279) );
NOR3xp33_ASAP7_75t_SL g280 ( .A(n_194), .B(n_5), .C(n_8), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_218), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_180), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_195), .B(n_119), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_183), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_206), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_210), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_187), .Y(n_289) );
BUFx4_ASAP7_75t_SL g290 ( .A(n_187), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_208), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_210), .Y(n_292) );
NOR2xp33_ASAP7_75t_R g293 ( .A(n_182), .B(n_184), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_286), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_240), .B(n_165), .Y(n_295) );
INVx3_ASAP7_75t_SL g296 ( .A(n_236), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_286), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_SL g298 ( .A1(n_267), .A2(n_178), .B(n_224), .C(n_222), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_278), .A2(n_213), .B(n_202), .Y(n_300) );
INVx5_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_260), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_244), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_226), .B(n_167), .Y(n_304) );
BUFx12f_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_226), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_290), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_236), .A2(n_162), .B1(n_165), .B2(n_219), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_263), .A2(n_200), .B(n_199), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_236), .A2(n_207), .B1(n_195), .B2(n_215), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_246), .Y(n_314) );
BUFx4f_ASAP7_75t_L g315 ( .A(n_236), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_291), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_230), .B(n_217), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_228), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_228), .A2(n_282), .B1(n_277), .B2(n_293), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_240), .B(n_176), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_260), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_291), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_240), .B(n_196), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_254), .B(n_185), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_229), .A2(n_211), .B1(n_208), .B2(n_183), .C(n_225), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_243), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_254), .B(n_183), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_273), .Y(n_329) );
BUFx10_ASAP7_75t_L g330 ( .A(n_241), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_275), .B(n_211), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_263), .A2(n_225), .B(n_191), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_284), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_234), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_242), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_279), .A2(n_223), .B1(n_198), .B2(n_197), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_265), .B(n_8), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_275), .B(n_9), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_279), .A2(n_223), .B1(n_198), .B2(n_197), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_260), .B(n_192), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_247), .B(n_252), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_274), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_315), .A2(n_279), .B1(n_251), .B2(n_245), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_255), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_294), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_257), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_341), .A2(n_279), .B(n_267), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_294), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_296), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_300), .A2(n_283), .B(n_249), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_297), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_318), .A2(n_319), .B1(n_304), .B2(n_306), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_304), .A2(n_237), .B1(n_233), .B2(n_232), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_343), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_332), .A2(n_289), .B1(n_234), .B2(n_268), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_297), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_308), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_332), .A2(n_289), .B1(n_266), .B2(n_264), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_330), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_308), .A2(n_249), .B1(n_266), .B2(n_292), .Y(n_366) );
AOI22xp5_ASAP7_75t_SL g367 ( .A1(n_311), .A2(n_263), .B1(n_272), .B2(n_238), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_309), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_343), .B(n_337), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_337), .B(n_274), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_303), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_339), .A2(n_235), .B1(n_266), .B2(n_238), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_313), .A2(n_270), .B1(n_288), .B2(n_250), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_301), .B(n_270), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_322), .A2(n_316), .B1(n_310), .B2(n_320), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_301), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_374), .A2(n_324), .B1(n_335), .B2(n_329), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_357), .A2(n_324), .B1(n_335), .B2(n_329), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_348), .B(n_322), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_373), .A2(n_280), .B(n_276), .C(n_269), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_369), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_356), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_362), .B(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_362), .B(n_330), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_359), .B(n_295), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_369), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_227), .B1(n_340), .B2(n_326), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_358), .A2(n_259), .B1(n_298), .B2(n_239), .C(n_336), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_376), .B(n_369), .Y(n_399) );
OAI21x1_ASAP7_75t_SL g400 ( .A1(n_366), .A2(n_312), .B(n_338), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_370), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_323), .B1(n_331), .B2(n_325), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_360), .A2(n_262), .B(n_248), .C(n_333), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_359), .A2(n_346), .B1(n_366), .B2(n_372), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_227), .B1(n_328), .B2(n_283), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_399), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_399), .B(n_361), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_380), .B(n_347), .Y(n_408) );
INVx4_ASAP7_75t_L g409 ( .A(n_395), .Y(n_409) );
OA211x2_ASAP7_75t_L g410 ( .A1(n_398), .A2(n_355), .B(n_262), .C(n_367), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_391), .B(n_361), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_391), .B(n_361), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_398), .B(n_351), .C(n_355), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_383), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_378), .B(n_365), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_391), .B(n_365), .Y(n_417) );
BUFx12f_ASAP7_75t_L g418 ( .A(n_395), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_383), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_385), .B(n_351), .C(n_365), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_403), .B(n_336), .Y(n_424) );
OAI332xp33_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_363), .A3(n_305), .B1(n_309), .B2(n_364), .B3(n_314), .C1(n_17), .C2(n_18), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_402), .A2(n_364), .B1(n_354), .B2(n_353), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_231), .B(n_327), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_391), .B(n_347), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_380), .B(n_349), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
AOI221xp5_ASAP7_75t_SL g431 ( .A1(n_404), .A2(n_354), .B1(n_353), .B2(n_349), .C(n_377), .Y(n_431) );
AOI211xp5_ASAP7_75t_L g432 ( .A1(n_404), .A2(n_377), .B(n_317), .C(n_314), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_389), .B(n_330), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_389), .B(n_317), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_403), .A2(n_317), .B1(n_371), .B2(n_328), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_391), .B(n_334), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_379), .A2(n_371), .B1(n_328), .B2(n_305), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_385), .A2(n_368), .B1(n_285), .B2(n_327), .C(n_334), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_413), .B(n_379), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_411), .B(n_388), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_422), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_388), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_425), .A2(n_405), .B1(n_401), .B2(n_394), .C(n_400), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_419), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_430), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_419), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_410), .A2(n_395), .B1(n_386), .B2(n_396), .Y(n_451) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_426), .A2(n_392), .A3(n_401), .B(n_394), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_417), .B(n_381), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_432), .A2(n_395), .B1(n_392), .B2(n_394), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_424), .A2(n_396), .B(n_386), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_406), .B(n_395), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_430), .B(n_390), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_418), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx4_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
INVx4_ASAP7_75t_SL g463 ( .A(n_418), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_437), .A2(n_393), .B1(n_382), .B2(n_390), .C(n_381), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_409), .B(n_390), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_371), .B(n_393), .C(n_375), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_439), .B(n_175), .C(n_171), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_407), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_425), .B(n_393), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_415), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_414), .A2(n_400), .B1(n_285), .B2(n_258), .C(n_281), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_441), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_9), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_438), .B(n_10), .Y(n_475) );
INVx4_ASAP7_75t_L g476 ( .A(n_409), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_407), .Y(n_477) );
OAI33xp33_ASAP7_75t_L g478 ( .A1(n_408), .A2(n_429), .A3(n_423), .B1(n_434), .B2(n_433), .B3(n_416), .Y(n_478) );
OAI22xp5_ASAP7_75t_SL g479 ( .A1(n_409), .A2(n_350), .B1(n_375), .B2(n_301), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_421), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_410), .B(n_12), .C(n_15), .D(n_17), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_440), .B(n_18), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_462), .B(n_409), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_444), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_455), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_468), .B(n_416), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_446), .B(n_428), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_470), .B(n_423), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_460), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_458), .A2(n_441), .B1(n_436), .B2(n_427), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_469), .B(n_436), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_453), .B(n_441), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_469), .B(n_435), .Y(n_497) );
INVxp33_ASAP7_75t_L g498 ( .A(n_479), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_477), .B(n_427), .Y(n_499) );
NAND2xp33_ASAP7_75t_SL g500 ( .A(n_473), .B(n_350), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_477), .B(n_20), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_473), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_483), .B(n_20), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_474), .B(n_350), .Y(n_505) );
NAND2xp33_ASAP7_75t_R g506 ( .A(n_471), .B(n_375), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_463), .B(n_350), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_463), .Y(n_509) );
OAI211xp5_ASAP7_75t_SL g510 ( .A1(n_447), .A2(n_168), .B(n_174), .C(n_189), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_481), .B(n_21), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_482), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_463), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_474), .B(n_281), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_442), .B(n_253), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_482), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_475), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_475), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_443), .B(n_25), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_445), .B(n_28), .Y(n_521) );
NOR2xp67_ASAP7_75t_L g522 ( .A(n_462), .B(n_29), .Y(n_522) );
NAND2xp33_ASAP7_75t_R g523 ( .A(n_471), .B(n_465), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_459), .Y(n_524) );
NAND2xp33_ASAP7_75t_R g525 ( .A(n_465), .B(n_32), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_453), .B(n_38), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_450), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_498), .A2(n_458), .B1(n_462), .B2(n_476), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_490), .B(n_480), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_488), .B(n_480), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_492), .B(n_452), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_502), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_503), .B(n_461), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_493), .B(n_478), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_494), .A2(n_454), .B1(n_466), .B2(n_451), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_512), .B(n_457), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_513), .A2(n_464), .B1(n_465), .B2(n_467), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_496), .B(n_461), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_525), .A2(n_456), .B1(n_457), .B2(n_463), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_511), .A2(n_472), .B(n_174), .Y(n_542) );
INVxp67_ASAP7_75t_L g543 ( .A(n_523), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_525), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_484), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_516), .B(n_41), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_517), .B(n_43), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_500), .A2(n_301), .B(n_302), .C(n_307), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_518), .B(n_44), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_491), .B(n_45), .Y(n_550) );
AOI32xp33_ASAP7_75t_L g551 ( .A1(n_500), .A2(n_307), .A3(n_299), .B1(n_321), .B2(n_344), .Y(n_551) );
AOI22xp5_ASAP7_75t_SL g552 ( .A1(n_509), .A2(n_307), .B1(n_299), .B2(n_302), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_487), .Y(n_554) );
AO22x1_ASAP7_75t_L g555 ( .A1(n_508), .A2(n_272), .B1(n_299), .B2(n_321), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_506), .A2(n_272), .B1(n_342), .B2(n_344), .Y(n_556) );
OAI21xp33_ASAP7_75t_SL g557 ( .A1(n_522), .A2(n_523), .B(n_520), .Y(n_557) );
AOI21xp5_ASAP7_75t_SL g558 ( .A1(n_508), .A2(n_345), .B(n_49), .Y(n_558) );
AOI321xp33_ASAP7_75t_L g559 ( .A1(n_497), .A2(n_189), .A3(n_168), .B1(n_192), .B2(n_191), .C(n_63), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_47), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_501), .B(n_50), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_53), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_511), .A2(n_344), .B1(n_321), .B2(n_345), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_489), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_505), .A2(n_345), .B(n_256), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_506), .A2(n_272), .B1(n_345), .B2(n_171), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_499), .B(n_65), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_526), .B(n_66), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_504), .B(n_171), .C(n_175), .Y(n_569) );
INVxp33_ASAP7_75t_SL g570 ( .A(n_529), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_535), .A2(n_510), .B(n_514), .C(n_515), .Y(n_571) );
NOR2xp33_ASAP7_75t_R g572 ( .A(n_544), .B(n_527), .Y(n_572) );
XOR2x2_ASAP7_75t_L g573 ( .A(n_532), .B(n_521), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_557), .B(n_519), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_535), .B(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_540), .B(n_507), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_537), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_545), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_543), .B(n_171), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_553), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_554), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_564), .Y(n_582) );
INVx6_ASAP7_75t_L g583 ( .A(n_531), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_534), .Y(n_584) );
BUFx4f_ASAP7_75t_SL g585 ( .A(n_550), .Y(n_585) );
NAND2xp33_ASAP7_75t_L g586 ( .A(n_539), .B(n_272), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_533), .B(n_175), .Y(n_587) );
CKINVDCx16_ASAP7_75t_R g588 ( .A(n_530), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_175), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_538), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_552), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_562), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_575), .B(n_536), .C(n_559), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_574), .A2(n_541), .B(n_558), .Y(n_594) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_587), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g596 ( .A(n_591), .B(n_551), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_570), .B(n_569), .Y(n_597) );
NOR3xp33_ASAP7_75t_L g598 ( .A(n_586), .B(n_542), .C(n_546), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_588), .B(n_584), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_570), .A2(n_561), .B1(n_563), .B2(n_560), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_573), .A2(n_566), .B(n_556), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_571), .A2(n_549), .B1(n_547), .B2(n_567), .C(n_565), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_590), .B(n_568), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_585), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_583), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_583), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_586), .A2(n_555), .B(n_548), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_573), .A2(n_345), .B(n_256), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_577), .Y(n_609) );
XNOR2x1_ASAP7_75t_L g610 ( .A(n_592), .B(n_578), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_578), .B(n_256), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_599), .B(n_579), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_593), .A2(n_581), .B1(n_580), .B2(n_582), .C(n_572), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_595), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_610), .Y(n_615) );
XNOR2x1_ASAP7_75t_L g616 ( .A(n_610), .B(n_576), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_604), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_597), .A2(n_589), .B(n_607), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_597), .A2(n_609), .B1(n_603), .B2(n_602), .C(n_605), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_600), .A2(n_606), .B1(n_611), .B2(n_598), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_606), .B(n_596), .C(n_593), .Y(n_621) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_610), .A2(n_570), .B(n_597), .Y(n_622) );
AOI221x1_ASAP7_75t_L g623 ( .A1(n_594), .A2(n_608), .B1(n_593), .B2(n_578), .C(n_601), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_615), .A2(n_621), .B1(n_620), .B2(n_618), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_614), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_617), .A2(n_616), .B1(n_612), .B2(n_623), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_622), .B(n_612), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_625), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_627), .Y(n_629) );
XNOR2xp5_ASAP7_75t_L g630 ( .A(n_624), .B(n_617), .Y(n_630) );
INVxp33_ASAP7_75t_L g631 ( .A(n_630), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_628), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_632), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_631), .Y(n_634) );
AOI22xp5_ASAP7_75t_SL g635 ( .A1(n_633), .A2(n_634), .B1(n_628), .B2(n_627), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_626), .B1(n_629), .B2(n_619), .C(n_613), .Y(n_636) );
endmodule