module real_jpeg_30175_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_300, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_300;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_197;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_216;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_73),
.B1(n_74),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_0),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_0),
.A2(n_32),
.B1(n_35),
.B2(n_99),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_99),
.Y(n_185)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_3),
.A2(n_32),
.B1(n_35),
.B2(n_54),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_73),
.B1(n_74),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_5),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_32),
.B1(n_35),
.B2(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_122),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_6),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_6),
.A2(n_73),
.B1(n_74),
.B2(n_147),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_46),
.B1(n_73),
.B2(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_9),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_10),
.A2(n_32),
.B1(n_35),
.B2(n_76),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_241)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_11),
.B(n_32),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_26),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_13),
.A2(n_25),
.B(n_26),
.C(n_135),
.D(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_13),
.B(n_48),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_84),
.B(n_152),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_44),
.B(n_47),
.C(n_183),
.D(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_44),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_69),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_13),
.A2(n_71),
.B(n_74),
.C(n_227),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_13),
.A2(n_73),
.B1(n_74),
.B2(n_167),
.Y(n_232)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

XNOR2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_56),
.B2(n_80),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_25),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_25),
.A2(n_31),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_26),
.A2(n_45),
.A3(n_183),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_27),
.A2(n_29),
.A3(n_35),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_27),
.B(n_50),
.Y(n_195)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_32),
.B(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_35),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_45),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_44),
.A2(n_70),
.B(n_167),
.Y(n_227)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_47),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_47),
.A2(n_48),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_79),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_63),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_62),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_62),
.A2(n_63),
.B1(n_114),
.B2(n_241),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_63),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_63),
.A2(n_148),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_68),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_68),
.A2(n_69),
.B1(n_121),
.B2(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_77),
.B(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_77),
.A2(n_97),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_95),
.B1(n_96),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_104),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_89),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_154),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_84),
.A2(n_88),
.B1(n_192),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_84),
.A2(n_86),
.B1(n_111),
.B2(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_87),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_87),
.A2(n_170),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_87),
.A2(n_160),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_88),
.A2(n_159),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_167),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_107),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_287)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_107),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_115),
.C(n_119),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_108),
.A2(n_109),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_110),
.B(n_113),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_115),
.B(n_119),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_116),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_117),
.A2(n_118),
.B(n_203),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_279),
.A3(n_288),
.B1(n_293),
.B2(n_298),
.C(n_300),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_243),
.C(n_275),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_217),
.B(n_242),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_197),
.B(n_216),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_178),
.B(n_196),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_155),
.B(n_177),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_133),
.B(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_137),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_145),
.C(n_150),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_164),
.B(n_176),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_163),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_175),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.C(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_193),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_199),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_212),
.C(n_213),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_206),
.C(n_209),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_222),
.C(n_230),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_236),
.C(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_262),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_245),
.B(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.C(n_261),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_249),
.C(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_256),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_271),
.C(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_277),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);


endmodule