module fake_jpeg_4054_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_20),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_39),
.B1(n_28),
.B2(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_20),
.B1(n_27),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_38),
.B1(n_27),
.B2(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_36),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_82),
.B1(n_26),
.B2(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_39),
.B1(n_41),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_35),
.B1(n_34),
.B2(n_48),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_68),
.Y(n_91)
);

OR2x4_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_79),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_34),
.B1(n_35),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_75),
.B1(n_29),
.B2(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_80),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_39),
.B(n_42),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_24),
.B(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_47),
.C(n_37),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_78),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_28),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_30),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp67_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_16),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_77),
.B(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_105),
.B1(n_107),
.B2(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_101),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_1),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_76),
.C(n_79),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_119),
.C(n_124),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_96),
.B(n_104),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_58),
.B1(n_82),
.B2(n_71),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_105),
.B1(n_86),
.B2(n_85),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_123),
.B1(n_125),
.B2(n_128),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_80),
.C(n_37),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_126),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_59),
.B1(n_62),
.B2(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_37),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_53),
.B1(n_37),
.B2(n_31),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_147),
.B(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_148),
.C(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_88),
.B(n_106),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_144),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_106),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_95),
.B1(n_90),
.B2(n_17),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_17),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_152),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_148),
.B(n_140),
.C(n_142),
.D(n_134),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_162),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_163),
.C(n_2),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_129),
.B1(n_127),
.B2(n_122),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_121),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_17),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_149),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_146),
.B1(n_144),
.B2(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_168),
.B1(n_172),
.B2(n_171),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_135),
.B1(n_22),
.B2(n_4),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_8),
.C(n_10),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_8),
.C(n_13),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_159),
.B1(n_160),
.B2(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_155),
.B(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_183),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_169),
.B(n_165),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_184),
.B(n_15),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_185),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_5),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_6),
.B1(n_185),
.B2(n_178),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_190),
.B(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_6),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_191),
.A2(n_182),
.B(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_178),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_196),
.B(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_192),
.C(n_199),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_201),
.Y(n_205)
);


endmodule