module fake_netlist_1_4530_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_2), .B(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_1), .B(n_6), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_9), .A2(n_7), .B1(n_0), .B2(n_1), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_9), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_8), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_11), .B(n_4), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_11), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_20) );
INVx5_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_13), .B(n_5), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_13), .Y(n_23) );
NAND2xp5_ASAP7_75t_SL g24 ( .A(n_15), .B(n_8), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_21), .B(n_16), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_22), .A2(n_17), .B1(n_18), .B2(n_14), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_28), .B(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_26), .Y(n_32) );
NAND4xp25_ASAP7_75t_SL g33 ( .A(n_31), .B(n_20), .C(n_12), .D(n_24), .Y(n_33) );
AOI21xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_31), .B(n_21), .Y(n_34) );
INVx1_ASAP7_75t_SL g35 ( .A(n_33), .Y(n_35) );
NOR4xp25_ASAP7_75t_SL g36 ( .A(n_34), .B(n_19), .C(n_10), .D(n_22), .Y(n_36) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_35), .B(n_22), .Y(n_37) );
OR5x1_ASAP7_75t_L g38 ( .A(n_37), .B(n_10), .C(n_21), .D(n_23), .E(n_36), .Y(n_38) );
AOI222xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_21), .B1(n_23), .B2(n_36), .C1(n_35), .C2(n_13), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_21), .B1(n_23), .B2(n_37), .Y(n_40) );
endmodule