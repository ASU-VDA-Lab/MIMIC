module fake_jpeg_9725_n_74 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_73;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_59;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_42),
.C(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_45),
.B1(n_15),
.B2(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_4),
.B(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_36),
.B1(n_8),
.B2(n_9),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_36),
.B1(n_10),
.B2(n_11),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_18),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_60),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_66),
.Y(n_71)
);

AOI21x1_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_62),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_59),
.A3(n_65),
.B1(n_51),
.B2(n_28),
.C1(n_23),
.C2(n_24),
.Y(n_74)
);


endmodule