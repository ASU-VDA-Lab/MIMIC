module real_aes_14835_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_372;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_0), .A2(n_100), .B1(n_885), .B2(n_893), .Y(n_99) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_1), .A2(n_49), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g240 ( .A(n_1), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_2), .B(n_187), .Y(n_536) );
AND2x2_ASAP7_75t_L g199 ( .A(n_3), .B(n_189), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_4), .B(n_266), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_5), .A2(n_95), .B1(n_220), .B2(n_233), .C(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_6), .B(n_600), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_7), .B(n_174), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_8), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_9), .B(n_143), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_10), .B(n_233), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_11), .B(n_143), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_12), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_13), .B(n_289), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_14), .Y(n_584) );
BUFx3_ASAP7_75t_L g145 ( .A(n_15), .Y(n_145) );
INVx1_ASAP7_75t_L g156 ( .A(n_15), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_16), .B(n_158), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_17), .B(n_180), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_18), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_19), .Y(n_282) );
BUFx10_ASAP7_75t_L g120 ( .A(n_20), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_21), .B(n_220), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_22), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_23), .B(n_166), .Y(n_279) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_23), .A2(n_69), .B(n_324), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_24), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_25), .B(n_187), .Y(n_594) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_26), .A2(n_191), .B(n_225), .C(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_27), .B(n_220), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_28), .B(n_180), .Y(n_628) );
NAND2xp33_ASAP7_75t_L g539 ( .A(n_29), .B(n_159), .Y(n_539) );
INVx1_ASAP7_75t_L g164 ( .A(n_30), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_31), .A2(n_160), .B(n_574), .C(n_576), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_32), .B(n_148), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_33), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_34), .B(n_225), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_35), .B(n_147), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_36), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
AND3x2_ASAP7_75t_L g884 ( .A(n_37), .B(n_117), .C(n_118), .Y(n_884) );
AO221x1_ASAP7_75t_L g545 ( .A1(n_38), .A2(n_85), .B1(n_178), .B2(n_189), .C(n_220), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_39), .B(n_284), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_40), .B(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g163 ( .A(n_41), .B(n_164), .Y(n_163) );
NAND2x1_ASAP7_75t_L g188 ( .A(n_42), .B(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_43), .Y(n_288) );
INVx1_ASAP7_75t_L g183 ( .A(n_44), .Y(n_183) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_45), .B(n_154), .C(n_160), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_46), .Y(n_257) );
AND2x2_ASAP7_75t_L g198 ( .A(n_47), .B(n_154), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_48), .B(n_147), .Y(n_304) );
INVx1_ASAP7_75t_L g239 ( .A(n_49), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_50), .A2(n_122), .B1(n_865), .B2(n_866), .Y(n_121) );
INVx1_ASAP7_75t_L g865 ( .A(n_50), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_51), .B(n_174), .Y(n_269) );
INVx1_ASAP7_75t_L g139 ( .A(n_52), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_53), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_54), .A2(n_200), .B(n_643), .C(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_55), .B(n_154), .Y(n_205) );
INVx2_ASAP7_75t_L g645 ( .A(n_56), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_57), .B(n_174), .Y(n_612) );
AND2x4_ASAP7_75t_L g891 ( .A(n_58), .B(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_59), .B(n_166), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_60), .B(n_187), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g111 ( .A(n_61), .B(n_77), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_62), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_63), .B(n_283), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_64), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g892 ( .A(n_65), .Y(n_892) );
AND2x2_ASAP7_75t_L g203 ( .A(n_66), .B(n_174), .Y(n_203) );
AND2x2_ASAP7_75t_L g601 ( .A(n_67), .B(n_174), .Y(n_601) );
INVx1_ASAP7_75t_L g550 ( .A(n_68), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_69), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_70), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_71), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_72), .B(n_147), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_73), .Y(n_237) );
INVx2_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
AND3x2_ASAP7_75t_L g887 ( .A(n_74), .B(n_117), .C(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_75), .B(n_310), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_76), .A2(n_80), .B1(n_143), .B2(n_187), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_78), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_79), .B(n_160), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_81), .B(n_167), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_82), .B(n_154), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_83), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_84), .B(n_219), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_86), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_87), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g651 ( .A(n_88), .B(n_167), .Y(n_651) );
INVx1_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
BUFx3_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
INVx1_ASAP7_75t_L g192 ( .A(n_89), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_90), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_91), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_92), .B(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_93), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
INVx1_ASAP7_75t_L g874 ( .A(n_93), .Y(n_874) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_94), .B(n_284), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_96), .B(n_174), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_97), .B(n_265), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_98), .Y(n_634) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_112), .Y(n_100) );
INVxp67_ASAP7_75t_L g879 ( .A(n_101), .Y(n_879) );
NOR2xp67_ASAP7_75t_SL g101 ( .A(n_102), .B(n_103), .Y(n_101) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g878 ( .A(n_106), .Y(n_878) );
NOR2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g118 ( .A(n_108), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
BUFx2_ASAP7_75t_L g126 ( .A(n_110), .Y(n_126) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_111), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_121), .B(n_867), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx5_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_120), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_120), .B(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g866 ( .A(n_122), .Y(n_866) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B(n_524), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_123), .B(n_525), .Y(n_524) );
CKINVDCx10_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g888 ( .A(n_126), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_453), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_400), .C(n_430), .Y(n_128) );
NAND4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_328), .C(n_367), .D(n_380), .Y(n_129) );
AOI332xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_228), .A3(n_245), .B1(n_270), .B2(n_275), .B3(n_296), .C1(n_314), .C2(n_318), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_194), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_169), .Y(n_132) );
INVx2_ASAP7_75t_L g271 ( .A(n_133), .Y(n_271) );
AND2x2_ASAP7_75t_L g385 ( .A(n_133), .B(n_170), .Y(n_385) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g340 ( .A(n_134), .Y(n_340) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_140), .B(n_165), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g324 ( .A(n_137), .Y(n_324) );
INVxp67_ASAP7_75t_L g635 ( .A(n_137), .Y(n_635) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_138), .Y(n_174) );
INVx1_ASAP7_75t_L g241 ( .A(n_139), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_162), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_143), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_144), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g254 ( .A(n_144), .Y(n_254) );
INVx2_ASAP7_75t_L g263 ( .A(n_144), .Y(n_263) );
INVx2_ASAP7_75t_L g289 ( .A(n_144), .Y(n_289) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_145), .Y(n_159) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
INVx2_ASAP7_75t_L g284 ( .A(n_148), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_149), .A2(n_216), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_149), .A2(n_261), .B(n_264), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_149), .A2(n_309), .B(n_311), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_149), .A2(n_598), .B(n_599), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_149), .A2(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g650 ( .A(n_149), .Y(n_650) );
BUFx10_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx3_ASAP7_75t_L g234 ( .A(n_151), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_160), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
INVx2_ASAP7_75t_L g225 ( .A(n_155), .Y(n_225) );
INVx2_ASAP7_75t_L g266 ( .A(n_155), .Y(n_266) );
INVx1_ASAP7_75t_L g582 ( .A(n_155), .Y(n_582) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
INVx3_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVx2_ASAP7_75t_L g559 ( .A(n_159), .Y(n_559) );
INVx2_ASAP7_75t_L g600 ( .A(n_159), .Y(n_600) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_161), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g286 ( .A(n_161), .Y(n_286) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_162), .A2(n_176), .B(n_185), .Y(n_175) );
INVx1_ASAP7_75t_L g227 ( .A(n_162), .Y(n_227) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_162), .A2(n_606), .B(n_609), .Y(n_605) );
BUFx6f_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx2_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
INVx1_ASAP7_75t_L g293 ( .A(n_163), .Y(n_293) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_167), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g391 ( .A(n_169), .B(n_340), .Y(n_391) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g274 ( .A(n_170), .Y(n_274) );
AND2x4_ASAP7_75t_SL g315 ( .A(n_170), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_170), .B(n_196), .Y(n_343) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_170), .Y(n_361) );
AND2x2_ASAP7_75t_L g387 ( .A(n_170), .B(n_340), .Y(n_387) );
INVx1_ASAP7_75t_L g434 ( .A(n_170), .Y(n_434) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_193), .Y(n_171) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_172), .A2(n_533), .B(n_540), .Y(n_532) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVxp33_ASAP7_75t_L g209 ( .A(n_174), .Y(n_209) );
INVx1_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_174), .Y(n_250) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_174), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_174), .B(n_211), .Y(n_564) );
INVx2_ASAP7_75t_L g592 ( .A(n_174), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_181), .Y(n_176) );
INVx1_ASAP7_75t_L g560 ( .A(n_178), .Y(n_560) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_184), .Y(n_181) );
AOI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_188), .B(n_190), .Y(n_185) );
INVx1_ASAP7_75t_L g306 ( .A(n_187), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_190), .A2(n_223), .B(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_190), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g307 ( .A(n_191), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_191), .A2(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx3_ASAP7_75t_L g201 ( .A(n_192), .Y(n_201) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g357 ( .A(n_195), .Y(n_357) );
INVx1_ASAP7_75t_L g488 ( .A(n_195), .Y(n_488) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_212), .Y(n_195) );
INVx2_ASAP7_75t_L g316 ( .A(n_196), .Y(n_316) );
AND2x2_ASAP7_75t_L g362 ( .A(n_196), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g417 ( .A(n_196), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_196), .B(n_434), .Y(n_465) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_202), .B(n_208), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g207 ( .A(n_201), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_201), .A2(n_538), .B(n_539), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AOI21xp33_ASAP7_75t_L g208 ( .A1(n_203), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_210), .A2(n_534), .B(n_537), .Y(n_533) );
AND2x4_ASAP7_75t_L g591 ( .A(n_210), .B(n_592), .Y(n_591) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_210), .A2(n_635), .B(n_651), .Y(n_652) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_211), .B(n_232), .C(n_235), .Y(n_231) );
NOR2xp33_ASAP7_75t_R g548 ( .A(n_211), .B(n_294), .Y(n_548) );
INVx1_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
AND2x2_ASAP7_75t_L g338 ( .A(n_212), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g363 ( .A(n_212), .Y(n_363) );
INVx1_ASAP7_75t_L g384 ( .A(n_212), .Y(n_384) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_212), .Y(n_388) );
AND2x2_ASAP7_75t_L g398 ( .A(n_212), .B(n_316), .Y(n_398) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_222), .B(n_226), .Y(n_214) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g233 ( .A(n_221), .Y(n_233) );
INVx1_ASAP7_75t_L g440 ( .A(n_228), .Y(n_440) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g298 ( .A(n_229), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g449 ( .A(n_229), .B(n_423), .Y(n_449) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g334 ( .A(n_230), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g373 ( .A(n_230), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g406 ( .A(n_230), .B(n_300), .Y(n_406) );
INVx1_ASAP7_75t_L g496 ( .A(n_230), .Y(n_496) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_238), .B(n_242), .Y(n_230) );
NAND2xp33_ASAP7_75t_L g325 ( .A(n_231), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g310 ( .A(n_233), .Y(n_310) );
INVx2_ASAP7_75t_L g575 ( .A(n_233), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_233), .B(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_234), .A2(n_253), .B1(n_255), .B2(n_259), .Y(n_252) );
INVx2_ASAP7_75t_SL g258 ( .A(n_234), .Y(n_258) );
INVx1_ASAP7_75t_L g291 ( .A(n_234), .Y(n_291) );
AOI21xp5_ASAP7_75t_SL g593 ( .A1(n_234), .A2(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_238), .B(n_267), .Y(n_571) );
INVx2_ASAP7_75t_L g586 ( .A(n_238), .Y(n_586) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_241), .Y(n_238) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_239), .A2(n_240), .B(n_241), .Y(n_294) );
NOR2xp33_ASAP7_75t_R g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_247), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g372 ( .A(n_247), .Y(n_372) );
INVx2_ASAP7_75t_L g394 ( .A(n_247), .Y(n_394) );
OR2x2_ASAP7_75t_L g468 ( .A(n_247), .B(n_322), .Y(n_468) );
AND2x2_ASAP7_75t_L g507 ( .A(n_247), .B(n_298), .Y(n_507) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .B(n_269), .Y(n_248) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_249), .A2(n_251), .B(n_269), .Y(n_295) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_249), .A2(n_302), .B(n_313), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_249), .A2(n_302), .B(n_313), .Y(n_335) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_260), .B(n_267), .Y(n_251) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_266), .A2(n_288), .B1(n_289), .B2(n_290), .C(n_291), .Y(n_287) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
NOR2x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g317 ( .A(n_271), .Y(n_317) );
AND2x2_ASAP7_75t_L g439 ( .A(n_271), .B(n_424), .Y(n_439) );
AND2x2_ASAP7_75t_L g444 ( .A(n_271), .B(n_315), .Y(n_444) );
AND2x2_ASAP7_75t_L g519 ( .A(n_271), .B(n_362), .Y(n_519) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g411 ( .A(n_273), .Y(n_411) );
INVx1_ASAP7_75t_L g470 ( .A(n_274), .Y(n_470) );
AND2x2_ASAP7_75t_L g485 ( .A(n_274), .B(n_486), .Y(n_485) );
OAI211xp5_ASAP7_75t_SL g503 ( .A1(n_275), .A2(n_504), .B(n_506), .C(n_508), .Y(n_503) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_276), .B(n_298), .Y(n_389) );
AND2x2_ASAP7_75t_L g429 ( .A(n_276), .B(n_334), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_276), .B(n_406), .Y(n_441) );
AND2x2_ASAP7_75t_L g448 ( .A(n_276), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_295), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g333 ( .A(n_278), .Y(n_333) );
AND2x2_ASAP7_75t_L g346 ( .A(n_278), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g375 ( .A(n_278), .Y(n_375) );
AND2x2_ASAP7_75t_L g478 ( .A(n_278), .B(n_295), .Y(n_478) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_280), .B(n_323), .C(n_325), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .C(n_292), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_285), .C(n_286), .Y(n_281) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_286), .A2(n_562), .B(n_563), .Y(n_561) );
O2A1O1Ixp5_ASAP7_75t_L g606 ( .A1(n_286), .A2(n_310), .B(n_607), .C(n_608), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_286), .A2(n_627), .B(n_628), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g327 ( .A(n_294), .Y(n_327) );
INVx1_ASAP7_75t_L g425 ( .A(n_295), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_296), .A2(n_424), .B(n_444), .C(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g348 ( .A(n_299), .Y(n_348) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_308), .B(n_312), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_307), .Y(n_303) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_L g482 ( .A(n_315), .Y(n_482) );
AND2x2_ASAP7_75t_L g502 ( .A(n_315), .B(n_388), .Y(n_502) );
BUFx2_ASAP7_75t_L g451 ( .A(n_316), .Y(n_451) );
OR2x2_ASAP7_75t_L g464 ( .A(n_317), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g512 ( .A(n_318), .Y(n_512) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g370 ( .A(n_319), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_319), .B(n_371), .Y(n_399) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
OR2x2_ASAP7_75t_L g393 ( .A(n_322), .B(n_394), .Y(n_393) );
OAI21x1_ASAP7_75t_L g604 ( .A1(n_324), .A2(n_605), .B(n_612), .Y(n_604) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_327), .B(n_550), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_336), .B1(n_344), .B2(n_349), .C(n_351), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g424 ( .A(n_333), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g435 ( .A(n_334), .B(n_372), .Y(n_435) );
AND2x2_ASAP7_75t_L g471 ( .A(n_334), .B(n_424), .Y(n_471) );
AND2x2_ASAP7_75t_L g518 ( .A(n_334), .B(n_478), .Y(n_518) );
INVx1_ASAP7_75t_L g423 ( .A(n_335), .Y(n_423) );
NOR2xp67_ASAP7_75t_SL g336 ( .A(n_337), .B(n_341), .Y(n_336) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_337), .B(n_416), .C(n_463), .D(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g349 ( .A(n_338), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_338), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
INVx1_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_339), .Y(n_452) );
AND2x2_ASAP7_75t_L g461 ( .A(n_339), .B(n_350), .Y(n_461) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g486 ( .A(n_340), .B(n_417), .Y(n_486) );
INVx1_ASAP7_75t_L g409 ( .A(n_341), .Y(n_409) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g427 ( .A(n_342), .B(n_384), .Y(n_427) );
AND2x4_ASAP7_75t_L g442 ( .A(n_342), .B(n_411), .Y(n_442) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g350 ( .A(n_343), .Y(n_350) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_346), .B(n_406), .Y(n_413) );
INVx1_ASAP7_75t_L g510 ( .A(n_346), .Y(n_510) );
BUFx3_ASAP7_75t_L g404 ( .A(n_347), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_348), .B(n_439), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B(n_358), .C(n_364), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_354), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g390 ( .A(n_357), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g432 ( .A(n_357), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g436 ( .A(n_357), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_359), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_361), .Y(n_419) );
INVx1_ASAP7_75t_L g401 ( .A(n_362), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_362), .B(n_379), .Y(n_476) );
OR2x2_ASAP7_75t_L g416 ( .A(n_363), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g491 ( .A(n_363), .Y(n_491) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_373), .B(n_376), .Y(n_367) );
INVxp33_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_373), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_431) );
AND2x2_ASAP7_75t_L g405 ( .A(n_374), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g459 ( .A(n_374), .Y(n_459) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_389), .B1(n_390), .B2(n_392), .C1(n_395), .C2(n_399), .Y(n_380) );
NAND2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x2_ASAP7_75t_L g428 ( .A(n_384), .B(n_387), .Y(n_428) );
AND2x2_ASAP7_75t_L g499 ( .A(n_384), .B(n_470), .Y(n_499) );
INVx1_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_387), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_391), .B(n_415), .Y(n_446) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_395), .A2(n_429), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_407), .C(n_426), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_405), .A2(n_444), .B1(n_448), .B2(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g505 ( .A(n_406), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_412), .B1(n_414), .B2(n_420), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g460 ( .A(n_410), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g523 ( .A(n_411), .B(n_482), .Y(n_523) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_415), .A2(n_439), .A3(n_440), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_422), .B(n_424), .Y(n_421) );
INVx2_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_424), .B(n_440), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_424), .B(n_458), .Y(n_513) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_429), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_427), .A2(n_502), .B1(n_503), .B2(n_511), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g430 ( .A(n_431), .B(n_438), .C(n_443), .D(n_447), .Y(n_430) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_440), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g489 ( .A(n_441), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_441), .A2(n_491), .B(n_492), .Y(n_490) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_500), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_472), .C(n_490), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_460), .B1(n_462), .B2(n_466), .C1(n_469), .C2(n_471), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OR2x2_ASAP7_75t_L g467 ( .A(n_458), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g477 ( .A(n_458), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g521 ( .A(n_468), .Y(n_521) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B1(n_477), .B2(n_479), .C(n_483), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g494 ( .A(n_478), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B(n_489), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_491), .A2(n_493), .B(n_497), .C(n_499), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_491), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_514), .C(n_517), .D(n_520), .Y(n_500) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g520 ( .A1(n_518), .A2(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g873 ( .A(n_525), .Y(n_873) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_526), .B(n_716), .C(n_783), .D(n_825), .Y(n_525) );
NOR3x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_669), .C(n_710), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI211x1_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_565), .B(n_613), .C(n_653), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_541), .Y(n_529) );
OAI32xp33_ASAP7_75t_L g613 ( .A1(n_530), .A2(n_614), .A3(n_618), .B1(n_621), .B2(n_637), .Y(n_613) );
INVx2_ASAP7_75t_SL g823 ( .A(n_530), .Y(n_823) );
AND2x4_ASAP7_75t_L g840 ( .A(n_530), .B(n_712), .Y(n_840) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g636 ( .A(n_532), .B(n_551), .Y(n_636) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_532), .Y(n_668) );
INVx1_ASAP7_75t_L g674 ( .A(n_532), .Y(n_674) );
INVx1_ASAP7_75t_L g690 ( .A(n_532), .Y(n_690) );
AND2x2_ASAP7_75t_L g698 ( .A(n_532), .B(n_624), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_532), .B(n_551), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_541), .A2(n_697), .B(n_778), .C(n_782), .Y(n_777) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
OR2x2_ASAP7_75t_L g688 ( .A(n_543), .B(n_689), .Y(n_688) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_543), .B(n_623), .Y(n_744) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_551), .Y(n_543) );
INVx2_ASAP7_75t_SL g662 ( .A(n_544), .Y(n_662) );
AND2x2_ASAP7_75t_L g675 ( .A(n_544), .B(n_666), .Y(n_675) );
AND2x2_ASAP7_75t_L g684 ( .A(n_544), .B(n_667), .Y(n_684) );
AND2x2_ASAP7_75t_L g701 ( .A(n_544), .B(n_664), .Y(n_701) );
BUFx3_ASAP7_75t_L g729 ( .A(n_544), .Y(n_729) );
AND2x2_ASAP7_75t_L g824 ( .A(n_544), .B(n_663), .Y(n_824) );
OR2x2_ASAP7_75t_L g857 ( .A(n_544), .B(n_674), .Y(n_857) );
AO31x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .A3(n_548), .B(n_549), .Y(n_544) );
INVx3_ASAP7_75t_L g664 ( .A(n_551), .Y(n_664) );
AND2x2_ASAP7_75t_L g673 ( .A(n_551), .B(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_561), .B(n_564), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_560), .Y(n_556) );
INVx2_ASAP7_75t_L g631 ( .A(n_559), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_560), .A2(n_580), .B(n_583), .Y(n_579) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_587), .Y(n_566) );
AND2x4_ASAP7_75t_L g694 ( .A(n_567), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g714 ( .A(n_567), .B(n_715), .Y(n_714) );
NAND2x1_ASAP7_75t_L g793 ( .A(n_567), .B(n_730), .Y(n_793) );
INVx5_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_SL g619 ( .A(n_568), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g734 ( .A(n_568), .B(n_729), .Y(n_734) );
AND2x4_ASAP7_75t_L g738 ( .A(n_568), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g763 ( .A(n_568), .B(n_640), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_568), .B(n_587), .Y(n_854) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVxp67_ASAP7_75t_L g709 ( .A(n_569), .Y(n_709) );
AO21x1_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_572), .B(n_578), .Y(n_569) );
AO21x2_ASAP7_75t_L g723 ( .A1(n_570), .A2(n_572), .B(n_578), .Y(n_723) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI21x1_ASAP7_75t_SL g578 ( .A1(n_571), .A2(n_579), .B(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g643 ( .A(n_582), .Y(n_643) );
INVx1_ASAP7_75t_L g681 ( .A(n_587), .Y(n_681) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_602), .Y(n_587) );
INVx3_ASAP7_75t_L g678 ( .A(n_588), .Y(n_678) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g616 ( .A(n_589), .Y(n_616) );
OR2x2_ASAP7_75t_L g656 ( .A(n_589), .B(n_641), .Y(n_656) );
AND2x2_ASAP7_75t_L g732 ( .A(n_589), .B(n_604), .Y(n_732) );
AND2x2_ASAP7_75t_L g850 ( .A(n_589), .B(n_603), .Y(n_850) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_590), .B(n_596), .Y(n_589) );
NAND2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
AOI21x1_ASAP7_75t_L g596 ( .A1(n_591), .A2(n_597), .B(n_601), .Y(n_596) );
O2A1O1Ixp5_ASAP7_75t_L g625 ( .A1(n_591), .A2(n_626), .B(n_629), .C(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g638 ( .A(n_602), .Y(n_638) );
OR2x2_ASAP7_75t_L g702 ( .A(n_602), .B(n_656), .Y(n_702) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g617 ( .A(n_603), .Y(n_617) );
INVx1_ASAP7_75t_L g658 ( .A(n_603), .Y(n_658) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVxp33_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
OR2x2_ASAP7_75t_L g782 ( .A(n_614), .B(n_776), .Y(n_782) );
INVx1_ASAP7_75t_L g815 ( .A(n_614), .Y(n_815) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g739 ( .A(n_615), .B(n_641), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_615), .B(n_680), .Y(n_781) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g640 ( .A(n_616), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g679 ( .A(n_617), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g796 ( .A(n_617), .B(n_723), .Y(n_796) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g788 ( .A(n_619), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g843 ( .A(n_620), .B(n_623), .Y(n_843) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g733 ( .A(n_622), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_636), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_623), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g787 ( .A(n_623), .Y(n_787) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g667 ( .A(n_624), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_624), .B(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_624), .Y(n_801) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_632), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
AND2x4_ASAP7_75t_SL g746 ( .A(n_636), .B(n_662), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_636), .B(n_729), .Y(n_772) );
AND2x2_ASAP7_75t_L g800 ( .A(n_636), .B(n_801), .Y(n_800) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g742 ( .A(n_638), .B(n_640), .Y(n_742) );
AND2x2_ASAP7_75t_L g750 ( .A(n_638), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g790 ( .A(n_638), .Y(n_790) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_640), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g680 ( .A(n_641), .Y(n_680) );
INVx2_ASAP7_75t_L g687 ( .A(n_641), .Y(n_687) );
INVx1_ASAP7_75t_L g753 ( .A(n_641), .Y(n_753) );
AND2x2_ASAP7_75t_L g859 ( .A(n_641), .B(n_722), .Y(n_859) );
AO21x2_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_646), .B(n_652), .Y(n_641) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_643), .B(n_645), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B(n_651), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AOI21x1_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_SL g715 ( .A(n_655), .B(n_658), .Y(n_715) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g720 ( .A(n_656), .Y(n_720) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_658), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g811 ( .A(n_658), .Y(n_811) );
OR2x2_ASAP7_75t_L g834 ( .A(n_658), .B(n_781), .Y(n_834) );
OR2x6_ASAP7_75t_L g659 ( .A(n_660), .B(n_665), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_661), .Y(n_827) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g806 ( .A(n_662), .B(n_769), .Y(n_806) );
INVx1_ASAP7_75t_L g726 ( .A(n_663), .Y(n_726) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_664), .B(n_667), .Y(n_713) );
INVx1_ASAP7_75t_L g829 ( .A(n_665), .Y(n_829) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g707 ( .A(n_666), .Y(n_707) );
AND2x2_ASAP7_75t_L g759 ( .A(n_666), .B(n_746), .Y(n_759) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_691), .Y(n_669) );
OA222x2_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_676), .B1(n_681), .B2(n_682), .C1(n_685), .C2(n_688), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_672), .A2(n_845), .B(n_847), .Y(n_844) );
AND2x4_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
AND2x4_ASAP7_75t_L g683 ( .A(n_673), .B(n_684), .Y(n_683) );
NAND2x1_ASAP7_75t_L g706 ( .A(n_673), .B(n_707), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_673), .A2(n_792), .B(n_794), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_676), .A2(n_741), .B1(n_743), .B2(n_745), .Y(n_740) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_678), .B(n_709), .Y(n_708) );
INVx4_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g704 ( .A(n_684), .B(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_684), .A2(n_794), .B1(n_861), .B2(n_862), .Y(n_860) );
NOR2xp33_ASAP7_75t_SL g820 ( .A(n_685), .B(n_811), .Y(n_820) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2x1_ASAP7_75t_L g804 ( .A(n_686), .B(n_730), .Y(n_804) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_687), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g755 ( .A(n_687), .B(n_722), .Y(n_755) );
OR2x2_ASAP7_75t_L g776 ( .A(n_687), .B(n_722), .Y(n_776) );
INVx2_ASAP7_75t_L g769 ( .A(n_689), .Y(n_769) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI322xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_697), .A3(n_699), .B1(n_702), .B2(n_703), .C1(n_706), .C2(n_708), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g721 ( .A(n_696), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g831 ( .A(n_697), .B(n_832), .Y(n_831) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g757 ( .A(n_698), .B(n_701), .Y(n_757) );
AO221x1_ASAP7_75t_L g826 ( .A1(n_699), .A2(n_823), .B1(n_827), .B2(n_828), .C(n_830), .Y(n_826) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g812 ( .A(n_701), .B(n_769), .Y(n_812) );
AOI21xp5_ASAP7_75t_SL g736 ( .A1(n_703), .A2(n_731), .B(n_737), .Y(n_736) );
INVx4_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_704), .A2(n_750), .B1(n_820), .B2(n_821), .Y(n_819) );
AND2x2_ASAP7_75t_L g861 ( .A(n_707), .B(n_824), .Y(n_861) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_715), .A2(n_808), .B(n_812), .Y(n_807) );
INVx2_ASAP7_75t_L g817 ( .A(n_715), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_715), .A2(n_837), .B1(n_838), .B2(n_841), .Y(n_836) );
NOR3x1_ASAP7_75t_L g716 ( .A(n_717), .B(n_747), .C(n_770), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_735), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_724), .B1(n_730), .B2(n_733), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g766 ( .A(n_720), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_721), .B(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_721), .B(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_721), .B(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g780 ( .A(n_722), .Y(n_780) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_723), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_726), .B(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_727), .Y(n_846) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g832 ( .A(n_729), .Y(n_832) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_729), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_730), .B(n_775), .Y(n_774) );
INVx6_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g858 ( .A(n_732), .B(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_734), .B(n_800), .Y(n_818) );
NOR2xp67_ASAP7_75t_SL g735 ( .A(n_736), .B(n_740), .Y(n_735) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_756), .B(n_758), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_754), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g810 ( .A(n_751), .Y(n_810) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g761 ( .A(n_755), .Y(n_761) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_764), .B2(n_767), .Y(n_758) );
INVx2_ASAP7_75t_L g816 ( .A(n_759), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AO21x1_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_773), .B(n_777), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g837 ( .A(n_778), .Y(n_837) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
OR2x2_ASAP7_75t_L g848 ( .A(n_779), .B(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
BUFx2_ASAP7_75t_SL g803 ( .A(n_780), .Y(n_803) );
OR2x2_ASAP7_75t_L g802 ( .A(n_781), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g864 ( .A(n_781), .Y(n_864) );
NOR2x1_ASAP7_75t_L g783 ( .A(n_784), .B(n_813), .Y(n_783) );
NAND4xp75_ASAP7_75t_L g784 ( .A(n_785), .B(n_791), .C(n_797), .D(n_807), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B1(n_804), .B2(n_805), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_812), .A2(n_853), .B1(n_855), .B2(n_858), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_816), .B1(n_817), .B2(n_818), .C(n_819), .Y(n_813) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
AOI211x1_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_833), .B(n_835), .C(n_851), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g835 ( .A(n_836), .B(n_844), .Y(n_835) );
AND2x4_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
INVxp67_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_852), .B(n_860), .Y(n_851) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_863), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_870), .B(n_880), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_869), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_875), .B(n_879), .Y(n_870) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR2xp33_ASAP7_75t_R g880 ( .A(n_881), .B(n_882), .Y(n_880) );
BUFx3_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_886), .Y(n_893) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
endmodule