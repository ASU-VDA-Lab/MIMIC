module real_aes_2027_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_386;
wire n_905;
wire n_673;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_936;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_417;
wire n_449;
wire n_1006;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_727;
wire n_1014;
wire n_649;
wire n_385;
wire n_749;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_429;
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_0), .A2(n_317), .B1(n_639), .B2(n_640), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_1), .A2(n_209), .B1(n_647), .B2(n_741), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_2), .A2(n_267), .B1(n_455), .B2(n_517), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_3), .A2(n_113), .B1(n_438), .B2(n_523), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_4), .A2(n_119), .B1(n_429), .B2(n_690), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_5), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_6), .A2(n_190), .B1(n_483), .B2(n_557), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_7), .B(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_8), .A2(n_247), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_9), .A2(n_47), .B1(n_438), .B2(n_523), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_10), .A2(n_91), .B1(n_599), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_11), .A2(n_182), .B1(n_491), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_12), .A2(n_272), .B1(n_389), .B2(n_507), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_13), .A2(n_349), .B1(n_445), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_14), .A2(n_194), .B1(n_643), .B2(n_650), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_15), .A2(n_229), .B1(n_798), .B2(n_800), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_16), .A2(n_76), .B1(n_435), .B2(n_722), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_17), .A2(n_95), .B1(n_416), .B2(n_491), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_18), .A2(n_137), .B1(n_453), .B2(n_545), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_19), .A2(n_314), .B1(n_423), .B2(n_802), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_20), .A2(n_187), .B1(n_438), .B2(n_811), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_21), .A2(n_78), .B1(n_554), .B2(n_557), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_22), .A2(n_175), .B1(n_609), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_23), .A2(n_172), .B1(n_646), .B2(n_647), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_24), .A2(n_337), .B1(n_433), .B2(n_563), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_25), .A2(n_147), .B1(n_447), .B2(n_478), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_26), .A2(n_60), .B1(n_517), .B2(n_545), .Y(n_963) );
XOR2x2_ASAP7_75t_L g906 ( .A(n_27), .B(n_907), .Y(n_906) );
AO222x2_ASAP7_75t_L g776 ( .A1(n_28), .A2(n_142), .B1(n_231), .B2(n_626), .C1(n_634), .C2(n_729), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_29), .A2(n_323), .B1(n_631), .B2(n_732), .Y(n_779) );
INVx1_ASAP7_75t_SL g399 ( .A(n_30), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_30), .B(n_40), .Y(n_988) );
OA22x2_ASAP7_75t_L g383 ( .A1(n_31), .A2(n_384), .B1(n_385), .B2(n_386), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_31), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_32), .A2(n_169), .B1(n_618), .B2(n_766), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_33), .A2(n_364), .B1(n_429), .B2(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_34), .B(n_475), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_35), .A2(n_280), .B1(n_643), .B2(n_650), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_36), .A2(n_114), .B1(n_631), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_37), .A2(n_181), .B1(n_867), .B2(n_965), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_38), .A2(n_354), .B1(n_445), .B2(n_447), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_39), .A2(n_316), .B1(n_416), .B2(n_487), .Y(n_571) );
AO22x2_ASAP7_75t_L g393 ( .A1(n_40), .A2(n_344), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_41), .A2(n_203), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_42), .A2(n_109), .B1(n_429), .B2(n_433), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_43), .A2(n_52), .B1(n_455), .B2(n_517), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_44), .A2(n_357), .B1(n_416), .B2(n_615), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_45), .A2(n_176), .B1(n_523), .B2(n_533), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_46), .A2(n_273), .B1(n_416), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_48), .A2(n_327), .B1(n_423), .B2(n_484), .Y(n_767) );
INVx1_ASAP7_75t_L g400 ( .A(n_49), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_50), .A2(n_300), .B1(n_649), .B2(n_650), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_51), .A2(n_235), .B1(n_416), .B2(n_618), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_53), .A2(n_287), .B1(n_478), .B2(n_795), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_54), .A2(n_285), .B1(n_423), .B2(n_512), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_55), .A2(n_296), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_56), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_57), .A2(n_127), .B1(n_574), .B2(n_802), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_58), .A2(n_341), .B1(n_889), .B2(n_890), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_59), .A2(n_292), .B1(n_419), .B2(n_661), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_61), .A2(n_241), .B1(n_438), .B2(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_62), .A2(n_205), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_63), .A2(n_331), .B1(n_423), .B2(n_425), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_64), .B(n_475), .Y(n_949) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_65), .A2(n_188), .B1(n_394), .B2(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_66), .A2(n_192), .B1(n_609), .B2(n_611), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_67), .A2(n_81), .B1(n_611), .B2(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_68), .A2(n_301), .B1(n_507), .B2(n_609), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_69), .A2(n_228), .B1(n_423), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_70), .A2(n_138), .B1(n_650), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_71), .A2(n_338), .B1(n_453), .B2(n_455), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_72), .A2(n_161), .B1(n_627), .B2(n_867), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_73), .A2(n_193), .B1(n_416), .B2(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_74), .A2(n_153), .B1(n_560), .B2(n_662), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_75), .A2(n_111), .B1(n_639), .B2(n_640), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_77), .A2(n_277), .B1(n_642), .B2(n_646), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_79), .A2(n_248), .B1(n_519), .B2(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_80), .A2(n_244), .B1(n_634), .B2(n_635), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_82), .B(n_666), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_83), .A2(n_189), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_84), .A2(n_227), .B1(n_419), .B2(n_506), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_85), .A2(n_355), .B1(n_438), .B2(n_523), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_86), .A2(n_293), .B1(n_445), .B2(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_87), .A2(n_269), .B1(n_484), .B2(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_88), .A2(n_133), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_89), .A2(n_312), .B1(n_447), .B2(n_548), .Y(n_547) );
AO222x2_ASAP7_75t_L g625 ( .A1(n_90), .A2(n_202), .B1(n_347), .B2(n_626), .C1(n_627), .C2(n_628), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_92), .A2(n_123), .B1(n_997), .B2(n_999), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_93), .A2(n_222), .B1(n_599), .B2(n_628), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_94), .A2(n_224), .B1(n_440), .B2(n_533), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_96), .A2(n_246), .B1(n_419), .B2(n_722), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_97), .A2(n_250), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_98), .A2(n_170), .B1(n_329), .B2(n_460), .C1(n_521), .C2(n_523), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_99), .Y(n_848) );
OA22x2_ASAP7_75t_L g817 ( .A1(n_100), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_100), .Y(n_818) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_101), .A2(n_139), .B1(n_265), .B2(n_460), .C1(n_478), .C2(n_479), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_102), .A2(n_155), .B1(n_627), .B2(n_632), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_103), .A2(n_261), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_104), .A2(n_226), .B1(n_574), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_105), .A2(n_120), .B1(n_563), .B2(n_917), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_106), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_107), .A2(n_230), .B1(n_423), .B2(n_425), .Y(n_422) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_108), .A2(n_276), .B1(n_394), .B2(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_110), .A2(n_291), .B1(n_447), .B2(n_683), .Y(n_682) );
OAI22x1_ASAP7_75t_L g960 ( .A1(n_112), .A2(n_961), .B1(n_975), .B2(n_976), .Y(n_960) );
CKINVDCx16_ASAP7_75t_R g976 ( .A(n_112), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_115), .A2(n_151), .B1(n_479), .B2(n_683), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_116), .A2(n_257), .B1(n_429), .B2(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_117), .A2(n_141), .B1(n_389), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_118), .A2(n_236), .B1(n_470), .B2(n_471), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_121), .A2(n_239), .B1(n_487), .B2(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g524 ( .A(n_122), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_124), .A2(n_336), .B1(n_640), .B2(n_737), .Y(n_736) );
OA22x2_ASAP7_75t_L g697 ( .A1(n_125), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_125), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_126), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_128), .A2(n_196), .B1(n_647), .B2(n_741), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_129), .A2(n_321), .B1(n_808), .B2(n_810), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_130), .B(n_475), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_131), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_132), .A2(n_221), .B1(n_453), .B2(n_455), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_134), .A2(n_225), .B1(n_435), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_135), .A2(n_166), .B1(n_719), .B2(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_136), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_140), .A2(n_313), .B1(n_506), .B2(n_618), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_143), .A2(n_164), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_144), .A2(n_152), .B1(n_642), .B2(n_646), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_145), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_146), .A2(n_320), .B1(n_470), .B2(n_471), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_148), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_149), .A2(n_214), .B1(n_506), .B2(n_509), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_150), .A2(n_234), .B1(n_438), .B2(n_440), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_154), .A2(n_211), .B1(n_509), .B2(n_969), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_156), .A2(n_363), .B1(n_487), .B2(n_552), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_157), .B(n_666), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_158), .A2(n_232), .B1(n_389), .B2(n_408), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_159), .A2(n_278), .B1(n_425), .B2(n_483), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_160), .A2(n_351), .B1(n_519), .B2(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_162), .B(n_536), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_163), .A2(n_332), .B1(n_478), .B2(n_580), .Y(n_910) );
OA22x2_ASAP7_75t_L g755 ( .A1(n_165), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_165), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_167), .A2(n_340), .B1(n_560), .B2(n_561), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_168), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_171), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_173), .A2(n_219), .B1(n_453), .B2(n_455), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_174), .A2(n_330), .B1(n_661), .B2(n_662), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_177), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_178), .A2(n_199), .B1(n_470), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_179), .A2(n_288), .B1(n_791), .B2(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_180), .A2(n_251), .B1(n_455), .B2(n_517), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_183), .A2(n_352), .B1(n_438), .B2(n_523), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_184), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_185), .A2(n_366), .B1(n_692), .B2(n_766), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_186), .A2(n_302), .B1(n_609), .B2(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g987 ( .A(n_188), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_191), .A2(n_220), .B1(n_643), .B2(n_650), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_195), .A2(n_345), .B1(n_517), .B2(n_545), .Y(n_883) );
INVx1_ASAP7_75t_L g1006 ( .A(n_197), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_198), .A2(n_309), .B1(n_631), .B2(n_632), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_200), .A2(n_946), .B1(n_947), .B2(n_958), .Y(n_945) );
INVxp67_ASAP7_75t_L g958 ( .A(n_200), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_201), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_204), .A2(n_258), .B1(n_438), .B2(n_440), .Y(n_437) );
OA22x2_ASAP7_75t_L g566 ( .A1(n_206), .A2(n_567), .B1(n_568), .B2(n_583), .Y(n_566) );
INVxp67_ASAP7_75t_L g583 ( .A(n_206), .Y(n_583) );
OA22x2_ASAP7_75t_L g585 ( .A1(n_206), .A2(n_567), .B1(n_568), .B2(n_583), .Y(n_585) );
XNOR2x1_ASAP7_75t_L g590 ( .A(n_207), .B(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_208), .A2(n_359), .B1(n_438), .B2(n_440), .Y(n_761) );
INVx2_ASAP7_75t_L g375 ( .A(n_210), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_212), .A2(n_356), .B1(n_647), .B2(n_649), .Y(n_785) );
OA22x2_ASAP7_75t_L g463 ( .A1(n_213), .A2(n_464), .B1(n_496), .B2(n_497), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_213), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_215), .A2(n_262), .B1(n_429), .B2(n_611), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_216), .A2(n_237), .B1(n_490), .B2(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_217), .A2(n_991), .B1(n_1011), .B2(n_1012), .Y(n_990) );
INVx1_ASAP7_75t_L g1011 ( .A(n_217), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_218), .A2(n_245), .B1(n_453), .B2(n_470), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_223), .A2(n_307), .B1(n_507), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_233), .A2(n_271), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_238), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_240), .A2(n_992), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_240), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_242), .A2(n_622), .B1(n_623), .B2(n_651), .Y(n_621) );
INVx1_ASAP7_75t_L g651 ( .A(n_242), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_243), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_249), .A2(n_324), .B1(n_634), .B2(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_252), .A2(n_259), .B1(n_438), .B2(n_523), .Y(n_929) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_253), .A2(n_368), .B(n_376), .C(n_989), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_254), .A2(n_274), .B1(n_627), .B2(n_632), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_255), .A2(n_335), .B1(n_416), .B2(n_419), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_256), .A2(n_289), .B1(n_523), .B2(n_533), .Y(n_880) );
XNOR2x1_ASAP7_75t_L g923 ( .A(n_260), .B(n_924), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_263), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_264), .A2(n_343), .B1(n_419), .B2(n_661), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_266), .A2(n_339), .B1(n_483), .B2(n_573), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_268), .B(n_475), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_270), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_275), .A2(n_319), .B1(n_389), .B2(n_618), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_276), .B(n_986), .Y(n_985) );
AOI222xp33_ASAP7_75t_L g973 ( .A1(n_279), .A2(n_290), .B1(n_325), .B2(n_626), .C1(n_729), .C2(n_974), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_281), .A2(n_328), .B1(n_647), .B2(n_649), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_282), .B(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_283), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_284), .A2(n_365), .B1(n_423), .B2(n_573), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_286), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_294), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_295), .A2(n_310), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_297), .A2(n_318), .B1(n_429), .B2(n_433), .Y(n_768) );
INVx1_ASAP7_75t_L g564 ( .A(n_298), .Y(n_564) );
INVx3_ASAP7_75t_L g394 ( .A(n_299), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_303), .A2(n_311), .B1(n_647), .B2(n_649), .Y(n_873) );
AOI222xp33_ASAP7_75t_L g807 ( .A1(n_304), .A2(n_342), .B1(n_350), .B2(n_475), .C1(n_808), .C2(n_810), .Y(n_807) );
OAI22x1_ASAP7_75t_L g678 ( .A1(n_305), .A2(n_679), .B1(n_693), .B2(n_694), .Y(n_678) );
INVx1_ASAP7_75t_L g694 ( .A(n_305), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_306), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_308), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_315), .Y(n_895) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_322), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_326), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_333), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_334), .A2(n_362), .B1(n_478), .B2(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_346), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g983 ( .A(n_346), .Y(n_983) );
INVx1_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
AND2x2_ASAP7_75t_R g1014 ( .A(n_348), .B(n_983), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_353), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_358), .B(n_626), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_360), .B(n_666), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_361), .Y(n_600) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_371), .B(n_373), .Y(n_1023) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_372), .B(n_983), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_749), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_376) );
INVx1_ASAP7_75t_L g978 ( .A(n_377), .Y(n_978) );
OAI22xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_586), .B1(n_587), .B2(n_748), .Y(n_377) );
INVx1_ASAP7_75t_L g748 ( .A(n_378), .Y(n_748) );
OA22x2_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_525), .B2(n_526), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OA22x2_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_501), .B2(n_502), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_463), .B1(n_499), .B2(n_500), .Y(n_382) );
INVx1_ASAP7_75t_L g499 ( .A(n_383), .Y(n_499) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_436), .Y(n_386) );
NAND4xp25_ASAP7_75t_L g387 ( .A(n_388), .B(n_415), .C(n_422), .D(n_428), .Y(n_387) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g493 ( .A(n_390), .Y(n_493) );
INVx2_ASAP7_75t_L g506 ( .A(n_390), .Y(n_506) );
INVx2_ASAP7_75t_SL g766 ( .A(n_390), .Y(n_766) );
INVx3_ASAP7_75t_L g889 ( .A(n_390), .Y(n_889) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g552 ( .A(n_391), .Y(n_552) );
BUFx2_ASAP7_75t_L g969 ( .A(n_391), .Y(n_969) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_401), .Y(n_391) );
AND2x2_ASAP7_75t_L g424 ( .A(n_392), .B(n_413), .Y(n_424) );
AND2x4_ASAP7_75t_L g446 ( .A(n_392), .B(n_421), .Y(n_446) );
AND2x2_ASAP7_75t_L g632 ( .A(n_392), .B(n_421), .Y(n_632) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_392), .B(n_413), .Y(n_639) );
AND2x6_ASAP7_75t_L g643 ( .A(n_392), .B(n_401), .Y(n_643) );
AND2x2_ASAP7_75t_L g737 ( .A(n_392), .B(n_413), .Y(n_737) );
AND2x2_ASAP7_75t_L g867 ( .A(n_392), .B(n_421), .Y(n_867) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
INVx2_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
BUFx2_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
AND2x2_ASAP7_75t_L g451 ( .A(n_393), .B(n_397), .Y(n_451) );
INVx1_ASAP7_75t_L g395 ( .A(n_394), .Y(n_395) );
OAI22x1_ASAP7_75t_L g397 ( .A1(n_394), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_394), .Y(n_398) );
INVx2_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_394), .Y(n_407) );
AND2x4_ASAP7_75t_L g411 ( .A(n_396), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_412), .Y(n_432) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
AND2x4_ASAP7_75t_L g418 ( .A(n_401), .B(n_411), .Y(n_418) );
AND2x4_ASAP7_75t_L g431 ( .A(n_401), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_451), .Y(n_462) );
AND2x4_ASAP7_75t_L g626 ( .A(n_401), .B(n_451), .Y(n_626) );
AND2x2_ASAP7_75t_L g642 ( .A(n_401), .B(n_411), .Y(n_642) );
AND2x2_ASAP7_75t_L g649 ( .A(n_401), .B(n_432), .Y(n_649) );
AND2x2_ASAP7_75t_L g741 ( .A(n_401), .B(n_432), .Y(n_741) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g414 ( .A(n_403), .Y(n_414) );
AND2x4_ASAP7_75t_L g421 ( .A(n_403), .B(n_405), .Y(n_421) );
AND2x2_ASAP7_75t_L g427 ( .A(n_403), .B(n_406), .Y(n_427) );
INVxp67_ASAP7_75t_L g450 ( .A(n_405), .Y(n_450) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g413 ( .A(n_406), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g487 ( .A(n_409), .Y(n_487) );
INVx2_ASAP7_75t_L g509 ( .A(n_409), .Y(n_509) );
INVx2_ASAP7_75t_SL g618 ( .A(n_409), .Y(n_618) );
INVx2_ASAP7_75t_L g692 ( .A(n_409), .Y(n_692) );
INVx2_ASAP7_75t_SL g890 ( .A(n_409), .Y(n_890) );
INVx8_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x4_ASAP7_75t_L g420 ( .A(n_411), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g435 ( .A(n_411), .B(n_427), .Y(n_435) );
AND2x2_ASAP7_75t_L g646 ( .A(n_411), .B(n_421), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_411), .B(n_427), .Y(n_647) );
AND2x6_ASAP7_75t_L g650 ( .A(n_411), .B(n_413), .Y(n_650) );
AND2x2_ASAP7_75t_L g454 ( .A(n_413), .B(n_432), .Y(n_454) );
AND2x4_ASAP7_75t_L g631 ( .A(n_413), .B(n_432), .Y(n_631) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_414), .Y(n_458) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx3_ASAP7_75t_SL g560 ( .A(n_417), .Y(n_560) );
INVx4_ASAP7_75t_L g610 ( .A(n_417), .Y(n_610) );
INVx2_ASAP7_75t_L g661 ( .A(n_417), .Y(n_661) );
INVx2_ASAP7_75t_SL g719 ( .A(n_417), .Y(n_719) );
INVx8_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_419), .Y(n_561) );
INVx1_ASAP7_75t_L g616 ( .A(n_419), .Y(n_616) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g495 ( .A(n_420), .Y(n_495) );
BUFx3_ASAP7_75t_L g507 ( .A(n_420), .Y(n_507) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_420), .Y(n_662) );
AND2x2_ASAP7_75t_L g439 ( .A(n_421), .B(n_432), .Y(n_439) );
AND2x4_ASAP7_75t_L g634 ( .A(n_421), .B(n_432), .Y(n_634) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
INVx2_ASAP7_75t_L g556 ( .A(n_424), .Y(n_556) );
INVx5_ASAP7_75t_SL g485 ( .A(n_425), .Y(n_485) );
BUFx3_ASAP7_75t_L g557 ( .A(n_425), .Y(n_557) );
BUFx2_ASAP7_75t_L g573 ( .A(n_425), .Y(n_573) );
BUFx2_ASAP7_75t_L g802 ( .A(n_425), .Y(n_802) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x4_ASAP7_75t_L g640 ( .A(n_426), .B(n_427), .Y(n_640) );
AND2x2_ASAP7_75t_L g442 ( .A(n_427), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_427), .B(n_443), .Y(n_635) );
AND2x2_ASAP7_75t_SL g729 ( .A(n_427), .B(n_443), .Y(n_729) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
INVx3_ASAP7_75t_L g563 ( .A(n_430), .Y(n_563) );
INVx2_ASAP7_75t_L g806 ( .A(n_430), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_430), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
INVx6_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g722 ( .A(n_431), .Y(n_722) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g917 ( .A(n_434), .Y(n_917) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g491 ( .A(n_435), .Y(n_491) );
BUFx3_ASAP7_75t_L g514 ( .A(n_435), .Y(n_514) );
BUFx2_ASAP7_75t_SL g611 ( .A(n_435), .Y(n_611) );
BUFx2_ASAP7_75t_SL g690 ( .A(n_435), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_437), .B(n_444), .C(n_452), .D(n_459), .Y(n_436) );
BUFx5_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
BUFx3_ASAP7_75t_L g809 ( .A(n_439), .Y(n_809) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g468 ( .A(n_441), .Y(n_468) );
INVx3_ASAP7_75t_L g811 ( .A(n_441), .Y(n_811) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx12f_ASAP7_75t_L g523 ( .A(n_442), .Y(n_523) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_446), .Y(n_548) );
BUFx2_ASAP7_75t_L g669 ( .A(n_446), .Y(n_669) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g479 ( .A(n_448), .Y(n_479) );
INVx2_ASAP7_75t_L g519 ( .A(n_448), .Y(n_519) );
INVx1_ASAP7_75t_L g580 ( .A(n_448), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_448), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_448), .A2(n_604), .B1(n_711), .B2(n_712), .Y(n_710) );
INVx2_ASAP7_75t_L g795 ( .A(n_448), .Y(n_795) );
INVx2_ASAP7_75t_L g885 ( .A(n_448), .Y(n_885) );
INVx6_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AND2x2_ASAP7_75t_L g627 ( .A(n_450), .B(n_451), .Y(n_627) );
AND2x2_ASAP7_75t_L g965 ( .A(n_450), .B(n_451), .Y(n_965) );
AND2x4_ASAP7_75t_L g456 ( .A(n_451), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g628 ( .A(n_451), .B(n_457), .Y(n_628) );
AND2x2_ASAP7_75t_L g732 ( .A(n_451), .B(n_457), .Y(n_732) );
INVx1_ASAP7_75t_L g707 ( .A(n_453), .Y(n_707) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g472 ( .A(n_454), .Y(n_472) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_454), .Y(n_517) );
INVxp67_ASAP7_75t_L g601 ( .A(n_455), .Y(n_601) );
BUFx4f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_SL g470 ( .A(n_456), .Y(n_470) );
INVx2_ASAP7_75t_L g546 ( .A(n_456), .Y(n_546) );
BUFx3_ASAP7_75t_L g792 ( .A(n_456), .Y(n_792) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g927 ( .A(n_460), .Y(n_927) );
INVx4_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g475 ( .A(n_461), .Y(n_475) );
INVx3_ASAP7_75t_SL g537 ( .A(n_461), .Y(n_537) );
INVx3_ASAP7_75t_L g666 ( .A(n_461), .Y(n_666) );
INVx4_ASAP7_75t_SL g862 ( .A(n_461), .Y(n_862) );
INVx6_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_480), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_473), .C(n_476), .Y(n_465) );
NOR4xp25_ASAP7_75t_L g497 ( .A(n_466), .B(n_481), .C(n_488), .D(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVxp67_ASAP7_75t_L g709 ( .A(n_470), .Y(n_709) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx4_ASAP7_75t_L g599 ( .A(n_472), .Y(n_599) );
INVx1_ASAP7_75t_L g828 ( .A(n_472), .Y(n_828) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_474), .B(n_477), .Y(n_498) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_488), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_486), .Y(n_481) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g512 ( .A(n_485), .Y(n_512) );
OAI22xp33_ASAP7_75t_SL g849 ( .A1(n_485), .A2(n_850), .B1(n_853), .B2(n_854), .Y(n_849) );
INVx2_ASAP7_75t_L g999 ( .A(n_485), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
BUFx2_ASAP7_75t_L g845 ( .A(n_493), .Y(n_845) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g720 ( .A(n_495), .Y(n_720) );
INVx1_ASAP7_75t_L g1002 ( .A(n_495), .Y(n_1002) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
XOR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_524), .Y(n_502) );
NAND4xp75_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .C(n_515), .D(n_520), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
BUFx6f_ASAP7_75t_SL g544 ( .A(n_517), .Y(n_544) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g533 ( .A(n_522), .Y(n_533) );
BUFx3_ASAP7_75t_L g540 ( .A(n_523), .Y(n_540) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_565), .B1(n_584), .B2(n_585), .Y(n_526) );
INVx3_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
XOR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_564), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_549), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_542), .Y(n_529) );
OAI222xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_534), .B1(n_535), .B2(n_538), .C1(n_539), .C2(n_541), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g822 ( .A1(n_535), .A2(n_823), .B(n_824), .Y(n_822) );
OAI21xp33_ASAP7_75t_L g1005 ( .A1(n_535), .A2(n_1006), .B(n_1007), .Y(n_1005) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g604 ( .A(n_548), .Y(n_604) );
BUFx4f_ASAP7_75t_SL g683 ( .A(n_548), .Y(n_683) );
BUFx2_ASAP7_75t_L g794 ( .A(n_548), .Y(n_794) );
BUFx2_ASAP7_75t_L g830 ( .A(n_548), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g575 ( .A(n_556), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_577), .Y(n_568) );
NAND4xp25_ASAP7_75t_SL g569 ( .A(n_570), .B(n_571), .C(n_572), .D(n_576), .Y(n_569) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g852 ( .A(n_575), .Y(n_852) );
INVx1_ASAP7_75t_L g998 ( .A(n_575), .Y(n_998) );
NAND4xp25_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .C(n_581), .D(n_582), .Y(n_577) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_674), .B2(n_747), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_619), .B1(n_671), .B2(n_672), .Y(n_589) );
INVx1_ASAP7_75t_L g671 ( .A(n_590), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_606), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .C(n_602), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_600), .B2(n_601), .Y(n_596) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g799 ( .A(n_610), .Y(n_799) );
INVx1_ASAP7_75t_L g841 ( .A(n_611), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g673 ( .A(n_619), .Y(n_673) );
OA22x2_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_652), .B2(n_653), .Y(n_619) );
AO22x2_ASAP7_75t_L g904 ( .A1(n_620), .A2(n_905), .B1(n_906), .B2(n_919), .Y(n_904) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g919 ( .A(n_621), .Y(n_919) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_636), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_633), .Y(n_629) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_634), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_644), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_664), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .C(n_660), .D(n_663), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_662), .Y(n_800) );
INVx2_ASAP7_75t_L g835 ( .A(n_662), .Y(n_835) );
NAND4xp25_ASAP7_75t_SL g664 ( .A(n_665), .B(n_667), .C(n_668), .D(n_670), .Y(n_664) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g747 ( .A(n_674), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_695), .B2(n_746), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g693 ( .A(n_679), .Y(n_693) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_686), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .C(n_684), .D(n_685), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .C(n_689), .D(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g847 ( .A(n_692), .Y(n_847) );
INVx1_ASAP7_75t_L g746 ( .A(n_695), .Y(n_746) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AO22x2_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_723), .B1(n_744), .B2(n_745), .Y(n_696) );
INVx1_ASAP7_75t_L g744 ( .A(n_697), .Y(n_744) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_713), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .C(n_710), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .Y(n_717) );
BUFx2_ASAP7_75t_L g839 ( .A(n_719), .Y(n_839) );
INVx1_ASAP7_75t_L g745 ( .A(n_723), .Y(n_745) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_723), .B(n_755), .Y(n_754) );
XOR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_743), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_725), .B(n_734), .Y(n_724) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_730), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_739), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g979 ( .A(n_749), .Y(n_979) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_901), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_814), .B(n_899), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_751), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
XNOR2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_769), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_763), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .C(n_762), .Y(n_759) );
NAND4xp25_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .C(n_767), .D(n_768), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_787), .B2(n_813), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
XNOR2x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_780), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx2_ASAP7_75t_SL g813 ( .A(n_787), .Y(n_813) );
XNOR2x1_ASAP7_75t_L g787 ( .A(n_788), .B(n_812), .Y(n_787) );
NAND4xp75_ASAP7_75t_L g788 ( .A(n_789), .B(n_796), .C(n_803), .D(n_807), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_793), .Y(n_789) );
BUFx6f_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
BUFx6f_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g900 ( .A(n_815), .Y(n_900) );
OAI22x1_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_855), .B1(n_856), .B2(n_898), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g898 ( .A(n_817), .Y(n_898) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AND3x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_831), .C(n_842), .Y(n_820) );
NOR2xp67_ASAP7_75t_SL g821 ( .A(n_822), .B(n_825), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_826), .B(n_829), .Y(n_825) );
BUFx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_836), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_840), .B2(n_841), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_849), .Y(n_842) );
OAI22xp33_ASAP7_75t_SL g843 ( .A1(n_844), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g936 ( .A(n_852), .Y(n_936) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AO22x2_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_876), .B1(n_896), .B2(n_897), .Y(n_856) );
INVx1_ASAP7_75t_SL g897 ( .A(n_857), .Y(n_897) );
XOR2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_875), .Y(n_857) );
NAND2xp5_ASAP7_75t_SL g858 ( .A(n_859), .B(n_868), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_864), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx2_ASAP7_75t_L g896 ( .A(n_876), .Y(n_896) );
XOR2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_895), .Y(n_876) );
NAND2x1p5_ASAP7_75t_L g877 ( .A(n_878), .B(n_886), .Y(n_877) );
NOR2x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_882), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NOR2x1_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
OAI22xp5_ASAP7_75t_SL g901 ( .A1(n_902), .A2(n_942), .B1(n_943), .B2(n_977), .Y(n_901) );
INVx1_ASAP7_75t_L g977 ( .A(n_902), .Y(n_977) );
OAI22xp5_ASAP7_75t_SL g902 ( .A1(n_903), .A2(n_904), .B1(n_920), .B2(n_941), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NOR2xp67_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .Y(n_907) );
NAND4xp25_ASAP7_75t_SL g908 ( .A(n_909), .B(n_910), .C(n_911), .D(n_912), .Y(n_908) );
NAND4xp25_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .C(n_916), .D(n_918), .Y(n_913) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g941 ( .A(n_922), .Y(n_941) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AND2x4_ASAP7_75t_L g924 ( .A(n_925), .B(n_933), .Y(n_924) );
NOR2xp67_ASAP7_75t_L g925 ( .A(n_926), .B(n_930), .Y(n_925) );
OAI21xp5_ASAP7_75t_SL g926 ( .A1(n_927), .A2(n_928), .B(n_929), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
NOR2x1_ASAP7_75t_L g933 ( .A(n_934), .B(n_938), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_937), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OA22x2_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_945), .B1(n_959), .B2(n_960), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NOR2xp67_ASAP7_75t_L g947 ( .A(n_948), .B(n_953), .Y(n_947) );
NAND4xp25_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .C(n_951), .D(n_952), .Y(n_948) );
NAND4xp25_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .C(n_956), .D(n_957), .Y(n_953) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND4xp25_ASAP7_75t_SL g961 ( .A(n_962), .B(n_966), .C(n_970), .D(n_973), .Y(n_961) );
AND4x1_ASAP7_75t_L g975 ( .A(n_962), .B(n_966), .C(n_970), .D(n_973), .Y(n_975) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_964), .Y(n_962) );
AND2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
AND2x2_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
INVx4_ASAP7_75t_R g980 ( .A(n_981), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_982), .B(n_985), .Y(n_1022) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
OAI222xp33_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_1013), .B1(n_1015), .B2(n_1018), .C1(n_1020), .C2(n_1023), .Y(n_989) );
CKINVDCx16_ASAP7_75t_R g1012 ( .A(n_991), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_SL g1019 ( .A(n_992), .Y(n_1019) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_1004), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_994), .B(n_1000), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1003), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1008), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
INVx1_ASAP7_75t_SL g1013 ( .A(n_1014), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVxp33_ASAP7_75t_SL g1016 ( .A(n_1017), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_1021), .Y(n_1020) );
CKINVDCx6p67_ASAP7_75t_R g1021 ( .A(n_1022), .Y(n_1021) );
endmodule