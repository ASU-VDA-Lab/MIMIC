module fake_jpeg_14441_n_584 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_584);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_59),
.Y(n_121)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_22),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_60),
.B(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_89),
.Y(n_133)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_78),
.Y(n_190)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_8),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_30),
.B(n_10),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_10),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_30),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_105),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_51),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_37),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_20),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_33),
.B(n_16),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_110),
.A2(n_43),
.B(n_33),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_116),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_36),
.B1(n_54),
.B2(n_28),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_124),
.A2(n_155),
.B1(n_184),
.B2(n_164),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_125),
.B(n_154),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_23),
.B1(n_29),
.B2(n_34),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_134),
.A2(n_165),
.B1(n_168),
.B2(n_71),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_38),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_152),
.B(n_174),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_87),
.B(n_51),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_99),
.A2(n_102),
.B1(n_101),
.B2(n_119),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_37),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_161),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_56),
.B(n_37),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_69),
.A2(n_28),
.B1(n_54),
.B2(n_35),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_164),
.A2(n_51),
.B(n_110),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_38),
.B1(n_34),
.B2(n_29),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_120),
.B1(n_70),
.B2(n_98),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_43),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_181),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_55),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_13),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_90),
.B(n_50),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_SL g183 ( 
.A(n_58),
.Y(n_183)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_61),
.A2(n_28),
.B1(n_54),
.B2(n_35),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_94),
.B(n_50),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_50),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_170),
.Y(n_197)
);

BUFx24_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_125),
.A2(n_154),
.B1(n_128),
.B2(n_161),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_198),
.Y(n_313)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_35),
.B1(n_112),
.B2(n_74),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_200),
.A2(n_244),
.B1(n_259),
.B2(n_260),
.Y(n_286)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_201),
.Y(n_303)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_203),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_256),
.B1(n_182),
.B2(n_126),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_124),
.A2(n_63),
.B1(n_107),
.B2(n_93),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_207),
.A2(n_210),
.B1(n_225),
.B2(n_188),
.Y(n_295)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_208),
.Y(n_267)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_209),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_83),
.B1(n_82),
.B2(n_77),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

BUFx4f_ASAP7_75t_SL g291 ( 
.A(n_213),
.Y(n_291)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_158),
.A2(n_79),
.B1(n_116),
.B2(n_50),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_216),
.B(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_41),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_217),
.B(n_238),
.Y(n_293)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_152),
.A2(n_73),
.B(n_78),
.C(n_81),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_50),
.B1(n_55),
.B2(n_39),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_224),
.A2(n_250),
.B1(n_262),
.B2(n_144),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_39),
.B1(n_41),
.B2(n_113),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_229),
.Y(n_269)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_191),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_232),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_195),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_234),
.Y(n_270)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_139),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_240),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_121),
.B(n_16),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_72),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_142),
.B(n_106),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_245),
.Y(n_280)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g278 ( 
.A(n_242),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_174),
.B(n_86),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_248),
.B(n_253),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_0),
.Y(n_284)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_145),
.B(n_71),
.Y(n_253)
);

AO22x2_ASAP7_75t_SL g254 ( 
.A1(n_184),
.A2(n_75),
.B1(n_100),
.B2(n_2),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_254),
.A2(n_149),
.B1(n_126),
.B2(n_132),
.Y(n_299)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_169),
.A2(n_27),
.B1(n_20),
.B2(n_75),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_153),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_257),
.Y(n_300)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_172),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_258),
.Y(n_317)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_122),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_261),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_136),
.A2(n_176),
.B1(n_189),
.B2(n_169),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_167),
.B(n_27),
.C(n_20),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_150),
.C(n_180),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_16),
.B(n_14),
.C(n_12),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_11),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_27),
.B1(n_14),
.B2(n_12),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_177),
.B1(n_144),
.B2(n_182),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_266),
.B(n_222),
.C(n_214),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_288),
.B1(n_295),
.B2(n_316),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_272),
.A2(n_273),
.B1(n_301),
.B2(n_305),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_275),
.A2(n_296),
.B(n_240),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_189),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_289),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_198),
.B(n_11),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_283),
.B(n_265),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_284),
.B(n_5),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_246),
.A2(n_180),
.B1(n_188),
.B2(n_185),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_160),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_228),
.A2(n_185),
.B1(n_160),
.B2(n_149),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_299),
.A2(n_253),
.B1(n_230),
.B2(n_220),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_254),
.A2(n_190),
.B1(n_132),
.B2(n_27),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_254),
.A2(n_190),
.B1(n_11),
.B2(n_2),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_204),
.B(n_0),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_284),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_207),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_319),
.A2(n_229),
.B1(n_234),
.B2(n_231),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_270),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_337),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_326),
.B(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_289),
.B(n_221),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_342),
.Y(n_370)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_228),
.B(n_235),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_335),
.A2(n_351),
.B(n_277),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_336),
.A2(n_338),
.B1(n_346),
.B2(n_357),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_295),
.A2(n_235),
.B1(n_232),
.B2(n_223),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_264),
.B(n_200),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_339),
.A2(n_272),
.B(n_286),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_340),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_265),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_278),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_277),
.A2(n_211),
.B1(n_239),
.B2(n_213),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_344),
.A2(n_361),
.B1(n_307),
.B2(n_282),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_308),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_345),
.B(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_307),
.Y(n_347)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_263),
.C(n_215),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_355),
.C(n_302),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_275),
.A2(n_224),
.B(n_262),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_243),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g353 ( 
.A1(n_301),
.A2(n_225),
.B1(n_203),
.B2(n_258),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_299),
.A2(n_252),
.B1(n_242),
.B2(n_219),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_273),
.A2(n_260),
.B1(n_202),
.B2(n_206),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_358),
.A2(n_319),
.B1(n_279),
.B2(n_297),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_300),
.B(n_11),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_6),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_282),
.Y(n_385)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_206),
.B1(n_227),
.B2(n_6),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_362),
.A2(n_307),
.B1(n_309),
.B2(n_267),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_316),
.B1(n_281),
.B2(n_266),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_367),
.A2(n_383),
.B1(n_397),
.B2(n_338),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_349),
.C(n_325),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_374),
.B(n_389),
.Y(n_412)
);

AO32x1_ASAP7_75t_L g374 ( 
.A1(n_335),
.A2(n_283),
.A3(n_302),
.B1(n_307),
.B2(n_297),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_297),
.B1(n_296),
.B2(n_317),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_385),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_390),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_339),
.A2(n_280),
.B(n_274),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_317),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_331),
.Y(n_392)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_274),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_398),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_394),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_332),
.A2(n_285),
.B1(n_298),
.B2(n_304),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_395),
.A2(n_344),
.B1(n_347),
.B2(n_340),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_293),
.B1(n_306),
.B2(n_267),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_306),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_345),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_374),
.C(n_373),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_390),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_401),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_385),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_355),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_411),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_421),
.B1(n_423),
.B2(n_426),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_410),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_393),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_349),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_413),
.A2(n_384),
.B1(n_386),
.B2(n_343),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_330),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_391),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_419),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_371),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_422),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_367),
.A2(n_321),
.B1(n_341),
.B2(n_346),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_381),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_380),
.A2(n_321),
.B1(n_336),
.B2(n_357),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_379),
.B(n_360),
.Y(n_424)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_424),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_389),
.A2(n_323),
.B(n_351),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_380),
.A2(n_353),
.B1(n_362),
.B2(n_358),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_359),
.Y(n_428)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_379),
.B(n_352),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_431),
.Y(n_459)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_371),
.A2(n_353),
.A3(n_350),
.B1(n_348),
.B2(n_333),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_436),
.B1(n_437),
.B2(n_441),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_384),
.B1(n_375),
.B2(n_364),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_402),
.B1(n_423),
.B2(n_408),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_365),
.B1(n_374),
.B2(n_372),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g489 ( 
.A(n_443),
.B(n_396),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_419),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_446),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_397),
.B1(n_383),
.B2(n_366),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_411),
.B(n_373),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_452),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_394),
.B(n_395),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_381),
.B(n_340),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_418),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_455),
.B(n_392),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_458),
.C(n_462),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_416),
.B(n_425),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_400),
.A2(n_410),
.B1(n_412),
.B2(n_406),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_413),
.B1(n_422),
.B2(n_427),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_377),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_399),
.B(n_293),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_460),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_414),
.B(n_382),
.Y(n_462)
);

AOI221xp5_ASAP7_75t_L g463 ( 
.A1(n_457),
.A2(n_420),
.B1(n_409),
.B2(n_403),
.C(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_463),
.B(n_486),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_434),
.A2(n_424),
.B1(n_401),
.B2(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_406),
.Y(n_471)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_434),
.A2(n_430),
.B1(n_415),
.B2(n_418),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_477),
.B1(n_488),
.B2(n_451),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_473),
.A2(n_481),
.B1(n_445),
.B2(n_448),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_475),
.B(n_478),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_363),
.Y(n_476)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_437),
.A2(n_392),
.B1(n_377),
.B2(n_382),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_455),
.A2(n_353),
.B(n_368),
.C(n_378),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_440),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_480),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_451),
.A2(n_459),
.B1(n_439),
.B2(n_456),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_456),
.A2(n_376),
.B(n_363),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_483),
.A2(n_484),
.B(n_435),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_SL g484 ( 
.A(n_441),
.B(n_353),
.C(n_378),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_368),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_433),
.Y(n_490)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_432),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_487),
.B(n_467),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_436),
.A2(n_392),
.B1(n_376),
.B2(n_396),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_442),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_499),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_433),
.C(n_458),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_492),
.B(n_493),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_471),
.Y(n_493)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_459),
.B1(n_453),
.B2(n_450),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_498),
.A2(n_511),
.B1(n_473),
.B2(n_469),
.Y(n_517)
);

XNOR2x1_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_454),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_449),
.C(n_462),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_505),
.C(n_507),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_504),
.A2(n_506),
.B1(n_488),
.B2(n_477),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_475),
.C(n_483),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_468),
.A2(n_445),
.B1(n_438),
.B2(n_327),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_324),
.C(n_328),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_354),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_478),
.C(n_474),
.Y(n_526)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_510),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_361),
.B1(n_347),
.B2(n_312),
.Y(n_511)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_513),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_476),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g541 ( 
.A1(n_514),
.A2(n_478),
.A3(n_491),
.B1(n_511),
.B2(n_499),
.C(n_500),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_504),
.A2(n_464),
.B1(n_472),
.B2(n_470),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_516),
.A2(n_527),
.B1(n_497),
.B2(n_502),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_517),
.A2(n_518),
.B1(n_496),
.B2(n_501),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_494),
.A2(n_480),
.B1(n_484),
.B2(n_489),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_498),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_521),
.B(n_529),
.Y(n_539)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_512),
.Y(n_524)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_508),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_509),
.A2(n_478),
.B1(n_465),
.B2(n_361),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_501),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_495),
.B(n_326),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_531),
.Y(n_546)
);

FAx1_ASAP7_75t_SL g533 ( 
.A(n_526),
.B(n_505),
.CI(n_491),
.CON(n_533),
.SN(n_533)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_523),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_520),
.B(n_490),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_538),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_530),
.A2(n_503),
.B(n_507),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_535),
.A2(n_543),
.B(n_515),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_536),
.A2(n_541),
.B1(n_514),
.B2(n_518),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_492),
.C(n_522),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_543),
.C(n_545),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_544),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_519),
.B(n_312),
.C(n_309),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_524),
.A2(n_320),
.B(n_291),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_294),
.C(n_303),
.Y(n_545)
);

AO21x1_ASAP7_75t_L g561 ( 
.A1(n_547),
.A2(n_533),
.B(n_542),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_516),
.C(n_523),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_550),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_525),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_552),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_520),
.C(n_513),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_528),
.C(n_527),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_555),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_536),
.B(n_303),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_544),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_561),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_556),
.C(n_552),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_563),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_554),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_534),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_566),
.C(n_564),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_553),
.C(n_554),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g567 ( 
.A1(n_558),
.A2(n_548),
.B(n_546),
.Y(n_567)
);

A2O1A1O1Ixp25_ASAP7_75t_L g576 ( 
.A1(n_567),
.A2(n_565),
.B(n_287),
.C(n_291),
.D(n_315),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_570),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_557),
.C(n_545),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_561),
.A2(n_533),
.B1(n_285),
.B2(n_304),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_572),
.B(n_560),
.Y(n_575)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_566),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_575),
.Y(n_578)
);

OAI321xp33_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_287),
.A3(n_572),
.B1(n_291),
.B2(n_320),
.C(n_315),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g579 ( 
.A1(n_577),
.A2(n_287),
.B(n_291),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_578),
.C(n_282),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_569),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_581),
.B(n_574),
.Y(n_582)
);

AO21x1_ASAP7_75t_L g583 ( 
.A1(n_582),
.A2(n_304),
.B(n_315),
.Y(n_583)
);

FAx1_ASAP7_75t_SL g584 ( 
.A(n_583),
.B(n_320),
.CI(n_227),
.CON(n_584),
.SN(n_584)
);


endmodule