module real_aes_170_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_454;
wire n_565;
wire n_443;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_582;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_250;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_531;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_361;
wire n_246;
wire n_412;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_536;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_589;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_349;
wire n_336;
wire n_420;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_241;
wire n_393;
wire n_294;
wire n_258;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_0), .A2(n_204), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_1), .A2(n_172), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_2), .A2(n_83), .B1(n_332), .B2(n_451), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_3), .A2(n_94), .B1(n_298), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_4), .A2(n_77), .B1(n_267), .B2(n_419), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g486 ( .A1(n_5), .A2(n_70), .B1(n_205), .B2(n_331), .C1(n_379), .C2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_6), .A2(n_49), .B1(n_324), .B2(n_325), .Y(n_323) );
OA22x2_ASAP7_75t_L g369 ( .A1(n_7), .A2(n_370), .B1(n_371), .B2(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_7), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_8), .A2(n_60), .B1(n_264), .B2(n_350), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_9), .A2(n_130), .B1(n_390), .B2(n_391), .Y(n_480) );
AO22x2_ASAP7_75t_L g232 ( .A1(n_10), .A2(n_156), .B1(n_233), .B2(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g572 ( .A(n_10), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_11), .A2(n_134), .B1(n_320), .B2(n_321), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_12), .A2(n_133), .B1(n_332), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_13), .A2(n_62), .B1(n_318), .B2(n_348), .Y(n_347) );
XOR2x2_ASAP7_75t_L g494 ( .A(n_14), .B(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_15), .A2(n_155), .B1(n_376), .B2(n_461), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_16), .A2(n_81), .B1(n_390), .B2(n_391), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_17), .A2(n_85), .B1(n_267), .B2(n_437), .Y(n_559) );
AO22x2_ASAP7_75t_L g236 ( .A1(n_18), .A2(n_48), .B1(n_233), .B2(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_18), .B(n_571), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_19), .A2(n_45), .B1(n_298), .B2(n_300), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_20), .A2(n_161), .B1(n_448), .B2(n_449), .Y(n_447) );
AOI22xp5_ASAP7_75t_SL g283 ( .A1(n_21), .A2(n_187), .B1(n_284), .B2(n_286), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_22), .A2(n_124), .B1(n_343), .B2(n_345), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_23), .A2(n_110), .B1(n_324), .B2(n_325), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_24), .B(n_356), .Y(n_355) );
OA22x2_ASAP7_75t_L g432 ( .A1(n_25), .A2(n_433), .B1(n_434), .B2(n_454), .Y(n_432) );
INVx1_ASAP7_75t_L g454 ( .A(n_25), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_26), .A2(n_34), .B1(n_386), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_27), .A2(n_184), .B1(n_273), .B2(n_318), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_28), .A2(n_576), .B1(n_589), .B2(n_590), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_28), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_29), .A2(n_120), .B1(n_264), .B2(n_499), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_30), .A2(n_152), .B1(n_271), .B2(n_537), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_31), .A2(n_145), .B1(n_252), .B2(n_260), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_32), .A2(n_196), .B1(n_298), .B2(n_511), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_33), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_35), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_36), .A2(n_66), .B1(n_252), .B2(n_315), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_37), .A2(n_167), .B1(n_413), .B2(n_415), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_38), .A2(n_139), .B1(n_314), .B2(n_315), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_39), .A2(n_141), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_40), .A2(n_127), .B1(n_327), .B2(n_328), .Y(n_326) );
OAI22x1_ASAP7_75t_SL g398 ( .A1(n_41), .A2(n_399), .B1(n_429), .B2(n_430), .Y(n_398) );
INVx1_ASAP7_75t_L g429 ( .A(n_41), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_42), .A2(n_46), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_43), .A2(n_84), .B1(n_320), .B2(n_321), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_44), .A2(n_165), .B1(n_405), .B2(n_407), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_47), .A2(n_50), .B1(n_437), .B2(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_51), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_52), .A2(n_162), .B1(n_327), .B2(n_328), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_53), .A2(n_73), .B1(n_229), .B2(n_246), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_54), .A2(n_123), .B1(n_176), .B2(n_291), .C1(n_330), .C2(n_332), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_55), .A2(n_150), .B1(n_469), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_56), .A2(n_114), .B1(n_286), .B2(n_363), .Y(n_512) );
INVx3_ASAP7_75t_L g233 ( .A(n_57), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_58), .A2(n_122), .B1(n_324), .B2(n_325), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_59), .A2(n_111), .B1(n_276), .B2(n_439), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_61), .A2(n_203), .B1(n_318), .B2(n_437), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_63), .A2(n_191), .B1(n_264), .B2(n_267), .Y(n_263) );
XNOR2x2_ASAP7_75t_L g455 ( .A(n_64), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_65), .B(n_403), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_67), .A2(n_181), .B1(n_376), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_68), .A2(n_86), .B1(n_261), .B2(n_271), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_69), .B(n_279), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_71), .A2(n_103), .B1(n_229), .B2(n_312), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_72), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_74), .A2(n_121), .B1(n_271), .B2(n_275), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_75), .A2(n_102), .B1(n_328), .B2(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_76), .A2(n_96), .B1(n_229), .B2(n_246), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_78), .A2(n_99), .B1(n_363), .B2(n_364), .Y(n_362) );
INVx1_ASAP7_75t_SL g244 ( .A(n_79), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_79), .B(n_100), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_80), .A2(n_171), .B1(n_260), .B2(n_498), .Y(n_560) );
INVx2_ASAP7_75t_L g217 ( .A(n_82), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_87), .A2(n_194), .B1(n_385), .B2(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_88), .B(n_279), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_89), .A2(n_117), .B1(n_298), .B2(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_90), .A2(n_170), .B1(n_376), .B2(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_91), .A2(n_182), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_92), .A2(n_200), .B1(n_414), .B2(n_511), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_93), .A2(n_183), .B1(n_261), .B2(n_264), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_95), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_97), .A2(n_157), .B1(n_324), .B2(n_325), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_98), .A2(n_180), .B1(n_252), .B2(n_350), .Y(n_349) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_100), .A2(n_163), .B1(n_233), .B2(n_240), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_101), .A2(n_175), .B1(n_291), .B2(n_332), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_104), .A2(n_208), .B(n_218), .C(n_574), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_105), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_106), .A2(n_195), .B1(n_332), .B2(n_514), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_107), .A2(n_154), .B1(n_320), .B2(n_321), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_108), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_109), .A2(n_142), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_112), .A2(n_179), .B1(n_298), .B2(n_446), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_113), .A2(n_197), .B1(n_229), .B2(n_312), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_115), .A2(n_148), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_116), .A2(n_199), .B1(n_409), .B2(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g245 ( .A(n_118), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_119), .A2(n_143), .B1(n_284), .B2(n_550), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_125), .A2(n_178), .B1(n_284), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_126), .A2(n_135), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_128), .A2(n_188), .B1(n_422), .B2(n_424), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_129), .A2(n_132), .B1(n_385), .B2(n_386), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_131), .A2(n_147), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_136), .A2(n_202), .B1(n_320), .B2(n_321), .Y(n_464) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_137), .B(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_138), .A2(n_166), .B1(n_252), .B2(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_140), .A2(n_164), .B1(n_229), .B2(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_144), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_146), .A2(n_151), .B1(n_284), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_149), .A2(n_201), .B1(n_529), .B2(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_153), .B(n_516), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g522 ( .A(n_158), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_159), .A2(n_189), .B1(n_248), .B2(n_343), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_160), .A2(n_206), .B1(n_509), .B2(n_511), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_168), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_169), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g568 ( .A(n_169), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_173), .A2(n_193), .B1(n_390), .B2(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
AND2x2_ASAP7_75t_R g592 ( .A(n_174), .B(n_568), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_177), .B(n_516), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_185), .A2(n_192), .B1(n_291), .B2(n_293), .Y(n_290) );
INVxp67_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_190), .B(n_332), .Y(n_358) );
AO22x1_ASAP7_75t_L g595 ( .A1(n_198), .A2(n_577), .B1(n_596), .B2(n_597), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_198), .Y(n_596) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AND2x4_ASAP7_75t_SL g210 ( .A(n_211), .B(n_214), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g603 ( .A(n_212), .B(n_214), .Y(n_603) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_213), .B(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_472), .B1(n_563), .B2(n_564), .C(n_565), .Y(n_218) );
INVx1_ASAP7_75t_L g563 ( .A(n_219), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B1(n_394), .B2(n_471), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_334), .B1(n_335), .B2(n_393), .Y(n_221) );
INVx1_ASAP7_75t_L g393 ( .A(n_222), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B1(n_306), .B2(n_307), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
XNOR2x1_ASAP7_75t_L g225 ( .A(n_226), .B(n_305), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_277), .Y(n_226) );
NAND4xp25_ASAP7_75t_L g227 ( .A(n_228), .B(n_251), .C(n_263), .D(n_270), .Y(n_227) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g344 ( .A(n_230), .Y(n_344) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_238), .Y(n_230) );
AND2x4_ASAP7_75t_L g269 ( .A(n_231), .B(n_258), .Y(n_269) );
AND2x2_ASAP7_75t_L g299 ( .A(n_231), .B(n_274), .Y(n_299) );
AND2x6_ASAP7_75t_L g321 ( .A(n_231), .B(n_258), .Y(n_321) );
AND2x4_ASAP7_75t_L g324 ( .A(n_231), .B(n_274), .Y(n_324) );
AND2x2_ASAP7_75t_L g385 ( .A(n_231), .B(n_238), .Y(n_385) );
AND2x2_ASAP7_75t_SL g482 ( .A(n_231), .B(n_238), .Y(n_482) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
AND2x2_ASAP7_75t_L g250 ( .A(n_232), .B(n_236), .Y(n_250) );
INVx2_ASAP7_75t_L g257 ( .A(n_232), .Y(n_257) );
INVx1_ASAP7_75t_L g234 ( .A(n_233), .Y(n_234) );
INVx2_ASAP7_75t_L g237 ( .A(n_233), .Y(n_237) );
INVx1_ASAP7_75t_L g240 ( .A(n_233), .Y(n_240) );
OAI22x1_ASAP7_75t_L g242 ( .A1(n_233), .A2(n_243), .B1(n_244), .B2(n_245), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_233), .Y(n_243) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_235), .Y(n_304) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g256 ( .A(n_236), .Y(n_256) );
AND2x4_ASAP7_75t_L g262 ( .A(n_236), .B(n_257), .Y(n_262) );
AND2x2_ASAP7_75t_L g266 ( .A(n_238), .B(n_255), .Y(n_266) );
AND2x4_ASAP7_75t_L g285 ( .A(n_238), .B(n_262), .Y(n_285) );
AND2x6_ASAP7_75t_L g320 ( .A(n_238), .B(n_255), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_238), .B(n_262), .Y(n_327) );
AND2x2_ASAP7_75t_L g379 ( .A(n_238), .B(n_262), .Y(n_379) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
BUFx2_ASAP7_75t_L g249 ( .A(n_239), .Y(n_249) );
INVx2_ASAP7_75t_L g259 ( .A(n_239), .Y(n_259) );
AND2x2_ASAP7_75t_L g282 ( .A(n_239), .B(n_242), .Y(n_282) );
AND2x4_ASAP7_75t_L g258 ( .A(n_241), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g274 ( .A(n_242), .B(n_259), .Y(n_274) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g345 ( .A(n_247), .Y(n_345) );
INVx2_ASAP7_75t_L g424 ( .A(n_247), .Y(n_424) );
INVx5_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
BUFx2_ASAP7_75t_L g534 ( .A(n_248), .Y(n_534) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x4_ASAP7_75t_L g386 ( .A(n_249), .B(n_250), .Y(n_386) );
AND2x4_ASAP7_75t_L g276 ( .A(n_250), .B(n_258), .Y(n_276) );
AND2x2_ASAP7_75t_L g295 ( .A(n_250), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_250), .B(n_296), .Y(n_377) );
AND2x4_ASAP7_75t_L g391 ( .A(n_250), .B(n_258), .Y(n_391) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_250), .B(n_296), .Y(n_461) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_SL g314 ( .A(n_253), .Y(n_314) );
INVx2_ASAP7_75t_L g426 ( .A(n_253), .Y(n_426) );
INVx2_ASAP7_75t_SL g437 ( .A(n_253), .Y(n_437) );
INVx4_ASAP7_75t_L g468 ( .A(n_253), .Y(n_468) );
INVx2_ASAP7_75t_SL g536 ( .A(n_253), .Y(n_536) );
INVx8_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
AND2x4_ASAP7_75t_L g273 ( .A(n_255), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_255), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g331 ( .A(n_255), .B(n_282), .Y(n_331) );
AND2x2_ASAP7_75t_L g390 ( .A(n_255), .B(n_274), .Y(n_390) );
AND2x2_ASAP7_75t_L g484 ( .A(n_255), .B(n_258), .Y(n_484) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVxp67_ASAP7_75t_L g289 ( .A(n_257), .Y(n_289) );
AND2x4_ASAP7_75t_L g261 ( .A(n_258), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g469 ( .A(n_258), .B(n_262), .Y(n_469) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_261), .Y(n_315) );
INVx2_ASAP7_75t_L g441 ( .A(n_261), .Y(n_441) );
BUFx3_ASAP7_75t_L g527 ( .A(n_261), .Y(n_527) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_261), .Y(n_588) );
AND2x2_ASAP7_75t_L g292 ( .A(n_262), .B(n_274), .Y(n_292) );
AND2x4_ASAP7_75t_L g376 ( .A(n_262), .B(n_274), .Y(n_376) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_SL g529 ( .A(n_265), .Y(n_529) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g420 ( .A(n_266), .Y(n_420) );
BUFx2_ASAP7_75t_L g498 ( .A(n_266), .Y(n_498) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g350 ( .A(n_268), .Y(n_350) );
INVx2_ASAP7_75t_L g499 ( .A(n_268), .Y(n_499) );
INVx1_ASAP7_75t_SL g530 ( .A(n_268), .Y(n_530) );
INVx8_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g501 ( .A(n_272), .Y(n_501) );
INVx2_ASAP7_75t_L g526 ( .A(n_272), .Y(n_526) );
INVx6_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g348 ( .A(n_273), .Y(n_348) );
BUFx3_ASAP7_75t_L g439 ( .A(n_273), .Y(n_439) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx3_ASAP7_75t_L g318 ( .A(n_276), .Y(n_318) );
INVx2_ASAP7_75t_L g503 ( .A(n_276), .Y(n_503) );
NAND4xp25_ASAP7_75t_SL g277 ( .A(n_278), .B(n_283), .C(n_290), .D(n_297), .Y(n_277) );
INVx4_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx3_ASAP7_75t_SL g381 ( .A(n_280), .Y(n_381) );
INVx4_ASAP7_75t_SL g403 ( .A(n_280), .Y(n_403) );
INVx3_ASAP7_75t_L g516 ( .A(n_280), .Y(n_516) );
INVx6_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g288 ( .A(n_282), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g302 ( .A(n_282), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g325 ( .A(n_282), .B(n_303), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_282), .B(n_289), .Y(n_328) );
AND2x2_ASAP7_75t_L g487 ( .A(n_282), .B(n_289), .Y(n_487) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g363 ( .A(n_285), .Y(n_363) );
BUFx2_ASAP7_75t_L g448 ( .A(n_285), .Y(n_448) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g364 ( .A(n_287), .Y(n_364) );
INVx2_ASAP7_75t_L g407 ( .A(n_287), .Y(n_407) );
INVx2_ASAP7_75t_L g449 ( .A(n_287), .Y(n_449) );
INVx2_ASAP7_75t_SL g541 ( .A(n_287), .Y(n_541) );
INVx2_ASAP7_75t_L g550 ( .A(n_287), .Y(n_550) );
INVx6_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_291), .Y(n_409) );
BUFx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g357 ( .A(n_292), .Y(n_357) );
BUFx5_ASAP7_75t_L g514 ( .A(n_292), .Y(n_514) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g411 ( .A(n_294), .Y(n_411) );
INVx2_ASAP7_75t_L g452 ( .A(n_294), .Y(n_452) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_299), .Y(n_414) );
INVx3_ASAP7_75t_L g510 ( .A(n_299), .Y(n_510) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_SL g361 ( .A(n_302), .Y(n_361) );
INVx2_ASAP7_75t_L g416 ( .A(n_302), .Y(n_416) );
BUFx3_ASAP7_75t_L g446 ( .A(n_302), .Y(n_446) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_302), .Y(n_511) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
XOR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_333), .Y(n_308) );
NAND4xp75_ASAP7_75t_L g309 ( .A(n_310), .B(n_316), .C(n_322), .D(n_329), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_318), .Y(n_427) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g354 ( .A(n_331), .Y(n_354) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_366), .B1(n_367), .B2(n_392), .Y(n_335) );
INVx1_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
XOR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_365), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_351), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g423 ( .A(n_344), .Y(n_423) );
INVx2_ASAP7_75t_L g533 ( .A(n_344), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_359), .Y(n_351) );
OAI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_355), .C(n_358), .Y(n_352) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g451 ( .A(n_357), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2x1_ASAP7_75t_L g372 ( .A(n_373), .B(n_382), .Y(n_372) );
NAND4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .C(n_378), .D(n_380), .Y(n_373) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_381), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_388), .C(n_389), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_431), .B2(n_470), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g430 ( .A(n_399), .Y(n_430) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_417), .Y(n_399) );
NAND4xp25_ASAP7_75t_SL g400 ( .A(n_401), .B(n_404), .C(n_408), .D(n_412), .Y(n_400) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g417 ( .A(n_418), .B(n_421), .C(n_425), .D(n_428), .Y(n_417) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g470 ( .A(n_431), .Y(n_470) );
XNOR2x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_455), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .C(n_442), .D(n_443), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g506 ( .A(n_441), .Y(n_506) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .C(n_450), .D(n_453), .Y(n_444) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_463), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .C(n_460), .D(n_462), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .C(n_466), .D(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g564 ( .A(n_472), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_520), .B2(n_562), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_491), .B1(n_517), .B2(n_518), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g517 ( .A(n_476), .Y(n_517) );
XNOR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_490), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .C(n_481), .D(n_483), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .C(n_489), .Y(n_485) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_494), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .C(n_504), .D(n_505), .Y(n_496) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g537 ( .A(n_503), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .C(n_513), .D(n_515), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g562 ( .A(n_520), .Y(n_562) );
AO22x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_545), .B2(n_561), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_538), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .C(n_531), .D(n_535), .Y(n_524) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .C(n_542), .D(n_543), .Y(n_538) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g561 ( .A(n_546), .Y(n_561) );
NAND4xp75_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .C(n_555), .D(n_558), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_567), .B(n_570), .Y(n_600) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI222xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_591), .B1(n_593), .B2(n_596), .C1(n_598), .C2(n_601), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_576), .Y(n_590) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g597 ( .A(n_577), .Y(n_597) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .C(n_581), .D(n_582), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .C(n_586), .D(n_587), .Y(n_583) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_599), .Y(n_598) );
CKINVDCx6p67_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_603), .Y(n_602) );
endmodule