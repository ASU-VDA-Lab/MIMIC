module real_jpeg_10294_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_304, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_304;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_244;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_40),
.B1(n_50),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_102),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_102),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_102),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_144),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_10),
.A2(n_40),
.B1(n_50),
.B2(n_144),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_11),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_153),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_13),
.A2(n_40),
.B1(n_50),
.B2(n_153),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_14),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_40),
.B1(n_50),
.B2(n_76),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_15),
.A2(n_58),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_58),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_15),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_15),
.A2(n_27),
.B1(n_33),
.B2(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_52),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_42),
.B(n_46),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_15),
.A2(n_40),
.B1(n_50),
.B2(n_162),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_20),
.B(n_110),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_21),
.B(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_21),
.B(n_295),
.Y(n_302)
);

FAx1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.CI(n_91),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_55),
.B2(n_71),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_25),
.A2(n_38),
.B(n_71),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_25),
.A2(n_26),
.B1(n_56),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_27),
.A2(n_33),
.B1(n_143),
.B2(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_27),
.A2(n_96),
.B(n_146),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_27),
.A2(n_34),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_27),
.A2(n_33),
.B1(n_209),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_27),
.A2(n_195),
.B(n_231),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_28),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_28),
.A2(n_32),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_29),
.A2(n_30),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_29),
.B(n_65),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_29),
.B(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_30),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_32),
.B(n_95),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_33),
.B(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_33),
.A2(n_94),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_48),
.B(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_39),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_39),
.A2(n_44),
.B1(n_245),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_39),
.A2(n_44),
.B1(n_101),
.B2(n_254),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_40),
.A2(n_41),
.B(n_162),
.C(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_44),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_78),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_46),
.B(n_162),
.CON(n_187),
.SN(n_187)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_52),
.A2(n_118),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_66),
.B(n_68),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_64),
.B1(n_66),
.B2(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_57),
.A2(n_64),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_57),
.A2(n_64),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_57),
.A2(n_64),
.B1(n_152),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_57),
.A2(n_64),
.B1(n_177),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_57),
.A2(n_84),
.B(n_185),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_59),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_58),
.B(n_78),
.Y(n_193)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_59),
.A2(n_80),
.B1(n_187),
.B2(n_193),
.Y(n_192)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_64),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_64),
.A2(n_87),
.B(n_98),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_69),
.A2(n_86),
.B(n_89),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_83),
.B(n_90),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_77),
.A2(n_81),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_77),
.A2(n_125),
.B(n_257),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_81),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_112),
.B1(n_113),
.B2(n_130),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_90),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_104),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_92),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_93),
.B(n_97),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_106),
.A2(n_122),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_106),
.A2(n_122),
.B1(n_205),
.B2(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_131),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B(n_124),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_122),
.A2(n_241),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI321xp33_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_282),
.A3(n_294),
.B1(n_296),
.B2(n_302),
.C(n_304),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_247),
.C(n_278),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_221),
.B(n_246),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_198),
.B(n_220),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_180),
.B(n_197),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_171),
.B(n_179),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_159),
.B(n_170),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_158),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_165),
.B(n_169),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_181),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.CI(n_178),
.CON(n_174),
.SN(n_174)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_191),
.B2(n_196),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_190),
.C(n_196),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_214),
.B2(n_215),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_217),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_213),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_208),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_223),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_234),
.C(n_235),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_239),
.C(n_242),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_265),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_248),
.B(n_265),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.C(n_263),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_252),
.C(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_258),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_274),
.C(n_275),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_270),
.C(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_297),
.B(n_301),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_291),
.C(n_293),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B(n_300),
.Y(n_297)
);


endmodule