module fake_jpeg_14206_n_527 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_527);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_17),
.B(n_1),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_67),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_51),
.B1(n_47),
.B2(n_45),
.Y(n_105)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_65),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_20),
.B(n_2),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_81),
.Y(n_110)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_42),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_100),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_5),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_28),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_101),
.Y(n_147)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_15),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_105),
.A2(n_134),
.B1(n_95),
.B2(n_62),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_35),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_148),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_146),
.B1(n_157),
.B2(n_161),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_40),
.B1(n_35),
.B2(n_45),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_40),
.B1(n_50),
.B2(n_41),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_21),
.B1(n_36),
.B2(n_44),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_51),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_80),
.A2(n_25),
.B1(n_41),
.B2(n_38),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_52),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_23),
.B(n_29),
.C(n_46),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_36),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_156),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_64),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_76),
.B(n_36),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_68),
.A2(n_50),
.B1(n_25),
.B2(n_26),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_71),
.A2(n_50),
.B1(n_26),
.B2(n_27),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_162),
.B(n_179),
.Y(n_234)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_164),
.Y(n_264)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_169),
.Y(n_242)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_114),
.A2(n_61),
.B1(n_60),
.B2(n_37),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_172),
.A2(n_180),
.B1(n_181),
.B2(n_194),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_173),
.B(n_197),
.Y(n_253)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_148),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_192),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_64),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_177),
.B(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_129),
.A2(n_37),
.B1(n_26),
.B2(n_27),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_120),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_182),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_47),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_121),
.B(n_44),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_128),
.B(n_23),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_103),
.B(n_21),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_195),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_113),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_96),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_143),
.B(n_30),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_113),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_207),
.B1(n_109),
.B2(n_158),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_55),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_218),
.C(n_146),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_201),
.A2(n_208),
.B1(n_46),
.B2(n_29),
.Y(n_256)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_206),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_94),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_204),
.B(n_209),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_5),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_93),
.B1(n_90),
.B2(n_87),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_126),
.A2(n_86),
.B1(n_56),
.B2(n_75),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_124),
.Y(n_210)
);

BUFx8_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_214),
.Y(n_266)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_216),
.Y(n_246)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_219),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_115),
.B(n_83),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_232),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_131),
.B1(n_161),
.B2(n_157),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_223),
.A2(n_168),
.B1(n_218),
.B2(n_210),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_227),
.B1(n_238),
.B2(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_133),
.B1(n_106),
.B2(n_140),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_183),
.B(n_128),
.CI(n_109),
.CON(n_229),
.SN(n_229)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_229),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_73),
.B1(n_74),
.B2(n_140),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_241),
.B1(n_256),
.B2(n_268),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_163),
.A2(n_155),
.B(n_122),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_235),
.A2(n_185),
.B(n_202),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_125),
.B1(n_160),
.B2(n_158),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_125),
.B1(n_160),
.B2(n_124),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_29),
.B1(n_46),
.B2(n_7),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_46),
.C(n_29),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_252),
.C(n_219),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_46),
.Y(n_252)
);

AO22x1_ASAP7_75t_SL g259 ( 
.A1(n_196),
.A2(n_46),
.B1(n_29),
.B2(n_8),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_193),
.B(n_10),
.C(n_11),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_166),
.B(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_175),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_188),
.A2(n_29),
.B1(n_8),
.B2(n_9),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_171),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_167),
.B1(n_184),
.B2(n_174),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_221),
.A2(n_169),
.B(n_204),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_271),
.A2(n_250),
.B(n_236),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_170),
.B(n_165),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_272),
.A2(n_276),
.B(n_306),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_182),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_281),
.B(n_284),
.Y(n_323)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_245),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_297),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_226),
.A2(n_213),
.B1(n_198),
.B2(n_192),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_220),
.A2(n_203),
.B1(n_209),
.B2(n_217),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_288),
.A2(n_308),
.B1(n_260),
.B2(n_243),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_301),
.B1(n_302),
.B2(n_312),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_186),
.A3(n_206),
.B1(n_178),
.B2(n_211),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_218),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_294),
.C(n_313),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_193),
.Y(n_294)
);

OA22x2_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_310),
.B1(n_260),
.B2(n_233),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_230),
.B(n_189),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_296),
.B(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_228),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_229),
.B(n_214),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_305),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_225),
.A2(n_227),
.B1(n_229),
.B2(n_259),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_251),
.A2(n_164),
.B1(n_216),
.B2(n_212),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_304),
.Y(n_342)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_307),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_232),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_259),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_12),
.Y(n_311)
);

NAND2x1_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_244),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_235),
.A2(n_13),
.B1(n_14),
.B2(n_231),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_13),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_236),
.A2(n_13),
.B1(n_14),
.B2(n_268),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_314),
.A2(n_315),
.B1(n_284),
.B2(n_305),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_236),
.A2(n_14),
.B1(n_241),
.B2(n_255),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_242),
.B(n_234),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_331),
.B(n_343),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_275),
.A2(n_269),
.B1(n_257),
.B2(n_246),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_321),
.A2(n_327),
.B1(n_328),
.B2(n_349),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_315),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_275),
.A2(n_258),
.B1(n_266),
.B2(n_262),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_276),
.A2(n_258),
.B1(n_228),
.B2(n_264),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_271),
.B(n_306),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_311),
.B(n_295),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_285),
.A2(n_273),
.B(n_299),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_341),
.C(n_356),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_282),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_347),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_301),
.A2(n_264),
.B1(n_249),
.B2(n_233),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_334),
.A2(n_339),
.B1(n_280),
.B2(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_355),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_293),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_243),
.B(n_222),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_287),
.A2(n_222),
.B(n_224),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_346),
.A2(n_351),
.B(n_355),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_311),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_274),
.A2(n_244),
.B(n_224),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_298),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_333),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_272),
.A2(n_254),
.B(n_244),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_290),
.B(n_254),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_323),
.B(n_313),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_368),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_SL g419 ( 
.A(n_361),
.B(n_326),
.Y(n_419)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_272),
.A3(n_312),
.B1(n_314),
.B2(n_295),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_322),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_366),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_379),
.B1(n_328),
.B2(n_324),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_369),
.Y(n_403)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_375),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_319),
.B(n_350),
.Y(n_399)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_332),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_382),
.C(n_384),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_325),
.A2(n_295),
.B1(n_310),
.B2(n_303),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_14),
.B1(n_310),
.B2(n_334),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_390),
.B1(n_339),
.B2(n_323),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_310),
.C(n_317),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_381),
.B1(n_373),
.B2(n_374),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_329),
.C(n_343),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_338),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_386),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_316),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_350),
.C(n_318),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_326),
.C(n_345),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_389),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_342),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_316),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_393),
.A2(n_377),
.B1(n_357),
.B2(n_358),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_327),
.B1(n_356),
.B2(n_335),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_398),
.A2(n_404),
.B1(n_417),
.B2(n_372),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_364),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_321),
.B1(n_349),
.B2(n_319),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_346),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_407),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_320),
.Y(n_407)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_381),
.A2(n_373),
.B1(n_391),
.B2(n_382),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_409),
.A2(n_412),
.B1(n_340),
.B2(n_365),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_351),
.B1(n_347),
.B2(n_340),
.Y(n_410)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_410),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_320),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_415),
.C(n_421),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_368),
.A2(n_340),
.B1(n_353),
.B2(n_345),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_385),
.A2(n_340),
.B1(n_342),
.B2(n_330),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_419),
.B(n_361),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_342),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_390),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_386),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_441),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_384),
.Y(n_427)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_362),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_439),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_417),
.A2(n_362),
.B(n_391),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_395),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_431),
.A2(n_435),
.B1(n_404),
.B2(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_421),
.C(n_411),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_446),
.C(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_369),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_413),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_442),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_359),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_444),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_363),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_445),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_371),
.C(n_375),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_392),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_403),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_448),
.A2(n_397),
.B1(n_400),
.B2(n_405),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_463),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_409),
.C(n_399),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_461),
.C(n_465),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_424),
.C(n_443),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_464),
.B(n_430),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_418),
.C(n_393),
.Y(n_465)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_467),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_436),
.A2(n_418),
.B(n_403),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_468),
.A2(n_445),
.B(n_447),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_472),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_453),
.B(n_436),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_482),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_464),
.B(n_428),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_476),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_440),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_438),
.C(n_440),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_480),
.C(n_458),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_459),
.A2(n_468),
.B(n_429),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_481),
.B(n_449),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_466),
.A2(n_431),
.B1(n_435),
.B2(n_423),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_479),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_438),
.C(n_432),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_454),
.A2(n_397),
.B1(n_400),
.B2(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_460),
.Y(n_483)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_483),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_451),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_465),
.C(n_454),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_492),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_487),
.Y(n_501)
);

BUFx24_ASAP7_75t_SL g488 ( 
.A(n_473),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_493),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_498),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g492 ( 
.A(n_477),
.B(n_450),
.CI(n_459),
.CON(n_492),
.SN(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_456),
.C(n_462),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_456),
.C(n_448),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_497),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_496),
.A2(n_478),
.B(n_475),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_452),
.C(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_479),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_506),
.Y(n_516)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_505),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_495),
.A2(n_472),
.B(n_470),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_508),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_482),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_491),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_491),
.B1(n_486),
.B2(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_514),
.A2(n_515),
.B(n_499),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_500),
.B(n_449),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_510),
.A2(n_503),
.B(n_509),
.Y(n_517)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_520),
.C(n_516),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_502),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_522),
.A2(n_516),
.B(n_518),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_515),
.C(n_521),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_524),
.A2(n_511),
.B(n_504),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_420),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_420),
.B1(n_376),
.B2(n_330),
.Y(n_527)
);


endmodule