module real_aes_4400_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_0), .A2(n_570), .B(n_572), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_1), .Y(n_505) );
INVx1_ASAP7_75t_L g244 ( .A(n_2), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_3), .A2(n_15), .B1(n_84), .B2(n_197), .Y(n_220) );
INVx2_ASAP7_75t_L g177 ( .A(n_4), .Y(n_177) );
INVx1_ASAP7_75t_SL g117 ( .A(n_5), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_6), .A2(n_20), .B1(n_511), .B2(n_533), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_7), .B(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_8), .A2(n_51), .B1(n_542), .B2(n_548), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_9), .B(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_10), .A2(n_23), .B1(n_551), .B2(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g530 ( .A(n_11), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_11), .B(n_57), .Y(n_580) );
INVxp67_ASAP7_75t_L g592 ( .A(n_11), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_12), .A2(n_43), .B1(n_249), .B2(n_250), .Y(n_248) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_13), .A2(n_55), .B(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_13), .A2(n_55), .B(n_111), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_14), .B(n_515), .Y(n_526) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_15), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_16), .A2(n_65), .B1(n_585), .B2(n_586), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_17), .B(n_155), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_18), .A2(n_62), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx2_ASAP7_75t_L g201 ( .A(n_19), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_21), .A2(n_26), .B1(n_115), .B2(n_152), .Y(n_221) );
BUFx3_ASAP7_75t_L g610 ( .A(n_22), .Y(n_610) );
O2A1O1Ixp5_ASAP7_75t_L g194 ( .A1(n_24), .A2(n_88), .B(n_195), .C(n_196), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_25), .A2(n_52), .B1(n_174), .B2(n_175), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_27), .Y(n_153) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_28), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_29), .A2(n_64), .B1(n_257), .B2(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g190 ( .A(n_30), .Y(n_190) );
INVx1_ASAP7_75t_L g516 ( .A(n_31), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_31), .B(n_56), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_32), .B(n_186), .Y(n_239) );
INVx2_ASAP7_75t_L g198 ( .A(n_33), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_34), .B(n_562), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_35), .Y(n_156) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_36), .Y(n_598) );
INVx2_ASAP7_75t_L g207 ( .A(n_37), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_38), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g124 ( .A(n_39), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_40), .Y(n_597) );
INVx1_ASAP7_75t_L g148 ( .A(n_41), .Y(n_148) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_44), .A2(n_45), .B1(n_558), .B2(n_559), .Y(n_557) );
AND2x4_ASAP7_75t_L g91 ( .A(n_46), .B(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_L g142 ( .A(n_46), .B(n_92), .Y(n_142) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_46), .Y(n_620) );
INVx1_ASAP7_75t_L g573 ( .A(n_47), .Y(n_573) );
INVx1_ASAP7_75t_L g132 ( .A(n_48), .Y(n_132) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_50), .A2(n_506), .B1(n_507), .B2(n_623), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_50), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_53), .B(n_119), .Y(n_211) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_53), .Y(n_634) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_54), .A2(n_57), .B1(n_515), .B2(n_519), .Y(n_520) );
INVx1_ASAP7_75t_L g538 ( .A(n_54), .Y(n_538) );
INVx1_ASAP7_75t_L g532 ( .A(n_56), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_56), .B(n_536), .Y(n_583) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_56), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_57), .A2(n_63), .B(n_540), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_58), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_59), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_60), .B(n_116), .Y(n_127) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_61), .Y(n_602) );
INVx1_ASAP7_75t_L g518 ( .A(n_63), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_63), .B(n_74), .Y(n_581) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
BUFx5_ASAP7_75t_L g126 ( .A(n_66), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_67), .B(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g210 ( .A(n_68), .Y(n_210) );
INVx1_ASAP7_75t_L g214 ( .A(n_69), .Y(n_214) );
INVx2_ASAP7_75t_L g160 ( .A(n_70), .Y(n_160) );
INVx2_ASAP7_75t_SL g92 ( .A(n_71), .Y(n_92) );
AOI22xp5_ASAP7_75t_SL g565 ( .A1(n_72), .A2(n_75), .B1(n_566), .B2(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_73), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_74), .B(n_525), .Y(n_524) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_76), .A2(n_90), .A3(n_199), .B1(n_219), .B2(n_223), .Y(n_218) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_76), .A2(n_219), .B1(n_313), .B2(n_315), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_500), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_90), .Y(n_79) );
OA21x2_ASAP7_75t_L g629 ( .A1(n_80), .A2(n_630), .B(n_631), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx2_ASAP7_75t_L g192 ( .A(n_84), .Y(n_192) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_84), .Y(n_259) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g116 ( .A(n_85), .Y(n_116) );
INVx2_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
INVx6_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_87), .B(n_141), .Y(n_150) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_88), .A2(n_220), .B1(n_221), .B2(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_88), .A2(n_234), .B(n_236), .Y(n_233) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx3_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
INVx4_ASAP7_75t_L g187 ( .A(n_89), .Y(n_187) );
INVx1_ASAP7_75t_L g261 ( .A(n_89), .Y(n_261) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx3_ASAP7_75t_L g112 ( .A(n_91), .Y(n_112) );
AND2x2_ASAP7_75t_L g166 ( .A(n_91), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g313 ( .A(n_91), .B(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_92), .Y(n_618) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
BUFx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_SL g97 ( .A(n_98), .Y(n_97) );
NAND2x1p5_ASAP7_75t_L g98 ( .A(n_99), .B(n_385), .Y(n_98) );
AND3x1_ASAP7_75t_L g99 ( .A(n_100), .B(n_341), .C(n_369), .Y(n_99) );
NOR3xp33_ASAP7_75t_SL g100 ( .A(n_101), .B(n_278), .C(n_317), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_262), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_162), .B(n_215), .C(n_227), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g305 ( .A(n_104), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g319 ( .A(n_104), .B(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_104), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g461 ( .A(n_104), .Y(n_461) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_133), .Y(n_104) );
INVxp67_ASAP7_75t_SL g272 ( .A(n_105), .Y(n_272) );
OR2x2_ASAP7_75t_L g345 ( .A(n_105), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g267 ( .A(n_106), .Y(n_267) );
AND2x2_ASAP7_75t_L g280 ( .A(n_106), .B(n_274), .Y(n_280) );
OR2x2_ASAP7_75t_L g288 ( .A(n_106), .B(n_133), .Y(n_288) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_106), .Y(n_292) );
INVx1_ASAP7_75t_L g332 ( .A(n_106), .Y(n_332) );
INVx1_ASAP7_75t_L g402 ( .A(n_106), .Y(n_402) );
AO31x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_113), .A3(n_123), .B(n_129), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx2_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g158 ( .A(n_110), .Y(n_158) );
INVx2_ASAP7_75t_L g178 ( .A(n_110), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_112), .B(n_131), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_112), .B(n_131), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_112), .B(n_131), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_117), .B(n_118), .C(n_122), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g171 ( .A(n_116), .Y(n_171) );
INVx1_ASAP7_75t_L g235 ( .A(n_116), .Y(n_235) );
INVx1_ASAP7_75t_L g250 ( .A(n_116), .Y(n_250) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g174 ( .A(n_120), .Y(n_174) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g139 ( .A(n_121), .Y(n_139) );
INVx1_ASAP7_75t_L g172 ( .A(n_122), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_122), .A2(n_138), .B(n_210), .C(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g222 ( .A(n_122), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_122), .B(n_252), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B(n_127), .C(n_128), .Y(n_123) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g152 ( .A(n_126), .Y(n_152) );
INVx2_ASAP7_75t_L g237 ( .A(n_126), .Y(n_237) );
INVx1_ASAP7_75t_L g241 ( .A(n_126), .Y(n_241) );
INVx2_ASAP7_75t_L g249 ( .A(n_126), .Y(n_249) );
INVx3_ASAP7_75t_L g143 ( .A(n_128), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_128), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_132), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_130), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
BUFx3_ASAP7_75t_L g254 ( .A(n_131), .Y(n_254) );
INVx1_ASAP7_75t_L g314 ( .A(n_131), .Y(n_314) );
INVx2_ASAP7_75t_L g265 ( .A(n_133), .Y(n_265) );
BUFx2_ASAP7_75t_L g447 ( .A(n_133), .Y(n_447) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_157), .B(n_159), .Y(n_133) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_134), .A2(n_159), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_149), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B1(n_144), .B2(n_147), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
NOR3xp33_ASAP7_75t_L g147 ( .A(n_141), .B(n_143), .C(n_148), .Y(n_147) );
AOI221x1_ASAP7_75t_L g181 ( .A1(n_141), .A2(n_182), .B1(n_185), .B2(n_189), .C(n_191), .Y(n_181) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_143), .A2(n_169), .B1(n_172), .B2(n_173), .Y(n_168) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g258 ( .A(n_146), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
OAI22xp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B1(n_154), .B2(n_156), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_154), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx2_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
INVx2_ASAP7_75t_SL g197 ( .A(n_155), .Y(n_197) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_179), .Y(n_162) );
INVx2_ASAP7_75t_L g310 ( .A(n_163), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_163), .B(n_179), .Y(n_326) );
INVx4_ASAP7_75t_L g354 ( .A(n_163), .Y(n_354) );
AND2x2_ASAP7_75t_L g494 ( .A(n_163), .B(n_339), .Y(n_494) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g300 ( .A(n_164), .Y(n_300) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
INVx1_ASAP7_75t_L g360 ( .A(n_165), .Y(n_360) );
AOI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_176), .Y(n_165) );
INVx3_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx1_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
BUFx3_ASAP7_75t_L g199 ( .A(n_178), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_178), .B(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
AND2x2_ASAP7_75t_L g276 ( .A(n_179), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g294 ( .A(n_179), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g297 ( .A(n_179), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g441 ( .A(n_179), .B(n_346), .Y(n_441) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_202), .Y(n_179) );
INVx2_ASAP7_75t_L g225 ( .A(n_180), .Y(n_225) );
INVx1_ASAP7_75t_L g340 ( .A(n_180), .Y(n_340) );
AND2x2_ASAP7_75t_L g373 ( .A(n_180), .B(n_203), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_180), .B(n_360), .Y(n_421) );
OR2x2_ASAP7_75t_L g469 ( .A(n_180), .B(n_360), .Y(n_469) );
AO31x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_193), .A3(n_199), .B(n_200), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
AND2x2_ASAP7_75t_L g189 ( .A(n_186), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_187), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx2_ASAP7_75t_L g315 ( .A(n_199), .Y(n_315) );
AND2x4_ASAP7_75t_L g350 ( .A(n_202), .B(n_312), .Y(n_350) );
AND2x2_ASAP7_75t_L g395 ( .A(n_202), .B(n_226), .Y(n_395) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x4_ASAP7_75t_L g216 ( .A(n_203), .B(n_217), .Y(n_216) );
BUFx3_ASAP7_75t_L g316 ( .A(n_203), .Y(n_316) );
AND2x4_ASAP7_75t_L g339 ( .A(n_203), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g366 ( .A(n_203), .Y(n_366) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_209), .A3(n_212), .B(n_213), .Y(n_204) );
AO22x1_ASAP7_75t_L g635 ( .A1(n_207), .A2(n_506), .B1(n_507), .B2(n_636), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_207), .Y(n_636) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_224), .Y(n_215) );
INVx2_ASAP7_75t_L g384 ( .A(n_216), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_216), .A2(n_404), .B(n_407), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_217), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g355 ( .A(n_217), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx8_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
AND2x2_ASAP7_75t_L g474 ( .A(n_218), .B(n_300), .Y(n_474) );
INVxp67_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_224), .B(n_350), .Y(n_436) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_SL g356 ( .A(n_225), .Y(n_356) );
BUFx3_ASAP7_75t_L g394 ( .A(n_225), .Y(n_394) );
INVx1_ASAP7_75t_L g473 ( .A(n_225), .Y(n_473) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_226), .Y(n_320) );
INVx2_ASAP7_75t_L g346 ( .A(n_226), .Y(n_346) );
INVx1_ASAP7_75t_L g357 ( .A(n_227), .Y(n_357) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g291 ( .A(n_228), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g471 ( .A(n_228), .B(n_280), .Y(n_471) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_246), .Y(n_228) );
INVx2_ASAP7_75t_L g269 ( .A(n_229), .Y(n_269) );
INVx1_ASAP7_75t_L g284 ( .A(n_229), .Y(n_284) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_229), .Y(n_290) );
INVx1_ASAP7_75t_L g308 ( .A(n_229), .Y(n_308) );
AND2x2_ASAP7_75t_L g465 ( .A(n_229), .B(n_267), .Y(n_465) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_238), .B(n_245), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .Y(n_238) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g303 ( .A(n_246), .Y(n_303) );
INVx1_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
INVx1_ASAP7_75t_L g379 ( .A(n_246), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_247), .B(n_255), .Y(n_246) );
AND2x2_ASAP7_75t_SL g283 ( .A(n_247), .B(n_255), .Y(n_283) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_251), .B(n_253), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_252), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_260), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_270), .B(n_276), .Y(n_262) );
INVx2_ASAP7_75t_L g368 ( .A(n_263), .Y(n_368) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
AND2x2_ASAP7_75t_L g301 ( .A(n_264), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g399 ( .A(n_264), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_264), .B(n_382), .Y(n_427) );
AND2x4_ASAP7_75t_L g435 ( .A(n_264), .B(n_307), .Y(n_435) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g492 ( .A(n_265), .B(n_303), .Y(n_492) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g425 ( .A(n_268), .B(n_280), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_268), .B(n_447), .Y(n_455) );
AND2x2_ASAP7_75t_L g476 ( .A(n_268), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g273 ( .A(n_269), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g410 ( .A(n_271), .Y(n_410) );
OR2x6_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_273), .Y(n_336) );
INVxp67_ASAP7_75t_L g380 ( .A(n_273), .Y(n_380) );
AND2x2_ASAP7_75t_L g329 ( .A(n_274), .B(n_303), .Y(n_329) );
AND2x2_ASAP7_75t_L g349 ( .A(n_274), .B(n_308), .Y(n_349) );
AND2x2_ASAP7_75t_L g486 ( .A(n_274), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
INVx1_ASAP7_75t_L g325 ( .A(n_277), .Y(n_325) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_277), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g372 ( .A(n_277), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_277), .B(n_420), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_277), .B(n_348), .C(n_349), .D(n_394), .Y(n_430) );
BUFx3_ASAP7_75t_L g440 ( .A(n_277), .Y(n_440) );
OR2x2_ASAP7_75t_L g449 ( .A(n_277), .B(n_450), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_293), .B(n_296), .C(n_304), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_285), .B2(n_289), .C(n_291), .Y(n_279) );
OAI322xp33_ASAP7_75t_L g351 ( .A1(n_280), .A2(n_352), .A3(n_357), .B1(n_358), .B2(n_361), .C1(n_362), .C2(n_368), .Y(n_351) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_L g400 ( .A(n_283), .B(n_284), .Y(n_400) );
INVx1_ASAP7_75t_L g452 ( .A(n_283), .Y(n_452) );
INVx2_ASAP7_75t_L g487 ( .A(n_283), .Y(n_487) );
INVx1_ASAP7_75t_L g383 ( .A(n_284), .Y(n_383) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g438 ( .A(n_287), .B(n_400), .Y(n_438) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g416 ( .A(n_288), .B(n_378), .Y(n_416) );
AND2x4_ASAP7_75t_L g491 ( .A(n_289), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g330 ( .A(n_290), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g406 ( .A(n_299), .Y(n_406) );
OR2x2_ASAP7_75t_L g413 ( .A(n_299), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_302), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g460 ( .A(n_302), .Y(n_460) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g488 ( .A(n_308), .B(n_402), .Y(n_488) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g397 ( .A(n_311), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_311), .B(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
AND2x2_ASAP7_75t_L g359 ( .A(n_312), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
INVx1_ASAP7_75t_L g391 ( .A(n_312), .Y(n_391) );
INVx2_ASAP7_75t_SL g490 ( .A(n_316), .Y(n_490) );
OAI322xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .A3(n_324), .B1(n_326), .B2(n_327), .C1(n_333), .C2(n_337), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_319), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g348 ( .A(n_323), .B(n_331), .Y(n_348) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_329), .A2(n_370), .B(n_374), .Y(n_369) );
INVxp67_ASAP7_75t_L g477 ( .A(n_331), .Y(n_477) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_334), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_339), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g450 ( .A(n_339), .Y(n_450) );
O2A1O1Ixp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_347), .B(n_350), .C(n_351), .Y(n_341) );
INVxp33_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI32xp33_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_375), .A3(n_376), .B1(n_381), .B2(n_384), .Y(n_374) );
INVx1_ASAP7_75t_L g364 ( .A(n_346), .Y(n_364) );
BUFx3_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
AND2x2_ASAP7_75t_L g489 ( .A(n_346), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_346), .B(n_356), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_347), .A2(n_388), .B(n_396), .Y(n_387) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVxp67_ASAP7_75t_R g361 ( .A(n_348), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_350), .B(n_354), .Y(n_443) );
AND2x4_ASAP7_75t_L g467 ( .A(n_350), .B(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g478 ( .A(n_350), .B(n_394), .Y(n_478) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g484 ( .A(n_356), .Y(n_484) );
AOI21xp33_ASAP7_75t_SL g442 ( .A1(n_358), .A2(n_443), .B(n_444), .Y(n_442) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_360), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_397), .B1(n_398), .B2(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_372), .Y(n_375) );
INVxp67_ASAP7_75t_L g422 ( .A(n_372), .Y(n_422) );
AND2x2_ASAP7_75t_L g390 ( .A(n_373), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
INVx2_ASAP7_75t_L g454 ( .A(n_373), .Y(n_454) );
INVx1_ASAP7_75t_L g462 ( .A(n_375), .Y(n_462) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_377), .A2(n_438), .B1(n_439), .B2(n_441), .Y(n_437) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g445 ( .A(n_382), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR3x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_431), .C(n_479), .Y(n_385) );
NAND3xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_403), .C(n_411), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g429 ( .A(n_391), .B(n_420), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_406), .B(n_454), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_407), .A2(n_494), .B(n_495), .Y(n_493) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B1(n_417), .B2(n_423), .C(n_426), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_424), .A2(n_481), .B(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_429), .A2(n_471), .B1(n_476), .B2(n_478), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_456), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_442), .C(n_448), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g498 ( .A(n_438), .B(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B1(n_453), .B2(n_455), .Y(n_448) );
INVx1_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_462), .B(n_463), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NOR2x1p5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B(n_470), .C(n_475), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_473), .B(n_474), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .C(n_497), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_489), .B2(n_491), .Y(n_483) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_604), .B1(n_621), .B2(n_624), .C(n_626), .Y(n_500) );
XOR2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_593), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_506), .B2(n_507), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVxp33_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_560), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_510), .B(n_541), .C(n_550), .D(n_557), .Y(n_509) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
AND2x4_ASAP7_75t_L g558 ( .A(n_512), .B(n_546), .Y(n_558) );
AND2x2_ASAP7_75t_L g564 ( .A(n_512), .B(n_555), .Y(n_564) );
AND2x4_ASAP7_75t_L g585 ( .A(n_512), .B(n_552), .Y(n_585) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
INVx1_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
NAND2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g519 ( .A(n_515), .Y(n_519) );
INVx3_ASAP7_75t_L g525 ( .A(n_515), .Y(n_525) );
NAND2xp33_ASAP7_75t_L g531 ( .A(n_515), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g540 ( .A(n_515), .Y(n_540) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_515), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_516), .B(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_L g614 ( .A(n_516), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_518), .A2(n_540), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g545 ( .A(n_520), .Y(n_545) );
AND2x2_ASAP7_75t_L g567 ( .A(n_520), .B(n_544), .Y(n_567) );
AND2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g533 ( .A(n_521), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g549 ( .A(n_522), .Y(n_549) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
AND2x4_ASAP7_75t_L g546 ( .A(n_523), .B(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g552 ( .A(n_523), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g556 ( .A(n_523), .Y(n_556) );
AND2x2_ASAP7_75t_L g587 ( .A(n_523), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_525), .B(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_L g536 ( .A(n_525), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_526), .B(n_535), .C(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g547 ( .A(n_527), .Y(n_547) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g553 ( .A(n_528), .Y(n_553) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
AND2x4_ASAP7_75t_L g559 ( .A(n_534), .B(n_546), .Y(n_559) );
AND2x4_ASAP7_75t_L g568 ( .A(n_534), .B(n_555), .Y(n_568) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_538), .Y(n_615) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
AND2x4_ASAP7_75t_L g548 ( .A(n_543), .B(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g551 ( .A(n_543), .B(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g554 ( .A(n_543), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x4_ASAP7_75t_L g566 ( .A(n_552), .B(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g555 ( .A(n_553), .B(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g571 ( .A(n_555), .B(n_567), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .C(n_569), .D(n_584), .Y(n_560) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_579), .B(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_578), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x4_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_589), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_599), .B1(n_600), .B2(n_603), .Y(n_593) );
INVx1_ASAP7_75t_L g603 ( .A(n_594), .Y(n_603) );
XOR2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
XOR2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
BUFx10_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_616), .Y(n_607) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g639 ( .A(n_609), .B(n_616), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_612), .C(n_615), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
OR2x2_ASAP7_75t_L g625 ( .A(n_617), .B(n_620), .Y(n_625) );
INVx1_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_617), .B(n_619), .Y(n_631) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_632), .B1(n_635), .B2(n_637), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
CKINVDCx14_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
endmodule