module fake_netlist_1_11433_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_7), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
BUFx6f_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
OR2x6_ASAP7_75t_L g16 ( .A(n_9), .B(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_17), .B(n_8), .Y(n_19) );
OAI21xp5_ASAP7_75t_L g20 ( .A1(n_14), .A2(n_13), .B(n_11), .Y(n_20) );
OR2x2_ASAP7_75t_SL g21 ( .A(n_16), .B(n_10), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_15), .A2(n_10), .B(n_3), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_20), .B(n_16), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_19), .B(n_16), .Y(n_24) );
A2O1A1Ixp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_22), .B(n_18), .C(n_19), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_24), .B(n_18), .C(n_10), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_21), .B1(n_15), .B2(n_14), .C(n_5), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_27), .Y(n_29) );
BUFx2_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
OAI22xp5_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_21), .B1(n_3), .B2(n_4), .Y(n_31) );
OAI31xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_2), .A3(n_6), .B(n_22), .Y(n_32) );
AOI22xp5_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_2), .B1(n_30), .B2(n_32), .Y(n_33) );
endmodule