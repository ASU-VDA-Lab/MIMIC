module fake_jpeg_15873_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_5),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_52),
.B1(n_50),
.B2(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_74),
.B1(n_60),
.B2(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_73),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_57),
.B1(n_61),
.B2(n_47),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_78),
.B(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_61),
.B1(n_47),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_0),
.Y(n_94)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_82),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_49),
.B1(n_55),
.B2(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_58),
.C(n_56),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_51),
.C(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_58),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_98),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_104)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_8),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_114),
.B1(n_100),
.B2(n_9),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_102),
.B1(n_86),
.B2(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_107),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_9),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_105),
.C(n_26),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_111),
.C(n_112),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_115),
.B(n_119),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_105),
.B1(n_110),
.B2(n_11),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_110),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_24),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_134),
.B1(n_127),
.B2(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_133),
.C(n_20),
.Y(n_137)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_19),
.B(n_40),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_136),
.B1(n_138),
.B2(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_18),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_17),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_28),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_97),
.C(n_16),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_15),
.B1(n_36),
.B2(n_35),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_13),
.B(n_29),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_12),
.Y(n_148)
);


endmodule