module real_jpeg_3968_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_0),
.A2(n_163),
.B1(n_167),
.B2(n_170),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_0),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_183),
.C(n_187),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_0),
.B(n_79),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_0),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_0),
.B(n_131),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_0),
.B(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_1),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_1),
.Y(n_297)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_1),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_2),
.A2(n_68),
.B1(n_215),
.B2(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_2),
.A2(n_68),
.B1(n_87),
.B2(n_223),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_2),
.A2(n_68),
.B1(n_382),
.B2(n_459),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_3),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_104),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_104),
.B1(n_141),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_3),
.A2(n_104),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_4),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_4),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_4),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_4),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g445 ( 
.A(n_4),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_5),
.A2(n_57),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_5),
.A2(n_57),
.B1(n_223),
.B2(n_407),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_5),
.A2(n_57),
.B1(n_299),
.B2(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_194),
.B1(n_199),
.B2(n_200),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_8),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_163),
.B1(n_199),
.B2(n_268),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_8),
.A2(n_199),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_8),
.A2(n_199),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_11),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_11),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_174),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_11),
.A2(n_174),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_11),
.A2(n_174),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_15),
.A2(n_92),
.B1(n_94),
.B2(n_98),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_15),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_98),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_15),
.A2(n_98),
.B1(n_245),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_15),
.A2(n_98),
.B1(n_386),
.B2(n_427),
.Y(n_426)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_17),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_17),
.A2(n_225),
.B1(n_244),
.B2(n_247),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_17),
.A2(n_225),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_17),
.A2(n_225),
.B1(n_444),
.B2(n_446),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_18),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_18),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_18),
.A2(n_111),
.B1(n_291),
.B2(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_18),
.A2(n_291),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g471 ( 
.A1(n_18),
.A2(n_291),
.B1(n_366),
.B2(n_472),
.Y(n_471)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_547),
.B(n_550),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_152),
.B(n_546),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_145),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_29),
.B(n_145),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_136),
.C(n_142),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_30),
.A2(n_31),
.B1(n_542),
.B2(n_543),
.Y(n_541)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_69),
.C(n_105),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_32),
.B(n_534),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_33),
.A2(n_58),
.B1(n_60),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_33),
.A2(n_58),
.B1(n_137),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_33),
.A2(n_370),
.B(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_33),
.A2(n_46),
.B1(n_419),
.B2(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_33),
.A2(n_56),
.B1(n_58),
.B2(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_34),
.A2(n_365),
.B(n_369),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_34),
.B(n_371),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_34),
.A2(n_59),
.B(n_549),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_45),
.Y(n_347)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_46),
.B(n_170),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_47),
.Y(n_345)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g282 ( 
.A(n_49),
.Y(n_282)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_50),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_51),
.Y(n_319)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_52),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_52),
.Y(n_350)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_52),
.Y(n_380)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_52),
.Y(n_383)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_53),
.Y(n_281)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_58),
.A2(n_443),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_59),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_59),
.B(n_471),
.Y(n_470)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_63),
.Y(n_447)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_69),
.A2(n_105),
.B1(n_106),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_69),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_91),
.B1(n_99),
.B2(n_100),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_70),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_70),
.A2(n_99),
.B1(n_317),
.B2(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_70),
.A2(n_99),
.B1(n_413),
.B2(n_416),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_70),
.A2(n_91),
.B1(n_99),
.B2(n_523),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_75),
.Y(n_414)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_76),
.Y(n_306)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g448 ( 
.A1(n_79),
.A2(n_143),
.B1(n_321),
.B2(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_79),
.A2(n_143),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_85),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_86),
.Y(n_409)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_92),
.Y(n_274)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_99),
.B(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_99),
.A2(n_317),
.B(n_320),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_101),
.Y(n_415)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_105),
.A2(n_106),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_105),
.B(n_518),
.C(n_521),
.Y(n_529)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_130),
.B(n_132),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_162),
.B(n_171),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_107),
.A2(n_130),
.B1(n_222),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_107),
.A2(n_171),
.B(n_267),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_107),
.A2(n_130),
.B1(n_385),
.B2(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_108),
.B(n_172),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_108),
.A2(n_131),
.B1(n_406),
.B2(n_410),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_108),
.A2(n_131),
.B1(n_410),
.B2(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_108),
.A2(n_131),
.B1(n_426),
.B2(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_112),
.Y(n_227)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_119),
.A2(n_222),
.B(n_228),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_124),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_127),
.Y(n_246)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_127),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_127),
.Y(n_402)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_130),
.A2(n_228),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_131),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_132),
.Y(n_462)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_136),
.B(n_142),
.Y(n_543)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_143),
.A2(n_273),
.B(n_279),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_143),
.B(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_143),
.A2(n_279),
.B(n_486),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_145),
.B(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_145),
.B(n_548),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_146),
.Y(n_549)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_149),
.B(n_170),
.Y(n_351)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_540),
.B(n_545),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_512),
.B(n_537),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_390),
.A3(n_488),
.B1(n_506),
.C1(n_507),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_335),
.B(n_389),
.Y(n_155)
);

AO21x1_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_308),
.B(n_334),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_261),
.B(n_307),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_231),
.B(n_260),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_191),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_160),
.B(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_177),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_161),
.A2(n_177),
.B1(n_178),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

INVx5_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_169),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_170),
.A2(n_203),
.B(n_211),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_SL g273 ( 
.A1(n_170),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_SL g365 ( 
.A1(n_170),
.A2(n_351),
.B(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_190),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_219),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_192),
.B(n_220),
.C(n_230),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_211),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_198),
.Y(n_399)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_202),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_203),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_203),
.A2(n_396),
.B1(n_400),
.B2(n_401),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_203),
.A2(n_401),
.B(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_214),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_204),
.A2(n_212),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_204),
.A2(n_286),
.B1(n_325),
.B2(n_331),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_204),
.A2(n_357),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_207),
.Y(n_332)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_207),
.Y(n_440)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_229),
.B2(n_230),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_226),
.B(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_253),
.B(n_259),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_241),
.B(n_252),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_237),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_239),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_251),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_249),
.B(n_250),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_285),
.B(n_295),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_257),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_263),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_283),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_271),
.B2(n_272),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_271),
.C(n_283),
.Y(n_309)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI32xp33_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_299),
.A3(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_298),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_298),
.Y(n_314)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_309),
.B(n_310),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_315),
.B2(n_333),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_314),
.C(n_333),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_322),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_323),
.C(n_324),
.Y(n_359)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_342),
.A3(n_344),
.B1(n_346),
.B2(n_351),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_336),
.B(n_337),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_362),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_338)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_352),
.B2(n_353),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_341),
.B(n_352),
.Y(n_484)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx6_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_359),
.B(n_360),
.C(n_362),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_376),
.B2(n_388),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_363),
.B(n_377),
.C(n_384),
.Y(n_497)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_368),
.Y(n_472)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx8_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_376),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx6_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_474),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g507 ( 
.A1(n_391),
.A2(n_474),
.B(n_508),
.C(n_511),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_450),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_392),
.B(n_450),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_423),
.C(n_433),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_393),
.B(n_423),
.CI(n_433),
.CON(n_487),
.SN(n_487)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_411),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_412),
.C(n_418),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_405),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_405),
.Y(n_480)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

INVx4_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_418),
.Y(n_411)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_429),
.B2(n_432),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_425),
.B(n_429),
.Y(n_466)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_429),
.A2(n_432),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_429),
.A2(n_466),
.B(n_469),
.Y(n_515)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_441),
.C(n_448),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_437),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_435),
.B(n_437),
.Y(n_496)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_441),
.A2(n_442),
.B1(n_448),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_454),
.C(n_464),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_464),
.B2(n_465),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_460),
.B(n_463),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_461),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_458),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_463),
.B(n_515),
.CI(n_516),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_463),
.B(n_515),
.C(n_516),
.Y(n_536)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_475),
.B(n_487),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.C(n_481),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_485),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_482),
.A2(n_483),
.B1(n_485),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_487),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_490),
.A2(n_509),
.B(n_510),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_498),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.C(n_497),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_496),
.B1(n_497),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_503),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_526),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_525),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_525),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g554 ( 
.A(n_514),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_518),
.B1(n_520),
.B2(n_524),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_518),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_528),
.C(n_532),
.Y(n_544)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_526),
.A2(n_538),
.B(n_539),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_536),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_536),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_544),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_544),
.Y(n_545)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);


endmodule