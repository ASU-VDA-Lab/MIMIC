module fake_jpeg_16704_n_293 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_14),
.B(n_19),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_41),
.B(n_19),
.C(n_16),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_14),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_25),
.B(n_17),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_27),
.B1(n_16),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_19),
.B1(n_16),
.B2(n_25),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_27),
.B1(n_47),
.B2(n_39),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_101)
);

OAI22x1_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_20),
.B1(n_21),
.B2(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_68),
.B1(n_17),
.B2(n_22),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_35),
.B1(n_22),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_23),
.B1(n_18),
.B2(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_74),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_28),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_75),
.C(n_76),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_17),
.B(n_21),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_20),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_17),
.B(n_21),
.C(n_28),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_87),
.Y(n_111)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_81),
.Y(n_124)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_62),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_20),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_92),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22x1_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_62),
.B1(n_75),
.B2(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_20),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_55),
.B1(n_68),
.B2(n_62),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_123),
.B1(n_98),
.B2(n_67),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_68),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_101),
.B(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_83),
.B(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_62),
.B1(n_64),
.B2(n_61),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_60),
.C(n_75),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_127),
.A2(n_131),
.B(n_135),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_128),
.B(n_130),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_114),
.B1(n_113),
.B2(n_83),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_140),
.B1(n_146),
.B2(n_95),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_87),
.B(n_86),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_90),
.C(n_99),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_145),
.C(n_127),
.Y(n_154)
);

NAND2x1p5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_86),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_141),
.B(n_109),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_117),
.B1(n_121),
.B2(n_125),
.Y(n_140)
);

NAND2x1_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_86),
.Y(n_141)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_57),
.B(n_81),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_144),
.B1(n_106),
.B2(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_79),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_84),
.B1(n_78),
.B2(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_103),
.B(n_79),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_103),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_162),
.C(n_163),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_181),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_110),
.B1(n_107),
.B2(n_116),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_160),
.B1(n_166),
.B2(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_111),
.C(n_119),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_111),
.C(n_119),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_109),
.B1(n_92),
.B2(n_91),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_169),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_91),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_135),
.C(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_89),
.B1(n_77),
.B2(n_42),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_44),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_21),
.B(n_44),
.C(n_30),
.D(n_3),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_180),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_44),
.B(n_30),
.C(n_2),
.D(n_3),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_140),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_193),
.C(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_143),
.B1(n_153),
.B2(n_144),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_205),
.B(n_179),
.C(n_166),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_162),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_146),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_143),
.B1(n_128),
.B2(n_40),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_40),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_40),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_51),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_51),
.C(n_42),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_193),
.C(n_196),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_189),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_171),
.Y(n_210)
);

XOR2x1_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_216),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_163),
.Y(n_220)
);

NAND2x1_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_176),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_223),
.C(n_202),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_175),
.C(n_157),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_178),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_164),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_219),
.C(n_225),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_204),
.C(n_203),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_185),
.C(n_191),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_200),
.C(n_188),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_210),
.C(n_211),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_182),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_200),
.C(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_164),
.C(n_50),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_0),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_0),
.Y(n_241)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_249),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_254),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_230),
.A2(n_211),
.B1(n_216),
.B2(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_216),
.B(n_215),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_229),
.B(n_227),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_4),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_1),
.B(n_3),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_259),
.B(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_264),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_233),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_232),
.B1(n_239),
.B2(n_6),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_251),
.B(n_252),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_4),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_250),
.B1(n_245),
.B2(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_4),
.C(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_6),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_268),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_274),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_260),
.A2(n_244),
.B(n_242),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_273),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_7),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_265),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_6),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_275),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_257),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_257),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_269),
.B(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_11),
.C(n_12),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_270),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_281),
.C(n_12),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_9),
.B(n_10),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_290),
.A2(n_13),
.B1(n_283),
.B2(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_13),
.B(n_268),
.Y(n_293)
);


endmodule