module fake_ariane_1756_n_464 (n_83, n_8, n_56, n_60, n_64, n_119, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_464);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_464;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_124;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_130;
wire n_391;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_301;
wire n_248;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_355;
wire n_212;
wire n_123;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_407;
wire n_254;
wire n_460;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_19),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_31),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_84),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_25),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_41),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_42),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_39),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_60),
.B(n_51),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_27),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_24),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_79),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_61),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_10),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_57),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_40),
.B(n_17),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_96),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_38),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_29),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_45),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_74),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_98),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_88),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_49),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_48),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_0),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_65),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_78),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_128),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_2),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_3),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_140),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_4),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_R g207 ( 
.A(n_142),
.B(n_178),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_5),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_124),
.B(n_5),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_138),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_189),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_149),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

AND3x4_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_160),
.C(n_174),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_150),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_211),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_151),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_154),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_175),
.Y(n_241)
);

BUFx4f_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_185),
.B1(n_188),
.B2(n_193),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_134),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_207),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_132),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_195),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_158),
.Y(n_253)
);

BUFx4f_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_153),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_161),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_157),
.Y(n_260)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_202),
.A2(n_166),
.B1(n_168),
.B2(n_191),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_202),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_219),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_210),
.B1(n_229),
.B2(n_223),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_210),
.B1(n_220),
.B2(n_225),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_232),
.B(n_162),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_205),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_261),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_167),
.B1(n_177),
.B2(n_156),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_222),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_199),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_155),
.B(n_147),
.C(n_182),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_235),
.B(n_159),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_235),
.A2(n_199),
.B1(n_169),
.B2(n_186),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_170),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_260),
.B(n_181),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_203),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_184),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_192),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_257),
.B(n_172),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_251),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_244),
.B1(n_251),
.B2(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

AO22x1_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_266),
.B1(n_173),
.B2(n_179),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_288),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_227),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_276),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_281),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

BUFx8_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_292),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_267),
.A2(n_254),
.B(n_180),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_240),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_240),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_194),
.Y(n_334)
);

BUFx2_ASAP7_75t_SL g335 ( 
.A(n_275),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_302),
.A2(n_190),
.B(n_242),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_300),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_242),
.B(n_239),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_274),
.A2(n_297),
.B1(n_269),
.B2(n_279),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_274),
.B(n_230),
.Y(n_341)
);

OR2x6_ASAP7_75t_SL g342 ( 
.A(n_273),
.B(n_7),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_239),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_273),
.A2(n_246),
.B(n_245),
.C(n_243),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_337),
.A2(n_278),
.B(n_301),
.C(n_304),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

AO31x2_ASAP7_75t_L g349 ( 
.A1(n_339),
.A2(n_301),
.A3(n_278),
.B(n_298),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_275),
.Y(n_350)
);

AND2x4_ASAP7_75t_SL g351 ( 
.A(n_332),
.B(n_270),
.Y(n_351)
);

AO21x2_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_237),
.B(n_164),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_135),
.B(n_164),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_344),
.A2(n_135),
.B(n_164),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_248),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_328),
.A2(n_135),
.B(n_164),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_345),
.A2(n_164),
.B(n_135),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

AO31x2_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_323),
.A3(n_346),
.B(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

NAND2x1p5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_230),
.Y(n_364)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_324),
.B(n_311),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_321),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_62),
.B(n_9),
.Y(n_368)
);

OAI221xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

AO21x2_ASAP7_75t_L g371 ( 
.A1(n_309),
.A2(n_18),
.B(n_20),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_30),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_355),
.A2(n_329),
.B(n_331),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g376 ( 
.A1(n_353),
.A2(n_326),
.B(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_360),
.B1(n_373),
.B2(n_354),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_347),
.A2(n_331),
.B(n_320),
.C(n_315),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_327),
.B1(n_319),
.B2(n_318),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_325),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_358),
.A2(n_318),
.B(n_325),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_373),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_365),
.A2(n_35),
.B(n_36),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_37),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_352),
.A2(n_43),
.B(n_44),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_366),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_53),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_54),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_348),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_357),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

AOI221xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_369),
.B1(n_371),
.B2(n_357),
.C(n_350),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_387),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_359),
.B(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_389),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_385),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_370),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_362),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

BUFx2_ASAP7_75t_SL g409 ( 
.A(n_398),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_379),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_402),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_362),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_400),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_382),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_371),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_361),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_370),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_361),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_397),
.A2(n_383),
.B(n_386),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_349),
.Y(n_423)
);

NOR2x1_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_364),
.Y(n_424)
);

OAI31xp33_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_405),
.A3(n_407),
.B(n_403),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_396),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_396),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_423),
.B(n_399),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_406),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_406),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_56),
.Y(n_433)
);

AND3x1_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_63),
.C(n_64),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_411),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_66),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_436),
.B(n_420),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_435),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_421),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_421),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_417),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_439),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_440),
.A2(n_434),
.B(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_448),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_449),
.A2(n_450),
.B1(n_443),
.B2(n_433),
.Y(n_452)
);

AOI211xp5_ASAP7_75t_SL g453 ( 
.A1(n_451),
.A2(n_431),
.B(n_441),
.C(n_442),
.Y(n_453)
);

OAI21xp33_ASAP7_75t_SL g454 ( 
.A1(n_452),
.A2(n_428),
.B(n_422),
.Y(n_454)
);

OAI311xp33_ASAP7_75t_L g455 ( 
.A1(n_453),
.A2(n_444),
.A3(n_431),
.B1(n_433),
.C1(n_430),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_454),
.A2(n_437),
.B1(n_70),
.B2(n_72),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_455),
.B(n_67),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_457),
.B(n_76),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_458),
.B(n_456),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_77),
.B(n_80),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_461)
);

OAI222xp33_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_94),
.B1(n_97),
.B2(n_101),
.C1(n_102),
.C2(n_103),
.Y(n_462)
);

OAI221xp5_ASAP7_75t_R g463 ( 
.A1(n_462),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.C(n_110),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_464)
);


endmodule