module fake_netlist_6_971_n_1890 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1890);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1890;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_10),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_30),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_132),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_17),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_59),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_62),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_48),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_1),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_34),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_86),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_45),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_97),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_52),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_91),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_172),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_16),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_25),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_47),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_55),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_147),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_36),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_95),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_32),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_63),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_175),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_67),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_93),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_82),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_21),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_30),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_120),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_21),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_180),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_174),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_46),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_148),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_154),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_2),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_40),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_129),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_28),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_11),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_92),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_179),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_69),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_5),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_22),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_173),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_66),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_4),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_3),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_159),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_75),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_78),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_10),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_49),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_128),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_182),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_106),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_117),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_134),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_89),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_28),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_42),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_29),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_74),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_142),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_22),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_50),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_146),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_72),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_112),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_46),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_166),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_158),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_38),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_133),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_121),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_139),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_31),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_23),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_42),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_83),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_113),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_164),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_18),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_163),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_16),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_126),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_96),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_11),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_171),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_73),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_169),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_58),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_37),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_31),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_181),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_48),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_54),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_35),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_17),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_140),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_39),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_85),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_131),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_53),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_39),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_14),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_55),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_122),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_12),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_77),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_87),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_127),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_33),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_165),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_4),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_155),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_64),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_118),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_18),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_226),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_217),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_228),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_230),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_236),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_0),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_198),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_231),
.B(n_6),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_237),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_231),
.B(n_6),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_240),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_243),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_290),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_272),
.B(n_7),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_187),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_235),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_247),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_290),
.B(n_7),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_239),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_330),
.B(n_8),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_213),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_248),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_251),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_257),
.Y(n_398)
);

BUFx6f_ASAP7_75t_SL g399 ( 
.A(n_212),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_229),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_195),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_302),
.B(n_9),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_195),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_260),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_261),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_256),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_260),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_206),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_264),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_268),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_277),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_324),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_277),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_269),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_302),
.B(n_12),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_279),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_252),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_295),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_189),
.B(n_15),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_186),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_229),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_229),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_229),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_296),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_300),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_229),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_367),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_317),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_309),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_317),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_263),
.B(n_19),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_218),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_266),
.B(n_282),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_317),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_317),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_219),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_222),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_323),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_220),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_220),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_254),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_323),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_189),
.B(n_250),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_323),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_305),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_323),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_306),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_223),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_323),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_273),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_284),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_307),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_224),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_308),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_192),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_227),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_273),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_312),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_199),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_202),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_400),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_443),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_284),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_434),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_408),
.B(n_206),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_399),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_R g476 ( 
.A(n_431),
.B(n_232),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_439),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_440),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_451),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_456),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_370),
.B(n_215),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_459),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_422),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_399),
.B(n_272),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_371),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_371),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_408),
.B(n_206),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_376),
.B(n_301),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_385),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_372),
.B(n_242),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_372),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_388),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_R g511 ( 
.A(n_373),
.B(n_244),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_389),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_392),
.A2(n_278),
.B(n_250),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_401),
.B(n_359),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_444),
.B(n_359),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_463),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_446),
.B(n_301),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_373),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_403),
.B(n_364),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_462),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_374),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_460),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_411),
.B(n_246),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_393),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_413),
.B(n_364),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_406),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_412),
.A2(n_335),
.B1(n_259),
.B2(n_289),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_379),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_378),
.B(n_246),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_381),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_386),
.B(n_278),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_510),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_387),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_484),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_518),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_374),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_468),
.B(n_387),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_541),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_505),
.B(n_188),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_537),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_510),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_541),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_505),
.B(n_191),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_504),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_504),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_512),
.Y(n_563)
);

INVxp33_ASAP7_75t_SL g564 ( 
.A(n_476),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_529),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_377),
.C(n_394),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_533),
.B(n_472),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_507),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_533),
.B(n_380),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_501),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_380),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_513),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_418),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_513),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_501),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_477),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_383),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_517),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_518),
.B(n_383),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_521),
.B(n_390),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_481),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_505),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_390),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_518),
.B(n_396),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_527),
.B(n_396),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_506),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_397),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_484),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_541),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_506),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_521),
.B(n_397),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_485),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_485),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_521),
.B(n_283),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_510),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_471),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_484),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_538),
.B(n_398),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_519),
.B(n_541),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_398),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_508),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_491),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_527),
.B(n_405),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_405),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_510),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_540),
.B(n_409),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_516),
.A2(n_433),
.B1(n_466),
.B2(n_533),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_501),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_527),
.B(n_409),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_478),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_488),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_464),
.B(n_410),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_515),
.B(n_410),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_524),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_528),
.B(n_205),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_516),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_497),
.B(n_414),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_464),
.B(n_414),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_487),
.A2(n_221),
.B1(n_429),
.B2(n_211),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_283),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_524),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_532),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_467),
.B(n_473),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_474),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_532),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_467),
.B(n_417),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_509),
.B(n_417),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_420),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_515),
.B(n_420),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_514),
.A2(n_342),
.B1(n_349),
.B2(n_234),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_491),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_480),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_487),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_533),
.B(n_426),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_482),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_491),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_479),
.B(n_426),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_479),
.B(n_486),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_500),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_486),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_539),
.B(n_342),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_534),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_533),
.B(n_427),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_525),
.B(n_206),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_531),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_531),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_523),
.Y(n_663)
);

CKINVDCx6p67_ASAP7_75t_R g664 ( 
.A(n_526),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_493),
.A2(n_461),
.B1(n_457),
.B2(n_455),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_472),
.B(n_427),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_491),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_491),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_523),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_489),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_489),
.B(n_448),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_483),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_522),
.B(n_349),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_495),
.B(n_448),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_475),
.B(n_450),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_530),
.B(n_450),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_514),
.A2(n_294),
.B1(n_298),
.B2(n_356),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_528),
.B(n_206),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_500),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_495),
.B(n_455),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_496),
.B(n_457),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_523),
.B(n_461),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_490),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_499),
.B(n_453),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_475),
.B(n_212),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_499),
.B(n_216),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_502),
.B(n_207),
.Y(n_689)
);

INVx6_ASAP7_75t_L g690 ( 
.A(n_523),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_511),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_610),
.B(n_514),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_609),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_660),
.B(n_207),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_550),
.B(n_514),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_627),
.B(n_526),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_627),
.B(n_273),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_553),
.B(n_503),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_645),
.B(n_615),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_543),
.A2(n_255),
.B1(n_253),
.B2(n_265),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_655),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_660),
.B(n_553),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_574),
.B(n_502),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_552),
.A2(n_288),
.B(n_285),
.C(n_276),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_558),
.A2(n_310),
.B1(n_270),
.B2(n_271),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_545),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_563),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_682),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_558),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_596),
.B(n_503),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_556),
.A2(n_267),
.B(n_241),
.C(n_311),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_596),
.B(n_503),
.Y(n_714)
);

OAI221xp5_ASAP7_75t_L g715 ( 
.A1(n_566),
.A2(n_225),
.B1(n_314),
.B2(n_326),
.C(n_343),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_556),
.B(n_503),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_551),
.A2(n_334),
.B1(n_293),
.B2(n_297),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_571),
.B(n_207),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_581),
.B(n_214),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_679),
.A2(n_249),
.B1(n_258),
.B2(n_262),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_590),
.B(n_233),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_SL g722 ( 
.A(n_585),
.B(n_207),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_574),
.A2(n_347),
.B(n_281),
.C(n_341),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_594),
.B(n_275),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_587),
.B(n_333),
.C(n_338),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_617),
.B(n_185),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_546),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_546),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_620),
.A2(n_470),
.B(n_316),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_548),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_560),
.B(n_304),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_583),
.B(n_207),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_642),
.A2(n_202),
.B1(n_366),
.B2(n_345),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_564),
.B(n_535),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_682),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_624),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_548),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_641),
.B(n_320),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_560),
.B(n_313),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_641),
.B(n_327),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_561),
.B(n_319),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_561),
.A2(n_202),
.B1(n_340),
.B2(n_321),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_623),
.B(n_185),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_583),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_575),
.B(n_592),
.Y(n_746)
);

AND2x6_ASAP7_75t_SL g747 ( 
.A(n_628),
.B(n_535),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_683),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_575),
.B(n_470),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_592),
.B(n_274),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_586),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_563),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_586),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_686),
.B(n_329),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_611),
.B(n_614),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_611),
.B(n_287),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_292),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_629),
.B(n_190),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_568),
.B(n_299),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_637),
.Y(n_760)
);

INVxp33_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_577),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_683),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_656),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_632),
.A2(n_187),
.B1(n_197),
.B2(n_201),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_659),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_572),
.B(n_303),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_573),
.B(n_315),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_639),
.B(n_318),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_555),
.A2(n_202),
.B1(n_211),
.B2(n_209),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_649),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_684),
.B(n_322),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_555),
.B(n_202),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_678),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_638),
.B(n_346),
.C(n_369),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_555),
.B(n_328),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_577),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_559),
.B(n_202),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_559),
.A2(n_202),
.B1(n_209),
.B2(n_197),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_584),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_612),
.B(n_331),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_612),
.B(n_212),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_559),
.B(n_332),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_625),
.B(n_190),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_626),
.A2(n_202),
.B1(n_201),
.B2(n_354),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_618),
.B(n_351),
.C(n_348),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_582),
.B(n_344),
.C(n_193),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_625),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_653),
.B(n_336),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_653),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_584),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_600),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_657),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_SL g794 ( 
.A(n_687),
.B(n_691),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_633),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_671),
.B(n_337),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_667),
.B(n_204),
.C(n_208),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_633),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_635),
.A2(n_350),
.B(n_339),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_680),
.B(n_474),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_632),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_691),
.B(n_204),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_634),
.B(n_498),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_589),
.B(n_193),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_626),
.A2(n_354),
.B1(n_355),
.B2(n_208),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_598),
.A2(n_353),
.B1(n_196),
.B2(n_368),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_661),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_353),
.B1(n_196),
.B2(n_368),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_593),
.B(n_498),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_600),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_632),
.B(n_355),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_570),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_597),
.B(n_474),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_585),
.B(n_194),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_602),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_632),
.B(n_238),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_662),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_602),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_607),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_570),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_585),
.B(n_194),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_650),
.B(n_498),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_665),
.B(n_200),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_672),
.B(n_200),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_676),
.B(n_605),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_651),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_578),
.B(n_474),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_238),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_578),
.B(n_498),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_688),
.Y(n_830)
);

BUFx6f_ASAP7_75t_SL g831 ( 
.A(n_647),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_603),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_680),
.B(n_498),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_580),
.B(n_498),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_605),
.B(n_203),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_688),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_603),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_605),
.B(n_203),
.Y(n_838)
);

NAND2x1_ASAP7_75t_L g839 ( 
.A(n_601),
.B(n_498),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_605),
.A2(n_210),
.B1(n_352),
.B2(n_362),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_570),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_604),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_604),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_210),
.B1(n_352),
.B2(n_362),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_622),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_622),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_652),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_652),
.Y(n_848)
);

AOI22x1_ASAP7_75t_L g849 ( 
.A1(n_663),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_654),
.A2(n_365),
.B1(n_363),
.B2(n_357),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_585),
.B(n_361),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_654),
.B(n_365),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_565),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_681),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_681),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_761),
.B(n_599),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_795),
.B(n_636),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_692),
.A2(n_616),
.B(n_542),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_755),
.A2(n_658),
.B(n_569),
.C(n_646),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_825),
.A2(n_567),
.B(n_677),
.C(n_666),
.Y(n_860)
);

O2A1O1Ixp5_ASAP7_75t_L g861 ( 
.A1(n_695),
.A2(n_608),
.B(n_544),
.C(n_547),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_826),
.B(n_654),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_761),
.B(n_599),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_710),
.B(n_564),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_746),
.B(n_675),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_711),
.A2(n_716),
.B(n_712),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_825),
.A2(n_675),
.B1(n_670),
.B2(n_673),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_699),
.A2(n_562),
.B(n_542),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_745),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_793),
.B(n_599),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_693),
.A2(n_675),
.B1(n_674),
.B2(n_685),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_745),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_745),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_754),
.B(n_647),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_704),
.A2(n_673),
.B1(n_670),
.B2(n_680),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_736),
.B(n_607),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_700),
.B(n_621),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_714),
.A2(n_606),
.B(n_562),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_748),
.B(n_621),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_745),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_822),
.A2(n_562),
.B(n_557),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_771),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_SL g883 ( 
.A(n_819),
.B(n_644),
.Y(n_883)
);

CKINVDCx10_ASAP7_75t_R g884 ( 
.A(n_831),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_774),
.B(n_644),
.C(n_360),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_698),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_694),
.B(n_565),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_795),
.B(n_544),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_718),
.A2(n_601),
.B(n_557),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_744),
.B(n_544),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_L g891 ( 
.A(n_744),
.B(n_631),
.C(n_357),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_763),
.Y(n_892)
);

INVx3_ASAP7_75t_SL g893 ( 
.A(n_709),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_728),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_836),
.B(n_547),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_695),
.A2(n_595),
.B(n_608),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_790),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_704),
.A2(n_601),
.B1(n_690),
.B2(n_664),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_830),
.B(n_547),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_705),
.B(n_549),
.Y(n_900)
);

CKINVDCx11_ASAP7_75t_R g901 ( 
.A(n_747),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_739),
.B(n_647),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_728),
.Y(n_903)
);

AND2x6_ASAP7_75t_SL g904 ( 
.A(n_782),
.B(n_664),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

CKINVDCx8_ASAP7_75t_R g906 ( 
.A(n_752),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_719),
.B(n_549),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_729),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_837),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_750),
.A2(n_601),
.B1(n_690),
.B2(n_595),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_721),
.A2(n_724),
.B(n_772),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_718),
.A2(n_690),
.B(n_608),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_758),
.A2(n_549),
.B(n_554),
.C(n_669),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_741),
.B(n_363),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_803),
.A2(n_636),
.B(n_630),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_756),
.B(n_554),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_788),
.B(n_636),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_812),
.A2(n_630),
.B(n_643),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_812),
.A2(n_630),
.B(n_643),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_757),
.B(n_554),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_802),
.B(n_238),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_751),
.B(n_595),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_706),
.A2(n_648),
.B(n_669),
.C(n_668),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_812),
.A2(n_643),
.B(n_570),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_788),
.B(n_570),
.Y(n_925)
);

O2A1O1Ixp5_ASAP7_75t_L g926 ( 
.A1(n_733),
.A2(n_804),
.B(n_773),
.C(n_778),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_697),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_842),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_758),
.B(n_613),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_777),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_737),
.B(n_613),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_788),
.B(n_619),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_SL g933 ( 
.A1(n_733),
.A2(n_648),
.B(n_669),
.C(n_668),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_791),
.Y(n_934)
);

BUFx12f_ASAP7_75t_SL g935 ( 
.A(n_782),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_706),
.A2(n_613),
.B(n_648),
.C(n_668),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_846),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_734),
.A2(n_690),
.B1(n_643),
.B2(n_591),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_820),
.A2(n_619),
.B(n_591),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_820),
.A2(n_619),
.B(n_591),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_734),
.A2(n_680),
.B(n_689),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_824),
.B(n_576),
.C(n_588),
.Y(n_942)
);

INVx11_ASAP7_75t_L g943 ( 
.A(n_831),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_827),
.A2(n_576),
.B(n_619),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_791),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_824),
.A2(n_576),
.B(n_588),
.C(n_591),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_737),
.B(n_576),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_832),
.B(n_619),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_820),
.A2(n_841),
.B(n_778),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_727),
.A2(n_753),
.B1(n_804),
.B2(n_835),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_703),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_727),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_832),
.B(n_591),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_781),
.B(n_588),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_715),
.A2(n_245),
.B(n_280),
.C(n_291),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_841),
.A2(n_588),
.B(n_689),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_835),
.A2(n_588),
.B(n_280),
.C(n_291),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_854),
.B(n_689),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_841),
.A2(n_689),
.B(n_100),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_787),
.B(n_94),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_773),
.A2(n_689),
.B(n_102),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_788),
.B(n_291),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_784),
.B(n_245),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_854),
.B(n_689),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_806),
.B(n_280),
.Y(n_965)
);

CKINVDCx10_ASAP7_75t_R g966 ( 
.A(n_782),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_829),
.A2(n_245),
.B(n_84),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_809),
.A2(n_81),
.B(n_168),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_760),
.B(n_76),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_751),
.A2(n_71),
.B1(n_167),
.B2(n_160),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_784),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_813),
.A2(n_70),
.B(n_153),
.Y(n_972)
);

OA22x2_ASAP7_75t_L g973 ( 
.A1(n_801),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_789),
.A2(n_88),
.B(n_149),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_852),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_838),
.A2(n_65),
.B1(n_145),
.B2(n_141),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_764),
.B(n_115),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_766),
.B(n_176),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_838),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_979)
);

AO21x1_ASAP7_75t_L g980 ( 
.A1(n_720),
.A2(n_27),
.B(n_32),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_735),
.B(n_34),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_785),
.B(n_104),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_785),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_SL g984 ( 
.A1(n_732),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_770),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_848),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_805),
.B(n_56),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_796),
.A2(n_111),
.B(n_105),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_723),
.A2(n_57),
.B(n_107),
.C(n_108),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_702),
.B(n_57),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_798),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_853),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_770),
.B(n_779),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_731),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_801),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_776),
.A2(n_109),
.B(n_116),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_779),
.B(n_119),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_798),
.B(n_855),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_798),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_738),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_783),
.A2(n_123),
.B(n_125),
.Y(n_1001)
);

AO32x2_ASAP7_75t_L g1002 ( 
.A1(n_713),
.A2(n_723),
.A3(n_765),
.B1(n_805),
.B2(n_850),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_L g1003 ( 
.A(n_794),
.B(n_775),
.C(n_725),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_850),
.B(n_811),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_834),
.A2(n_767),
.B(n_759),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_768),
.A2(n_749),
.B(n_847),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_844),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_762),
.B(n_815),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_780),
.B(n_818),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_792),
.B(n_845),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_843),
.B(n_810),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_769),
.B(n_765),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_701),
.A2(n_708),
.B(n_833),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_839),
.Y(n_1014)
);

AO22x1_ASAP7_75t_L g1015 ( 
.A1(n_797),
.A2(n_786),
.B1(n_807),
.B2(n_817),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_823),
.B(n_828),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_808),
.B(n_840),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_717),
.B(n_707),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_800),
.A2(n_851),
.B(n_821),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_816),
.B(n_828),
.Y(n_1020)
);

AO21x1_ASAP7_75t_L g1021 ( 
.A1(n_740),
.A2(n_742),
.B(n_730),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_814),
.A2(n_851),
.B(n_821),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_814),
.A2(n_810),
.B(n_799),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_849),
.B(n_713),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_743),
.B(n_816),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_743),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_816),
.B(n_828),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_722),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_696),
.A2(n_550),
.B(n_553),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_793),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_737),
.A2(n_552),
.B(n_543),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_755),
.A2(n_704),
.B(n_706),
.C(n_695),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_692),
.A2(n_718),
.B(n_822),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_825),
.A2(n_755),
.B1(n_826),
.B2(n_704),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_696),
.A2(n_550),
.B(n_553),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1034),
.B(n_865),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_993),
.A2(n_1017),
.B1(n_982),
.B2(n_997),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_SL g1038 ( 
.A1(n_946),
.A2(n_859),
.B(n_1032),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_865),
.B(n_993),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_982),
.A2(n_997),
.B1(n_1026),
.B2(n_990),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_1012),
.A2(n_1018),
.B1(n_987),
.B2(n_965),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_952),
.B(n_1031),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_952),
.B(n_950),
.Y(n_1043)
);

AOI221x1_ASAP7_75t_L g1044 ( 
.A1(n_957),
.A2(n_860),
.B1(n_1003),
.B2(n_942),
.C(n_913),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_926),
.A2(n_1035),
.B(n_861),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_889),
.A2(n_858),
.B(n_1033),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_868),
.A2(n_878),
.B(n_949),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_897),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_1021),
.A2(n_980),
.A3(n_929),
.B(n_920),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_916),
.A2(n_920),
.B(n_866),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_900),
.B(n_862),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1030),
.B(n_870),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1019),
.A2(n_1005),
.B(n_1006),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_L g1055 ( 
.A1(n_1024),
.A2(n_1015),
.B(n_1023),
.C(n_1022),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_884),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_SL g1057 ( 
.A1(n_862),
.A2(n_1025),
.B(n_929),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_899),
.Y(n_1058)
);

BUFx4f_ASAP7_75t_SL g1059 ( 
.A(n_992),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_890),
.A2(n_910),
.A3(n_979),
.B(n_983),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_954),
.A2(n_1025),
.B(n_1004),
.C(n_977),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_877),
.B(n_887),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_931),
.B(n_914),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_969),
.A2(n_978),
.B(n_977),
.C(n_925),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_905),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_907),
.A2(n_953),
.B(n_948),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_888),
.A2(n_938),
.B(n_998),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_947),
.B(n_886),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_883),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_895),
.B(n_921),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_895),
.B(n_874),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_902),
.B(n_909),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_899),
.B(n_928),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_894),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_906),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_937),
.B(n_986),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_969),
.A2(n_978),
.B(n_975),
.C(n_955),
.Y(n_1077)
);

AOI211x1_ASAP7_75t_L g1078 ( 
.A1(n_891),
.A2(n_996),
.B(n_1001),
.C(n_896),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_951),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_985),
.A2(n_867),
.B(n_981),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_918),
.A2(n_919),
.B(n_924),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1013),
.A2(n_936),
.B(n_923),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_948),
.A2(n_953),
.B(n_998),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_873),
.B(n_880),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_903),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1007),
.A2(n_871),
.B1(n_885),
.B2(n_927),
.C(n_995),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_856),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_893),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_873),
.B(n_880),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_939),
.A2(n_940),
.B(n_915),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_908),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_971),
.A2(n_963),
.B(n_989),
.C(n_960),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_941),
.A2(n_964),
.B(n_958),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_863),
.B(n_922),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_892),
.B(n_864),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1016),
.A2(n_976),
.B(n_1000),
.C(n_994),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_876),
.B(n_879),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_SL g1098 ( 
.A1(n_974),
.A2(n_988),
.B(n_972),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_991),
.B(n_1014),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_922),
.B(n_934),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_999),
.Y(n_1101)
);

AND2x2_ASAP7_75t_SL g1102 ( 
.A(n_1020),
.B(n_1027),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1020),
.B(n_1002),
.Y(n_1103)
);

AO21x1_ASAP7_75t_L g1104 ( 
.A1(n_970),
.A2(n_968),
.B(n_898),
.Y(n_1104)
);

CKINVDCx8_ASAP7_75t_R g1105 ( 
.A(n_904),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_961),
.A2(n_967),
.B(n_1027),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_999),
.A2(n_932),
.B(n_1011),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_956),
.A2(n_1011),
.B(n_1010),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_935),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_930),
.B(n_945),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1008),
.A2(n_1010),
.B(n_1009),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_984),
.A2(n_875),
.B(n_964),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_958),
.A2(n_933),
.B(n_973),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_991),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_869),
.B(n_872),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_999),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_973),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_869),
.A2(n_872),
.A3(n_959),
.B(n_1002),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_962),
.B(n_1014),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1014),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_943),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1028),
.B(n_966),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_917),
.B(n_857),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1002),
.A2(n_692),
.B(n_1032),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_901),
.A2(n_692),
.B(n_929),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1030),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_914),
.B(n_761),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_877),
.B(n_793),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1031),
.B(n_755),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1030),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_991),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_877),
.B(n_819),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1136)
);

OAI22x1_ASAP7_75t_L g1137 ( 
.A1(n_965),
.A2(n_987),
.B1(n_1017),
.B2(n_487),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1032),
.A2(n_692),
.B(n_926),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_1030),
.B(n_1020),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_971),
.B(n_975),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1030),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_929),
.A2(n_692),
.B(n_889),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1032),
.A2(n_692),
.B(n_926),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1034),
.B(n_755),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_914),
.B(n_761),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_971),
.B(n_975),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1030),
.B(n_1020),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1031),
.B(n_755),
.Y(n_1151)
);

BUFx12f_ASAP7_75t_L g1152 ( 
.A(n_904),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1031),
.B(n_755),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_894),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_971),
.B(n_975),
.Y(n_1157)
);

AND3x4_ASAP7_75t_L g1158 ( 
.A(n_885),
.B(n_992),
.C(n_1030),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_999),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_911),
.A2(n_696),
.B(n_1029),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_991),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_911),
.A2(n_696),
.B(n_1029),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_982),
.A2(n_997),
.B(n_993),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1030),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_L g1166 ( 
.A(n_993),
.B(n_755),
.Y(n_1166)
);

AO22x1_ASAP7_75t_L g1167 ( 
.A1(n_990),
.A2(n_987),
.B1(n_965),
.B2(n_1017),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1016),
.B(n_831),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1017),
.A2(n_990),
.B(n_1031),
.C(n_965),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_991),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1032),
.A2(n_692),
.B(n_926),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1017),
.A2(n_993),
.B(n_1012),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1034),
.B(n_755),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1034),
.B(n_755),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_SL g1178 ( 
.A1(n_946),
.A2(n_550),
.B(n_755),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_944),
.A2(n_881),
.B(n_912),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_882),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_911),
.A2(n_696),
.B(n_1029),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_911),
.A2(n_696),
.B(n_1029),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_991),
.Y(n_1183)
);

CKINVDCx14_ASAP7_75t_R g1184 ( 
.A(n_870),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1129),
.B(n_1146),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1041),
.A2(n_1141),
.B1(n_1169),
.B2(n_1136),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1049),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1174),
.A2(n_1137),
.B1(n_1080),
.B2(n_1040),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1037),
.A2(n_1055),
.B(n_1057),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1164),
.Y(n_1191)
);

OAI321xp33_ASAP7_75t_L g1192 ( 
.A1(n_1150),
.A2(n_1154),
.A3(n_1171),
.B1(n_1040),
.B2(n_1037),
.C(n_1043),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1164),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1059),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1128),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1062),
.B(n_1167),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_SL g1198 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1198)
);

OR2x4_ASAP7_75t_L g1199 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_L g1200 ( 
.A(n_1121),
.B(n_1071),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1087),
.B(n_1130),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1063),
.B(n_1042),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1159),
.B(n_1118),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1153),
.B(n_1174),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1087),
.B(n_1184),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1123),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1132),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1180),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1088),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1157),
.B(n_1139),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1065),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1052),
.B(n_1039),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1088),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1133),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1038),
.A2(n_1082),
.B(n_1114),
.C(n_1054),
.Y(n_1216)
);

BUFx12f_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

BUFx2_ASAP7_75t_R g1218 ( 
.A(n_1105),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1142),
.B(n_1103),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1139),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1079),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1152),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1139),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1148),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1068),
.B(n_1072),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1046),
.A2(n_1156),
.B(n_1165),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1148),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1125),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1133),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1052),
.B(n_1039),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_1157),
.B1(n_1102),
.B2(n_1086),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1119),
.A2(n_1176),
.B1(n_1175),
.B2(n_1145),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1148),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1076),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1125),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1094),
.B(n_1053),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1161),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1058),
.B(n_1036),
.Y(n_1238)
);

INVx4_ASAP7_75t_SL g1239 ( 
.A(n_1161),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_1099),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1110),
.B(n_1135),
.Y(n_1241)
);

INVx3_ASAP7_75t_SL g1242 ( 
.A(n_1124),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1168),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1070),
.B(n_1158),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1161),
.B(n_1183),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1182),
.A2(n_1054),
.B(n_1051),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1074),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1145),
.A2(n_1175),
.B1(n_1176),
.B2(n_1073),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1107),
.B(n_1172),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1122),
.B(n_1100),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1085),
.Y(n_1251)
);

OR2x6_ASAP7_75t_SL g1252 ( 
.A(n_1036),
.B(n_1117),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1124),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1183),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_SL g1255 ( 
.A(n_1092),
.B(n_1061),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1116),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1091),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1116),
.Y(n_1258)
);

BUFx4_ASAP7_75t_SL g1259 ( 
.A(n_1127),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1138),
.A2(n_1173),
.B(n_1144),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1112),
.B(n_1073),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1138),
.A2(n_1144),
.B(n_1173),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1178),
.A2(n_1064),
.B(n_1045),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1084),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1045),
.A2(n_1166),
.B(n_1112),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1155),
.B(n_1077),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1104),
.A2(n_1115),
.B1(n_1126),
.B2(n_1106),
.Y(n_1267)
);

BUFx4_ASAP7_75t_SL g1268 ( 
.A(n_1078),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1096),
.A2(n_1117),
.B1(n_1089),
.B2(n_1111),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1120),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1115),
.B(n_1113),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1126),
.A2(n_1082),
.B1(n_1114),
.B2(n_1067),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1098),
.A2(n_1048),
.B(n_1044),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1066),
.B1(n_1093),
.B2(n_1083),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1047),
.A2(n_1090),
.B(n_1081),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1109),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1093),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1050),
.B(n_1060),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1060),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1143),
.B(n_1134),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1179),
.B(n_1149),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1170),
.A2(n_1177),
.B(n_1163),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1136),
.B(n_774),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1049),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1049),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_L g1286 ( 
.A1(n_1167),
.A2(n_1136),
.B(n_1150),
.C(n_1141),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1132),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1059),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1137),
.A2(n_735),
.B1(n_1012),
.B2(n_883),
.Y(n_1291)
);

BUFx4_ASAP7_75t_SL g1292 ( 
.A(n_1056),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1059),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1136),
.B(n_1141),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1049),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1101),
.B(n_999),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1129),
.B(n_1146),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1059),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1130),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1049),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1302)
);

AOI21xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1137),
.A2(n_1167),
.B(n_535),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1136),
.A2(n_1141),
.B(n_1154),
.C(n_1150),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1059),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1130),
.B(n_853),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1136),
.A2(n_1141),
.B(n_1154),
.C(n_1150),
.Y(n_1310)
);

CKINVDCx6p67_ASAP7_75t_R g1311 ( 
.A(n_1069),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1129),
.B(n_1146),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1075),
.Y(n_1314)
);

INVx5_ASAP7_75t_L g1315 ( 
.A(n_1101),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1133),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1037),
.A2(n_1055),
.B(n_1057),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1160),
.A2(n_1181),
.B(n_1162),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1131),
.B(n_1151),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1191),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1187),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1219),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1282),
.A2(n_1226),
.B(n_1275),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1284),
.Y(n_1324)
);

INVx3_ASAP7_75t_SL g1325 ( 
.A(n_1314),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1285),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1287),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1242),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1194),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1294),
.A2(n_1283),
.B1(n_1291),
.B2(n_1186),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1228),
.B(n_1235),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1294),
.A2(n_1199),
.B1(n_1303),
.B2(n_1186),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1217),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1193),
.B(n_1300),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1199),
.A2(n_1231),
.B1(n_1189),
.B2(n_1197),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1306),
.B(n_1205),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1205),
.B(n_1319),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1288),
.Y(n_1338)
);

NAND2x1_ASAP7_75t_L g1339 ( 
.A(n_1276),
.B(n_1266),
.Y(n_1339)
);

INVx6_ASAP7_75t_L g1340 ( 
.A(n_1315),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1244),
.A2(n_1203),
.B1(n_1255),
.B2(n_1200),
.Y(n_1341)
);

AO21x1_ASAP7_75t_L g1342 ( 
.A1(n_1255),
.A2(n_1310),
.B(n_1272),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1222),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1209),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1258),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1191),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1190),
.A2(n_1317),
.B1(n_1225),
.B2(n_1243),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1207),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1319),
.B(n_1193),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1295),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1201),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1279),
.B(n_1315),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1301),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1299),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1188),
.Y(n_1355)
);

INVx6_ASAP7_75t_L g1356 ( 
.A(n_1315),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1221),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1192),
.A2(n_1302),
.B1(n_1304),
.B2(n_1300),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1212),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1247),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1315),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1195),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1251),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1296),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1277),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1308),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1257),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1238),
.A2(n_1230),
.B(n_1213),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1188),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1293),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1202),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1234),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1264),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1260),
.B(n_1262),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1264),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1228),
.B(n_1235),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1263),
.A2(n_1246),
.B(n_1318),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1185),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1297),
.A2(n_1313),
.B1(n_1309),
.B2(n_1305),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1250),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1311),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1289),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1261),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1250),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1239),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1236),
.Y(n_1388)
);

BUFx4_ASAP7_75t_R g1389 ( 
.A(n_1210),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1252),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1240),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1281),
.A2(n_1274),
.B(n_1265),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1206),
.A2(n_1272),
.B1(n_1232),
.B2(n_1223),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1202),
.B(n_1312),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1211),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1270),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1216),
.A2(n_1192),
.B(n_1274),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1232),
.A2(n_1248),
.B(n_1278),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1289),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1271),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1213),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1204),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1230),
.B(n_1278),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1267),
.A2(n_1286),
.B(n_1280),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1248),
.B(n_1269),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1211),
.B(n_1224),
.Y(n_1406)
);

BUFx2_ASAP7_75t_R g1407 ( 
.A(n_1253),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1220),
.B(n_1227),
.Y(n_1408)
);

BUFx2_ASAP7_75t_R g1409 ( 
.A(n_1214),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1249),
.B(n_1290),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1249),
.B(n_1290),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1268),
.A2(n_1259),
.B(n_1312),
.Y(n_1412)
);

BUFx2_ASAP7_75t_R g1413 ( 
.A(n_1233),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1292),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1254),
.A2(n_1241),
.B(n_1208),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1298),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1241),
.A2(n_1198),
.B1(n_1196),
.B2(n_1256),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1307),
.A2(n_1256),
.B1(n_1215),
.B2(n_1237),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1316),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1245),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1316),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1239),
.Y(n_1422)
);

NAND2x1p5_ASAP7_75t_L g1423 ( 
.A(n_1215),
.B(n_1229),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1316),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1239),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1229),
.A2(n_1237),
.B(n_1218),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1187),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1294),
.A2(n_1041),
.B1(n_1137),
.B2(n_1186),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1219),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1217),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1286),
.A2(n_1141),
.B(n_1136),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1187),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1294),
.A2(n_1041),
.B1(n_1137),
.B2(n_1186),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1282),
.A2(n_1226),
.B(n_1275),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1187),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1217),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1217),
.Y(n_1437)
);

BUFx2_ASAP7_75t_R g1438 ( 
.A(n_1314),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1286),
.A2(n_1141),
.B(n_1136),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1190),
.A2(n_1317),
.B(n_1273),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1199),
.A2(n_1136),
.B1(n_1150),
.B2(n_1141),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1282),
.A2(n_1263),
.B(n_1275),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1315),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1294),
.A2(n_1041),
.B1(n_1137),
.B2(n_1186),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1294),
.A2(n_1012),
.B1(n_735),
.B2(n_1199),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1415),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1349),
.B(n_1366),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1346),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1323),
.A2(n_1434),
.B(n_1442),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1323),
.A2(n_1434),
.B(n_1442),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1414),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1396),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1337),
.B(n_1400),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1339),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1415),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1339),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1337),
.B(n_1400),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1329),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1398),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1396),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1398),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1375),
.B(n_1342),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1415),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1428),
.A2(n_1444),
.B1(n_1433),
.B2(n_1330),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1405),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1405),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1383),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1403),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1357),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1329),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1331),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1431),
.A2(n_1439),
.B(n_1441),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1336),
.B(n_1349),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1332),
.B(n_1367),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1440),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1336),
.B(n_1388),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1440),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1320),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1440),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1375),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1365),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1378),
.A2(n_1392),
.B(n_1342),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1445),
.B(n_1394),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1375),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1366),
.B(n_1386),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1386),
.B(n_1322),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1335),
.A2(n_1347),
.B1(n_1341),
.B2(n_1393),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1378),
.A2(n_1397),
.B(n_1369),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1397),
.A2(n_1358),
.B(n_1353),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1322),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1352),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1374),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1429),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1334),
.B(n_1380),
.Y(n_1495)
);

AOI21xp33_ASAP7_75t_L g1496 ( 
.A1(n_1397),
.A2(n_1391),
.B(n_1381),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1351),
.B(n_1384),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1344),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1383),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1331),
.B(n_1377),
.Y(n_1500)
);

AOI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1404),
.A2(n_1390),
.B(n_1402),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1429),
.B(n_1390),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1443),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1426),
.A2(n_1361),
.B(n_1401),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1350),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1360),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1443),
.B(n_1361),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1363),
.A2(n_1368),
.B(n_1373),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1432),
.B(n_1379),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1376),
.B(n_1385),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1321),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1324),
.Y(n_1512)
);

NAND2x1_ASAP7_75t_L g1513 ( 
.A(n_1340),
.B(n_1356),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1326),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1414),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1427),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1435),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1443),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1377),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1377),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1340),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1364),
.A2(n_1423),
.B(n_1425),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1417),
.A2(n_1354),
.B(n_1359),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1340),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1340),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1356),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1356),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1356),
.Y(n_1530)
);

INVx5_ASAP7_75t_SL g1531 ( 
.A(n_1412),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1419),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1455),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1465),
.A2(n_1412),
.B1(n_1406),
.B2(n_1372),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1463),
.B(n_1412),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1463),
.B(n_1406),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1463),
.B(n_1424),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1476),
.A2(n_1421),
.B(n_1408),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1481),
.B(n_1485),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1446),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1463),
.B(n_1395),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1463),
.B(n_1478),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1480),
.B(n_1327),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1481),
.B(n_1485),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1464),
.B(n_1408),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1473),
.A2(n_1488),
.B1(n_1475),
.B2(n_1484),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1327),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1488),
.A2(n_1343),
.B1(n_1389),
.B2(n_1382),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1489),
.B(n_1420),
.Y(n_1549)
);

NAND2xp33_ASAP7_75t_SL g1550 ( 
.A(n_1513),
.B(n_1389),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1489),
.B(n_1483),
.Y(n_1551)
);

AND2x4_ASAP7_75t_SL g1552 ( 
.A(n_1503),
.B(n_1518),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1460),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1525),
.A2(n_1418),
.B(n_1364),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1483),
.B(n_1466),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1483),
.B(n_1466),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1469),
.B(n_1420),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1558)
);

OAI222xp33_ASAP7_75t_L g1559 ( 
.A1(n_1495),
.A2(n_1382),
.B1(n_1364),
.B2(n_1355),
.C1(n_1372),
.C2(n_1370),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1462),
.B(n_1453),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1459),
.B(n_1370),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1515),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1508),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1453),
.B(n_1419),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1457),
.B(n_1474),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1459),
.B(n_1355),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1457),
.B(n_1423),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1474),
.B(n_1423),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1469),
.B(n_1422),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1454),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1454),
.B(n_1345),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1468),
.A2(n_1345),
.B(n_1338),
.Y(n_1572)
);

NAND2x1_ASAP7_75t_L g1573 ( 
.A(n_1454),
.B(n_1456),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1565),
.B(n_1482),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1546),
.B(n_1482),
.C(n_1496),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1565),
.B(n_1448),
.Y(n_1576)
);

AOI211xp5_ASAP7_75t_L g1577 ( 
.A1(n_1554),
.A2(n_1572),
.B(n_1559),
.C(n_1535),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1546),
.A2(n_1490),
.B1(n_1502),
.B2(n_1477),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1548),
.A2(n_1524),
.B(n_1504),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1548),
.B(n_1521),
.C(n_1502),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1554),
.A2(n_1470),
.B1(n_1499),
.B2(n_1468),
.C(n_1513),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_1487),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1534),
.B(n_1521),
.C(n_1493),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1534),
.B(n_1522),
.C(n_1492),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1560),
.B(n_1501),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1535),
.A2(n_1559),
.B(n_1536),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1547),
.B(n_1522),
.C(n_1492),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1547),
.B(n_1529),
.C(n_1530),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1529),
.C(n_1530),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1567),
.B(n_1491),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1447),
.Y(n_1591)
);

NAND4xp25_ASAP7_75t_L g1592 ( 
.A(n_1569),
.B(n_1479),
.C(n_1497),
.D(n_1510),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1544),
.A2(n_1458),
.B1(n_1471),
.B2(n_1477),
.C(n_1494),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1535),
.A2(n_1486),
.B1(n_1494),
.B2(n_1491),
.C(n_1520),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_R g1595 ( 
.A(n_1550),
.B(n_1451),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1523),
.C(n_1526),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1562),
.A2(n_1490),
.B1(n_1477),
.B2(n_1500),
.Y(n_1597)
);

OAI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1561),
.A2(n_1499),
.B1(n_1523),
.B2(n_1528),
.C(n_1526),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1543),
.B(n_1498),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1551),
.B(n_1545),
.C(n_1569),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1543),
.B(n_1498),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1551),
.B(n_1528),
.C(n_1477),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1544),
.A2(n_1509),
.B1(n_1510),
.B2(n_1516),
.C(n_1506),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1563),
.A2(n_1449),
.B(n_1450),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1560),
.B(n_1543),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1571),
.B(n_1472),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1567),
.B(n_1505),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1536),
.A2(n_1519),
.B(n_1520),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1564),
.B(n_1568),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1564),
.B(n_1506),
.Y(n_1612)
);

NAND4xp25_ASAP7_75t_L g1613 ( 
.A(n_1545),
.B(n_1516),
.C(n_1514),
.D(n_1517),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1551),
.B(n_1545),
.C(n_1561),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1452),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1561),
.B(n_1566),
.C(n_1549),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1568),
.B(n_1461),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1558),
.B(n_1511),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1571),
.A2(n_1519),
.B(n_1500),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1537),
.B(n_1531),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1544),
.B(n_1531),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1566),
.A2(n_1451),
.B1(n_1325),
.B2(n_1338),
.C(n_1553),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1558),
.B(n_1512),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1574),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1605),
.B(n_1540),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1621),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1585),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1605),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1555),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1614),
.B(n_1538),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1591),
.B(n_1555),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1599),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1538),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1580),
.A2(n_1539),
.B1(n_1571),
.B2(n_1541),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1619),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1624),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1538),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1612),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1582),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1577),
.B(n_1571),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1604),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1571),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1606),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1587),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1606),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1538),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1622),
.B(n_1549),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1602),
.B(n_1573),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1617),
.B(n_1533),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1621),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1622),
.B(n_1570),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1603),
.B(n_1556),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1611),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1645),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1645),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1658),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1654),
.B(n_1609),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1646),
.A2(n_1586),
.B1(n_1581),
.B2(n_1575),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1654),
.B(n_1609),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1662),
.B(n_1590),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1657),
.B(n_1579),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1662),
.B(n_1592),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1627),
.B(n_1620),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1650),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1597),
.Y(n_1677)
);

OAI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1651),
.A2(n_1578),
.B(n_1597),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1593),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1627),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1629),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1665),
.B(n_1610),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1629),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1632),
.B(n_1578),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1641),
.B(n_1549),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1635),
.B(n_1566),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1552),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1641),
.B(n_1539),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1552),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1630),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1631),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1648),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1657),
.B(n_1596),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1650),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1642),
.B(n_1539),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1642),
.B(n_1539),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1655),
.B(n_1533),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1652),
.B(n_1539),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1638),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1628),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1639),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1674),
.B(n_1664),
.Y(n_1706)
);

O2A1O1Ixp33_ASAP7_75t_SL g1707 ( 
.A1(n_1702),
.A2(n_1562),
.B(n_1664),
.C(n_1633),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

AOI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1678),
.A2(n_1583),
.B(n_1584),
.C(n_1633),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1667),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1681),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1713)
);

NOR2xp67_ASAP7_75t_L g1714 ( 
.A(n_1702),
.B(n_1639),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1688),
.B(n_1653),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1674),
.B(n_1644),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1688),
.B(n_1663),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1668),
.B(n_1643),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1691),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1670),
.A2(n_1634),
.B(n_1640),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1703),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1673),
.B(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1693),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1673),
.B(n_1660),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_SL g1730 ( 
.A(n_1684),
.B(n_1343),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1676),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1676),
.Y(n_1735)
);

INVxp33_ASAP7_75t_L g1736 ( 
.A(n_1672),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1695),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1694),
.B(n_1636),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1695),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1696),
.B(n_1643),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1673),
.B(n_1661),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1697),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1696),
.B(n_1655),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1680),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1697),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1700),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1700),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1677),
.B(n_1634),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1686),
.Y(n_1749)
);

NAND2x1_ASAP7_75t_L g1750 ( 
.A(n_1731),
.B(n_1673),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1661),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1729),
.B(n_1687),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1744),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1708),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1731),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1717),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1669),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1706),
.B(n_1671),
.Y(n_1759)
);

AND3x2_ASAP7_75t_L g1760 ( 
.A(n_1709),
.B(n_1704),
.C(n_1705),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1726),
.Y(n_1762)
);

AND3x1_ASAP7_75t_L g1763 ( 
.A(n_1709),
.B(n_1731),
.C(n_1723),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1731),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1736),
.B(n_1636),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1708),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1726),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1738),
.B(n_1637),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1730),
.B(n_1430),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1730),
.A2(n_1595),
.B1(n_1531),
.B2(n_1705),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1710),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1713),
.B(n_1638),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1710),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1637),
.Y(n_1775)
);

NOR2xp67_ASAP7_75t_L g1776 ( 
.A(n_1714),
.B(n_1734),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1727),
.B(n_1689),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1712),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1728),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1712),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1718),
.B(n_1626),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1716),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1728),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1714),
.B(n_1625),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1718),
.B(n_1626),
.Y(n_1785)
);

AO22x1_ASAP7_75t_L g1786 ( 
.A1(n_1764),
.A2(n_1734),
.B1(n_1333),
.B2(n_1741),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1763),
.A2(n_1707),
.B1(n_1734),
.B2(n_1743),
.C(n_1746),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1754),
.B(n_1783),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_SL g1789 ( 
.A(n_1784),
.B(n_1743),
.C(n_1740),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1778),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1755),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1779),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1750),
.A2(n_1740),
.B(n_1748),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1755),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1766),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1756),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1760),
.A2(n_1734),
.B1(n_1748),
.B2(n_1741),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1766),
.Y(n_1799)
);

OAI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1763),
.A2(n_1749),
.B1(n_1747),
.B2(n_1746),
.C(n_1719),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1772),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1779),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1752),
.B(n_1720),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1776),
.A2(n_1747),
.B(n_1722),
.C(n_1720),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1776),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1753),
.Y(n_1806)
);

CKINVDCx16_ASAP7_75t_R g1807 ( 
.A(n_1770),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1756),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1772),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1753),
.Y(n_1810)
);

AOI31xp33_ASAP7_75t_L g1811 ( 
.A1(n_1771),
.A2(n_1438),
.A3(n_1328),
.B(n_1407),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1796),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1788),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1808),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1792),
.B(n_1762),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1791),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1796),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1802),
.B(n_1767),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1791),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1806),
.B(n_1759),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1789),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1803),
.B(n_1752),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1803),
.B(n_1781),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1787),
.A2(n_1768),
.B(n_1758),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1790),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1794),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1810),
.B(n_1758),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1800),
.B(n_1750),
.C(n_1756),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1798),
.B(n_1769),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1805),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_SL g1832 ( 
.A(n_1821),
.B(n_1797),
.C(n_1804),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1825),
.A2(n_1797),
.B(n_1793),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1815),
.B(n_1777),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1813),
.B(n_1786),
.C(n_1795),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1813),
.A2(n_1786),
.B1(n_1768),
.B2(n_1751),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_SL g1837 ( 
.A(n_1829),
.B(n_1799),
.C(n_1801),
.D(n_1809),
.Y(n_1837)
);

AOI32xp33_ASAP7_75t_L g1838 ( 
.A1(n_1820),
.A2(n_1751),
.A3(n_1774),
.B1(n_1782),
.B2(n_1780),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1822),
.A2(n_1773),
.B1(n_1765),
.B2(n_1774),
.Y(n_1839)
);

AOI221x1_ASAP7_75t_L g1840 ( 
.A1(n_1831),
.A2(n_1780),
.B1(n_1782),
.B2(n_1761),
.C(n_1775),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1831),
.B(n_1362),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1814),
.B(n_1761),
.C(n_1781),
.D(n_1785),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1814),
.Y(n_1843)
);

AO22x2_ASAP7_75t_L g1844 ( 
.A1(n_1832),
.A2(n_1824),
.B1(n_1826),
.B2(n_1819),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_SL g1845 ( 
.A1(n_1833),
.A2(n_1818),
.B(n_1817),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1835),
.B(n_1820),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1843),
.B(n_1828),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1841),
.B(n_1838),
.C(n_1828),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1836),
.B(n_1822),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1837),
.B(n_1812),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_SL g1851 ( 
.A(n_1842),
.B(n_1827),
.C(n_1816),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

NAND4xp25_ASAP7_75t_L g1853 ( 
.A(n_1834),
.B(n_1830),
.C(n_1817),
.D(n_1812),
.Y(n_1853)
);

NAND4xp25_ASAP7_75t_L g1854 ( 
.A(n_1839),
.B(n_1823),
.C(n_1773),
.D(n_1722),
.Y(n_1854)
);

OAI21x1_ASAP7_75t_L g1855 ( 
.A1(n_1850),
.A2(n_1852),
.B(n_1845),
.Y(n_1855)
);

AOI211xp5_ASAP7_75t_L g1856 ( 
.A1(n_1846),
.A2(n_1325),
.B(n_1773),
.C(n_1333),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1844),
.A2(n_1773),
.B1(n_1732),
.B2(n_1724),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1847),
.B(n_1719),
.Y(n_1858)
);

AOI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1848),
.A2(n_1333),
.B(n_1811),
.C(n_1436),
.Y(n_1859)
);

OAI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1851),
.A2(n_1430),
.B(n_1437),
.C(n_1436),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1853),
.B(n_1437),
.C(n_1724),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1844),
.A2(n_1732),
.B(n_1716),
.C(n_1725),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1859),
.A2(n_1849),
.B1(n_1721),
.B2(n_1725),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_L g1864 ( 
.A(n_1860),
.B(n_1854),
.C(n_1348),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1858),
.Y(n_1865)
);

AND3x4_ASAP7_75t_L g1866 ( 
.A(n_1861),
.B(n_1348),
.C(n_1413),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1855),
.B(n_1362),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1857),
.B(n_1856),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1862),
.B(n_1785),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1865),
.B(n_1721),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1864),
.A2(n_1732),
.B1(n_1735),
.B2(n_1739),
.C(n_1742),
.Y(n_1871)
);

NOR2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1869),
.B(n_1399),
.Y(n_1872)
);

INVx3_ASAP7_75t_SL g1873 ( 
.A(n_1868),
.Y(n_1873)
);

AND3x4_ASAP7_75t_L g1874 ( 
.A(n_1866),
.B(n_1399),
.C(n_1409),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_SL g1875 ( 
.A(n_1867),
.B(n_1371),
.C(n_1416),
.Y(n_1875)
);

XOR2x2_ASAP7_75t_L g1876 ( 
.A(n_1874),
.B(n_1863),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1873),
.A2(n_1735),
.B1(n_1742),
.B2(n_1739),
.Y(n_1877)
);

OR3x2_ASAP7_75t_L g1878 ( 
.A(n_1870),
.B(n_1416),
.C(n_1371),
.Y(n_1878)
);

XOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1878),
.B(n_1875),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_L g1880 ( 
.A(n_1879),
.B(n_1876),
.C(n_1872),
.Y(n_1880)
);

AOI22x1_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1877),
.B1(n_1871),
.B2(n_1739),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1880),
.A2(n_1742),
.B(n_1735),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1881),
.A2(n_1745),
.B1(n_1737),
.B2(n_1733),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1882),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1884),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1883),
.A2(n_1745),
.B1(n_1737),
.B2(n_1733),
.C(n_1715),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1885),
.A2(n_1598),
.B(n_1507),
.Y(n_1887)
);

AOI322xp5_ASAP7_75t_L g1888 ( 
.A1(n_1887),
.A2(n_1886),
.A3(n_1685),
.B1(n_1701),
.B2(n_1699),
.C1(n_1698),
.C2(n_1638),
.Y(n_1888)
);

OAI221xp5_ASAP7_75t_R g1889 ( 
.A1(n_1888),
.A2(n_1387),
.B1(n_1531),
.B2(n_1647),
.C(n_1649),
.Y(n_1889)
);

AOI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1889),
.A2(n_1527),
.B(n_1532),
.C(n_1647),
.Y(n_1890)
);


endmodule