module real_aes_8734_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_162;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_1), .A2(n_139), .B(n_143), .C(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_2), .A2(n_173), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g513 ( .A(n_3), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_4), .B(n_240), .Y(n_259) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_173), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g139 ( .A(n_6), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g214 ( .A(n_7), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_42), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_9), .A2(n_172), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_10), .B(n_151), .Y(n_226) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_12), .B(n_254), .Y(n_538) );
INVx1_ASAP7_75t_L g159 ( .A(n_13), .Y(n_159) );
INVx1_ASAP7_75t_L g550 ( .A(n_14), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_15), .A2(n_149), .B(n_236), .C(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_16), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_17), .B(n_501), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_18), .B(n_173), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_19), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_20), .A2(n_254), .B(n_269), .C(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_21), .B(n_240), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_22), .B(n_151), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_23), .A2(n_181), .B(n_238), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_24), .B(n_151), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_25), .Y(n_190) );
INVx1_ASAP7_75t_L g147 ( .A(n_26), .Y(n_147) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_28), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_29), .B(n_151), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_30), .A2(n_31), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_30), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_31), .Y(n_748) );
INVx1_ASAP7_75t_L g179 ( .A(n_32), .Y(n_179) );
INVx1_ASAP7_75t_L g492 ( .A(n_33), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_34), .A2(n_104), .B1(n_117), .B2(n_757), .Y(n_103) );
INVx2_ASAP7_75t_L g137 ( .A(n_35), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_36), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_37), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
INVxp67_ASAP7_75t_L g180 ( .A(n_38), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_39), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_40), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_41), .A2(n_139), .B(n_143), .C(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g491 ( .A(n_43), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_44), .A2(n_198), .B(n_212), .C(n_213), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_45), .B(n_151), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_46), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_46), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_47), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_48), .Y(n_175) );
INVx1_ASAP7_75t_L g267 ( .A(n_49), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_50), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_51), .B(n_173), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_52), .B(n_459), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_53), .A2(n_143), .B1(n_271), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_54), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_55), .Y(n_510) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_56), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_212), .B(n_257), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_58), .Y(n_566) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_60), .A2(n_89), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_60), .Y(n_454) );
INVx1_ASAP7_75t_L g140 ( .A(n_61), .Y(n_140) );
INVx1_ASAP7_75t_L g158 ( .A(n_62), .Y(n_158) );
INVx1_ASAP7_75t_SL g256 ( .A(n_63), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_65), .B(n_240), .Y(n_273) );
INVx1_ASAP7_75t_L g193 ( .A(n_66), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_67), .A2(n_257), .B(n_501), .C(n_502), .Y(n_500) );
INVxp67_ASAP7_75t_L g503 ( .A(n_68), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_69), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_69), .Y(n_124) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_71), .A2(n_173), .B(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_72), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_73), .A2(n_173), .B(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_74), .Y(n_495) );
INVx1_ASAP7_75t_L g560 ( .A(n_75), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_76), .A2(n_172), .B(n_174), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_77), .Y(n_141) );
INVx1_ASAP7_75t_L g234 ( .A(n_78), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_79), .A2(n_139), .B(n_143), .C(n_562), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_80), .A2(n_173), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g237 ( .A(n_81), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_82), .B(n_148), .Y(n_526) );
INVx2_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
INVx1_ASAP7_75t_L g225 ( .A(n_84), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_85), .B(n_501), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_86), .A2(n_139), .B(n_143), .C(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OR2x2_ASAP7_75t_L g457 ( .A(n_87), .B(n_113), .Y(n_457) );
OR2x2_ASAP7_75t_L g466 ( .A(n_87), .B(n_114), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_88), .A2(n_143), .B(n_192), .C(n_200), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_89), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_90), .B(n_155), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_91), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_92), .A2(n_139), .B(n_143), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_93), .Y(n_542) );
INVx1_ASAP7_75t_L g499 ( .A(n_94), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_95), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_96), .B(n_148), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_97), .B(n_163), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_98), .B(n_163), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_99), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g270 ( .A(n_100), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_101), .A2(n_173), .B(n_498), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_102), .A2(n_463), .B1(n_744), .B2(n_745), .C1(n_751), .C2(n_754), .Y(n_462) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g757 ( .A(n_107), .Y(n_757) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_SL g754 ( .A(n_110), .Y(n_754) );
INVx3_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
NOR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g469 ( .A(n_112), .B(n_114), .Y(n_469) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_461), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g756 ( .A(n_120), .Y(n_756) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_455), .B(n_458), .Y(n_122) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_452), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_127), .A2(n_464), .B1(n_467), .B2(n_470), .Y(n_463) );
INVx1_ASAP7_75t_L g752 ( .A(n_127), .Y(n_752) );
OR4x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_342), .C(n_389), .D(n_429), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_288), .C(n_317), .Y(n_128) );
AOI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_203), .B(n_241), .C(n_281), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_130), .A2(n_301), .B(n_318), .C(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_132), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_SL g284 ( .A(n_132), .Y(n_284) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_132), .Y(n_296) );
AND2x4_ASAP7_75t_L g300 ( .A(n_132), .B(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_132), .B(n_188), .Y(n_311) );
OR2x2_ASAP7_75t_L g335 ( .A(n_132), .B(n_244), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_132), .B(n_249), .Y(n_348) );
AND2x2_ASAP7_75t_L g388 ( .A(n_132), .B(n_374), .Y(n_388) );
AND2x2_ASAP7_75t_L g395 ( .A(n_132), .B(n_358), .Y(n_395) );
AND2x2_ASAP7_75t_L g425 ( .A(n_132), .B(n_166), .Y(n_425) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_160), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_142), .C(n_155), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_134), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_134), .A2(n_222), .B(n_223), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_134), .A2(n_183), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_134), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_134), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
AND2x4_ASAP7_75t_L g173 ( .A(n_135), .B(n_139), .Y(n_173) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx1_ASAP7_75t_L g272 ( .A(n_137), .Y(n_272) );
INVx1_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_138), .Y(n_151) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
INVx1_ASAP7_75t_L g501 ( .A(n_138), .Y(n_501) );
BUFx3_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx4_ASAP7_75t_SL g183 ( .A(n_139), .Y(n_183) );
INVx5_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_144), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_152), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_148), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_148), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_149), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_149), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_149), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx4_ASAP7_75t_L g254 ( .A(n_151), .Y(n_254) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_153), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_155), .A2(n_208), .B(n_215), .Y(n_207) );
INVx1_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_155), .A2(n_545), .B(n_551), .Y(n_544) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g164 ( .A(n_156), .B(n_157), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_201), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_162), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_162), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_163), .Y(n_231) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_163), .A2(n_497), .B(n_504), .Y(n_496) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_165), .B(n_352), .Y(n_364) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_187), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_166), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g302 ( .A(n_166), .B(n_187), .Y(n_302) );
BUFx3_ASAP7_75t_L g310 ( .A(n_166), .Y(n_310) );
OR2x2_ASAP7_75t_L g331 ( .A(n_166), .B(n_206), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_166), .B(n_352), .Y(n_442) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_184), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_245), .B(n_246), .Y(n_244) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_168), .A2(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_169), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_170), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_170), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_170), .A2(n_509), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_176), .A2(n_183), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_176), .A2(n_183), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_176), .A2(n_183), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_176), .A2(n_183), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_176), .A2(n_183), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_176), .A2(n_183), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_176), .A2(n_183), .B(n_547), .C(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_181), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_181), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_181), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_182), .A2(n_195), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
INVx1_ASAP7_75t_L g246 ( .A(n_184), .Y(n_246) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_186), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_186), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_L g247 ( .A(n_187), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g295 ( .A(n_187), .Y(n_295) );
AND2x2_ASAP7_75t_L g358 ( .A(n_187), .B(n_249), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_187), .A2(n_361), .B1(n_363), .B2(n_365), .C(n_366), .Y(n_360) );
AND2x2_ASAP7_75t_L g374 ( .A(n_187), .B(n_244), .Y(n_374) );
AND2x2_ASAP7_75t_L g400 ( .A(n_187), .B(n_284), .Y(n_400) );
INVx2_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g280 ( .A(n_188), .B(n_249), .Y(n_280) );
BUFx2_ASAP7_75t_L g414 ( .A(n_188), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_194), .A2(n_197), .B(n_225), .C(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_197), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_197), .A2(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_204), .A2(n_341), .A3(n_355), .B1(n_381), .B2(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
AND2x2_ASAP7_75t_L g321 ( .A(n_205), .B(n_263), .Y(n_321) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g303 ( .A(n_206), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_206), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g375 ( .A(n_206), .B(n_263), .Y(n_375) );
AND2x2_ASAP7_75t_L g386 ( .A(n_206), .B(n_278), .Y(n_386) );
BUFx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g287 ( .A(n_207), .B(n_264), .Y(n_287) );
AND2x2_ASAP7_75t_L g291 ( .A(n_207), .B(n_264), .Y(n_291) );
AND2x2_ASAP7_75t_L g326 ( .A(n_207), .B(n_277), .Y(n_326) );
AND2x2_ASAP7_75t_L g333 ( .A(n_207), .B(n_229), .Y(n_333) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_207), .A2(n_284), .B(n_295), .C(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g392 ( .A(n_207), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_207), .B(n_218), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_275), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_216), .B(n_291), .Y(n_381) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g286 ( .A(n_217), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
AND2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_230), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_218), .B(n_230), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_218), .B(n_277), .Y(n_316) );
INVx1_ASAP7_75t_L g320 ( .A(n_218), .Y(n_320) );
AND2x2_ASAP7_75t_L g339 ( .A(n_218), .B(n_276), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_218), .A2(n_304), .B1(n_350), .B2(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_218), .B(n_392), .Y(n_416) );
AND2x2_ASAP7_75t_L g431 ( .A(n_218), .B(n_291), .Y(n_431) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx3_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
AND2x2_ASAP7_75t_L g305 ( .A(n_219), .B(n_230), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_219), .B(n_263), .Y(n_307) );
AND3x2_ASAP7_75t_L g369 ( .A(n_219), .B(n_333), .C(n_370), .Y(n_369) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_220), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_220), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_220), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g404 ( .A(n_229), .B(n_276), .Y(n_404) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g263 ( .A(n_230), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_230), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_230), .B(n_275), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_230), .B(n_316), .C(n_392), .Y(n_444) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_239), .Y(n_230) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_231), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_231), .A2(n_265), .B(n_273), .Y(n_264) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_240), .A2(n_478), .B(n_484), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_260), .B1(n_274), .B2(n_279), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_244), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g356 ( .A(n_244), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_247), .A2(n_373), .A3(n_374), .B(n_375), .Y(n_372) );
AND2x2_ASAP7_75t_L g397 ( .A(n_247), .B(n_284), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_247), .B(n_310), .Y(n_443) );
AND2x2_ASAP7_75t_L g352 ( .A(n_248), .B(n_284), .Y(n_352) );
AND2x2_ASAP7_75t_L g413 ( .A(n_248), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g283 ( .A(n_249), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g341 ( .A(n_249), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_258), .Y(n_539) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_261), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_262), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AOI221x1_ASAP7_75t_SL g329 ( .A1(n_263), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_336), .Y(n_329) );
INVx2_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_264), .Y(n_371) );
INVx2_ASAP7_75t_L g515 ( .A(n_271), .Y(n_515) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g359 ( .A(n_274), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_275), .B(n_292), .Y(n_384) );
INVx1_ASAP7_75t_SL g447 ( .A(n_275), .Y(n_447) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g365 ( .A(n_278), .B(n_291), .Y(n_365) );
INVx1_ASAP7_75t_L g433 ( .A(n_279), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_279), .B(n_362), .Y(n_446) );
INVx2_ASAP7_75t_SL g285 ( .A(n_280), .Y(n_285) );
AND2x2_ASAP7_75t_L g328 ( .A(n_280), .B(n_284), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_280), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_280), .B(n_355), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_285), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_283), .B(n_355), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_283), .B(n_310), .Y(n_451) );
OR2x2_ASAP7_75t_L g323 ( .A(n_284), .B(n_302), .Y(n_323) );
AND2x2_ASAP7_75t_L g422 ( .A(n_284), .B(n_413), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g297 ( .A1(n_285), .A2(n_298), .B1(n_303), .B2(n_306), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_285), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g409 ( .A(n_287), .Y(n_409) );
AOI311xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .A3(n_296), .B(n_297), .C(n_308), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_292), .A2(n_424), .B1(n_436), .B2(n_439), .C(n_441), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_292), .B(n_447), .Y(n_449) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_337), .B(n_338), .C(n_340), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_SL g405 ( .A1(n_299), .A2(n_301), .B(n_406), .C(n_407), .Y(n_405) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_300), .B(n_374), .Y(n_440) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_303), .A2(n_323), .B1(n_324), .B2(n_327), .C(n_329), .Y(n_322) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g408 ( .A(n_305), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_309), .A2(n_367), .B(n_368), .C(n_372), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_310), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_310), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_316), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_320), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g434 ( .A(n_323), .Y(n_434) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_326), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_326), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g438 ( .A(n_326), .Y(n_438) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g379 ( .A(n_328), .B(n_355), .Y(n_379) );
INVx1_ASAP7_75t_SL g373 ( .A(n_335), .Y(n_373) );
INVx1_ASAP7_75t_L g350 ( .A(n_341), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_360), .C(n_376), .Y(n_342) );
AOI322xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .A3(n_347), .B1(n_349), .B2(n_353), .C1(n_357), .C2(n_359), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_344), .A2(n_397), .B(n_398), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_347), .A2(n_368), .B1(n_399), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_355), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_355), .B(n_395), .Y(n_394) );
AOI32xp33_ASAP7_75t_L g445 ( .A1(n_355), .A2(n_446), .A3(n_447), .B1(n_448), .B2(n_450), .Y(n_445) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g367 ( .A(n_358), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_358), .A2(n_411), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_410) );
AND2x2_ASAP7_75t_L g424 ( .A(n_358), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g427 ( .A(n_362), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g437 ( .A(n_362), .B(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g428 ( .A(n_371), .B(n_392), .Y(n_428) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .C(n_383), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_393), .B(n_396), .C(n_410), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_404), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_416), .Y(n_419) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_426), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI211xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B(n_435), .C(n_445), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_457), .Y(n_460) );
AOI21xp33_ASAP7_75t_L g461 ( .A1(n_458), .A2(n_462), .B(n_755), .Y(n_461) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_464), .A2(n_467), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g753 ( .A(n_471), .Y(n_753) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_666), .C(n_711), .Y(n_472) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_589), .C(n_630), .D(n_647), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_505), .B(n_519), .C(n_552), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_476), .B(n_506), .Y(n_505) );
NOR4xp25_ASAP7_75t_L g613 ( .A(n_476), .B(n_607), .C(n_614), .D(n_620), .Y(n_613) );
AND2x2_ASAP7_75t_L g686 ( .A(n_476), .B(n_575), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_476), .B(n_651), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_476), .B(n_700), .Y(n_714) );
AND2x2_ASAP7_75t_L g727 ( .A(n_476), .B(n_518), .Y(n_727) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g572 ( .A(n_477), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_477), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g629 ( .A(n_477), .B(n_486), .Y(n_629) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_477), .B(n_575), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_477), .B(n_486), .Y(n_644) );
AND2x2_ASAP7_75t_L g653 ( .A(n_477), .B(n_578), .Y(n_653) );
BUFx2_ASAP7_75t_L g676 ( .A(n_477), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_477), .B(n_496), .Y(n_680) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_496), .Y(n_518) );
BUFx2_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_486), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g636 ( .A(n_486), .B(n_508), .Y(n_636) );
AND2x2_ASAP7_75t_L g700 ( .A(n_486), .B(n_578), .Y(n_700) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g568 ( .A(n_487), .B(n_508), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_487), .B(n_496), .Y(n_575) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_487), .Y(n_617) );
OR2x2_ASAP7_75t_L g652 ( .A(n_487), .B(n_507), .Y(n_652) );
INVx1_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
INVx3_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
BUFx2_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_496), .B(n_572), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_505), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_580), .Y(n_584) );
INVx1_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
INVx1_ASAP7_75t_L g590 ( .A(n_518), .Y(n_590) );
NAND2x1_ASAP7_75t_SL g519 ( .A(n_520), .B(n_530), .Y(n_519) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_543), .Y(n_588) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_520), .Y(n_662) );
AND2x2_ASAP7_75t_L g689 ( .A(n_520), .B(n_609), .Y(n_689) );
AND2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_659), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_520), .B(n_555), .Y(n_724) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g556 ( .A(n_521), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g573 ( .A(n_521), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g594 ( .A(n_521), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_521), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g633 ( .A(n_521), .B(n_558), .Y(n_633) );
OR2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_626), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g683 ( .A1(n_521), .A2(n_684), .A3(n_687), .B1(n_688), .B2(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_521), .B(n_659), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_521), .B(n_619), .Y(n_734) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_543), .Y(n_531) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_532), .B(n_557), .Y(n_626) );
AND2x2_ASAP7_75t_L g659 ( .A(n_532), .B(n_635), .Y(n_659) );
AND2x2_ASAP7_75t_L g696 ( .A(n_532), .B(n_558), .Y(n_696) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g555 ( .A(n_533), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_533), .B(n_557), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g634 ( .A(n_533), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g610 ( .A(n_543), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_543), .B(n_557), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_543), .B(n_601), .Y(n_682) );
INVx1_ASAP7_75t_L g704 ( .A(n_543), .Y(n_704) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_557), .Y(n_574) );
AND2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g635 ( .A(n_544), .Y(n_635) );
AOI221x1_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_567), .B1(n_573), .B2(n_575), .C(n_576), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_553), .A2(n_640), .B1(n_707), .B2(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g693 ( .A(n_554), .B(n_573), .Y(n_693) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_574), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
AND2x2_ASAP7_75t_L g672 ( .A(n_556), .B(n_659), .Y(n_672) );
AND2x2_ASAP7_75t_L g739 ( .A(n_556), .B(n_634), .Y(n_739) );
INVx2_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_568), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g691 ( .A(n_568), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_569), .B(n_652), .Y(n_655) );
INVx3_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_570), .A2(n_691), .B(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_573), .B(n_599), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_574), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g665 ( .A(n_574), .B(n_593), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_574), .B(n_600), .Y(n_742) );
AND2x2_ASAP7_75t_L g611 ( .A(n_575), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g678 ( .A(n_575), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B(n_585), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g639 ( .A(n_578), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_578), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g663 ( .A(n_579), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_579), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_582), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_582), .A2(n_621), .B(n_651), .C(n_653), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_582), .A2(n_669), .B1(n_672), .B2(n_673), .C(n_677), .Y(n_668) );
AND2x2_ASAP7_75t_L g664 ( .A(n_583), .B(n_617), .Y(n_664) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_597), .C(n_622), .Y(n_589) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_590), .B(n_709), .C(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
OR2x2_ASAP7_75t_L g681 ( .A(n_592), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_602), .B1(n_605), .B2(n_611), .C(n_613), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_599), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g621 ( .A(n_604), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
OR2x2_ASAP7_75t_L g741 ( .A(n_604), .B(n_652), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVxp67_ASAP7_75t_L g715 ( .A(n_607), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_609), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g616 ( .A(n_610), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_612), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_612), .B(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_612), .B(n_679), .Y(n_718) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g732 ( .A(n_621), .B(n_652), .Y(n_732) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g710 ( .A(n_627), .Y(n_710) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI322xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_636), .A3(n_637), .B1(n_638), .B2(n_641), .C1(n_643), .C2(n_645), .Y(n_630) );
OAI322xp33_ASAP7_75t_L g712 ( .A1(n_631), .A2(n_713), .A3(n_714), .B1(n_715), .B2(n_716), .C1(n_717), .C2(n_719), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx4_ASAP7_75t_L g646 ( .A(n_633), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_633), .B(n_659), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_633), .B(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_636), .Y(n_731) );
INVx1_ASAP7_75t_L g709 ( .A(n_637), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g726 ( .A(n_639), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_639), .B(n_680), .Y(n_737) );
OR2x2_ASAP7_75t_L g670 ( .A(n_642), .B(n_671), .Y(n_670) );
INVxp33_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_654), .C(n_656), .Y(n_647) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_646), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g730 ( .A(n_646), .Y(n_730) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_678), .A3(n_695), .B1(n_697), .B2(n_698), .C1(n_701), .C2(n_705), .Y(n_694) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_690), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_683), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_671), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
NAND2xp33_ASAP7_75t_SL g688 ( .A(n_674), .B(n_685), .Y(n_688) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
OAI322xp33_ASAP7_75t_L g728 ( .A1(n_676), .A2(n_729), .A3(n_731), .B1(n_732), .B2(n_733), .C1(n_735), .C2(n_738), .Y(n_728) );
AOI21xp33_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_686), .B(n_734), .Y(n_743) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_694), .C(n_706), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_722), .C(n_728), .D(n_740), .Y(n_711) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_742), .B(n_743), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule