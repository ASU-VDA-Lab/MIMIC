module fake_jpeg_27194_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_51),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_58),
.B1(n_43),
.B2(n_36),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_63),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_18),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_40),
.B(n_22),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_27),
.C(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_27),
.C(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_41),
.B(n_17),
.C(n_28),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_64),
.B(n_91),
.C(n_39),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_76),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_78),
.Y(n_103)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_42),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_42),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_83),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_42),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_40),
.B(n_1),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_89),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_34),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_71),
.B(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_43),
.B1(n_36),
.B2(n_37),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_61),
.B1(n_36),
.B2(n_43),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_98),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_44),
.B1(n_28),
.B2(n_36),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_95),
.B(n_114),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_60),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_60),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.C(n_102),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_67),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_25),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_117),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_84),
.B1(n_76),
.B2(n_73),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_115),
.B1(n_37),
.B2(n_34),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_37),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_17),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_77),
.C(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_61),
.B1(n_43),
.B2(n_49),
.Y(n_128)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_23),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_16),
.CON(n_117),
.SN(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_127),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_85),
.B1(n_75),
.B2(n_92),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_71),
.B(n_87),
.C(n_64),
.D(n_83),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_16),
.B(n_20),
.Y(n_181)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_131),
.B1(n_61),
.B2(n_116),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_71),
.B1(n_87),
.B2(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_137),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_43),
.B1(n_49),
.B2(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_139),
.B1(n_47),
.B2(n_50),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_86),
.B1(n_108),
.B2(n_88),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_49),
.B1(n_90),
.B2(n_63),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_34),
.C(n_37),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_149),
.C(n_99),
.Y(n_155)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_35),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_34),
.C(n_35),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_96),
.B(n_105),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_153),
.B(n_164),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_96),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_163),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_125),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_97),
.A3(n_119),
.B1(n_102),
.B2(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_161),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_143),
.B(n_145),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_181),
.B(n_135),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_172),
.B1(n_174),
.B2(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_88),
.B1(n_116),
.B2(n_45),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_139),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_88),
.B1(n_45),
.B2(n_85),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_179),
.B1(n_123),
.B2(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_111),
.B1(n_106),
.B2(n_47),
.Y(n_177)
);

CKINVDCx12_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_123),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_132),
.B1(n_131),
.B2(n_135),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_126),
.C(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_198),
.C(n_211),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_139),
.B1(n_149),
.B2(n_126),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_201),
.B1(n_162),
.B2(n_39),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_161),
.B(n_181),
.C(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_202),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_205),
.B1(n_210),
.B2(n_32),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_207),
.B(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_136),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_200),
.B(n_180),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_135),
.B1(n_22),
.B2(n_47),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_30),
.B1(n_50),
.B2(n_23),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_39),
.C(n_35),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_39),
.B(n_25),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_150),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_216),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_175),
.B1(n_160),
.B2(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_232),
.B1(n_191),
.B2(n_210),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_164),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_171),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_166),
.C(n_153),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_156),
.C(n_167),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_172),
.C(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_188),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_39),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_209),
.C(n_189),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_27),
.C(n_19),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_39),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_24),
.B(n_26),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_201),
.B1(n_209),
.B2(n_194),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_238),
.A2(n_246),
.B1(n_233),
.B2(n_236),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_243),
.B1(n_248),
.B2(n_237),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_189),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_245),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_191),
.B1(n_205),
.B2(n_193),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_212),
.B1(n_199),
.B2(n_185),
.Y(n_246)
);

AND3x1_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_212),
.C(n_185),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_255),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_230),
.C(n_235),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_26),
.C(n_25),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_252),
.C(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_24),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_216),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_225),
.B(n_223),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_250),
.B(n_241),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_262),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_229),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_271),
.C(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_214),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_242),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_220),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_274),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_236),
.C(n_26),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_247),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_24),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_8),
.C(n_14),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_249),
.B(n_241),
.C(n_246),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_9),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.C(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_283),
.C(n_270),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_257),
.C(n_253),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_248),
.B(n_8),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_9),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_15),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_276),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_300),
.C(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_273),
.B1(n_1),
.B2(n_2),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_297),
.B1(n_1),
.B2(n_2),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_286),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_15),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_11),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_280),
.C(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_307),
.C(n_7),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_309),
.B(n_3),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_279),
.A3(n_281),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_5),
.B(n_6),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_292),
.B(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_300),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_5),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_303),
.B(n_302),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_318),
.B1(n_320),
.B2(n_317),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_6),
.B(n_7),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_7),
.Y(n_324)
);


endmodule