module fake_aes_642_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
NOR2xp33_ASAP7_75t_R g3 ( .A(n_2), .B(n_0), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
AOI22xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
CKINVDCx9p33_ASAP7_75t_R g7 ( .A(n_4), .Y(n_7) );
OA21x2_ASAP7_75t_L g8 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_8) );
BUFx3_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_9), .Y(n_11) );
OR2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_6), .Y(n_12) );
NOR4xp25_ASAP7_75t_L g13 ( .A(n_12), .B(n_7), .C(n_2), .D(n_1), .Y(n_13) );
AOI211xp5_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_7), .B(n_9), .C(n_11), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_14), .B(n_9), .Y(n_15) );
NOR3xp33_ASAP7_75t_SL g16 ( .A(n_13), .B(n_0), .C(n_1), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
OAI222xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_0), .B1(n_16), .B2(n_15), .C1(n_6), .C2(n_13), .Y(n_18) );
endmodule