module fake_netlist_1_8506_n_677 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_677);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_677;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g77 ( .A(n_73), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_32), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_44), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_49), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_41), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_1), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_38), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_7), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_57), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_5), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_39), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_48), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_33), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_35), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_53), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_64), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_16), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_36), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_43), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_68), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_51), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_61), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_14), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_23), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_67), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_46), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_86), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_90), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_90), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_106), .B(n_0), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_108), .B(n_1), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_84), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_96), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_117), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_100), .Y(n_140) );
NOR2xp33_ASAP7_75t_R g141 ( .A(n_104), .B(n_31), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_102), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_98), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_98), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_82), .B(n_4), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_91), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_114), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_82), .B(n_6), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_85), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_83), .B(n_9), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_79), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_79), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
NOR3xp33_ASAP7_75t_L g164 ( .A(n_83), .B(n_9), .C(n_10), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_99), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_80), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_80), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_87), .B(n_10), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_156), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_135), .A2(n_115), .B1(n_94), .B2(n_103), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_166), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
NAND3xp33_ASAP7_75t_L g174 ( .A(n_134), .B(n_94), .C(n_103), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_144), .B(n_125), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_139), .A2(n_112), .B1(n_87), .B2(n_88), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_144), .B(n_112), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_167), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_144), .B(n_113), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_130), .B(n_111), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_145), .B(n_119), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_151), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_169), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_131), .B(n_111), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_137), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_135), .B(n_115), .Y(n_197) );
OR2x2_ASAP7_75t_SL g198 ( .A(n_145), .B(n_119), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_135), .B(n_88), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_129), .B(n_105), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_132), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
INVxp67_ASAP7_75t_SL g205 ( .A(n_137), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_133), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_169), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_160), .A2(n_105), .B1(n_120), .B2(n_118), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
NAND3x1_ASAP7_75t_L g212 ( .A(n_164), .B(n_120), .C(n_118), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_160), .B(n_124), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_146), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_162), .B(n_97), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_146), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_156), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_162), .B(n_124), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_129), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_161), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_161), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g229 ( .A1(n_139), .A2(n_97), .B1(n_122), .B2(n_109), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_142), .B(n_122), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_142), .B(n_123), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_147), .B(n_123), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_126), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_160), .B(n_97), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_195), .Y(n_235) );
OR2x2_ASAP7_75t_SL g236 ( .A(n_175), .B(n_136), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_234), .Y(n_237) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_187), .B(n_164), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_234), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_213), .B(n_158), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_176), .B(n_158), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_213), .B(n_147), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_187), .B(n_168), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_199), .B(n_154), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_180), .B(n_153), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_180), .B(n_168), .Y(n_252) );
NOR2x1_ASAP7_75t_L g253 ( .A(n_174), .B(n_168), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
AND3x2_ASAP7_75t_SL g256 ( .A(n_170), .B(n_140), .C(n_143), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_195), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_193), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_182), .B(n_165), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_177), .B(n_138), .C(n_134), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_219), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
NAND2xp33_ASAP7_75t_SL g264 ( .A(n_226), .B(n_141), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_201), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_199), .B(n_148), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_193), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_197), .B(n_165), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_197), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_195), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_201), .B(n_163), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_171), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_198), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_201), .B(n_163), .Y(n_274) );
OR2x6_ASAP7_75t_L g275 ( .A(n_229), .B(n_148), .Y(n_275) );
AND2x4_ASAP7_75t_SL g276 ( .A(n_171), .B(n_159), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_177), .B(n_157), .C(n_77), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_198), .A2(n_157), .B1(n_159), .B2(n_155), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_230), .B(n_155), .Y(n_280) );
NAND2xp33_ASAP7_75t_SL g281 ( .A(n_226), .B(n_141), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_230), .B(n_153), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_172), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_181), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_217), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_230), .B(n_152), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_230), .Y(n_289) );
OAI22xp5_ASAP7_75t_SL g290 ( .A1(n_209), .A2(n_185), .B1(n_192), .B2(n_212), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_196), .B(n_152), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_223), .B(n_150), .Y(n_292) );
BUFx8_ASAP7_75t_L g293 ( .A(n_178), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_196), .B(n_150), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_212), .B(n_97), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_178), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_196), .B(n_116), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_205), .B(n_109), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_231), .B(n_78), .Y(n_299) );
XNOR2xp5_ASAP7_75t_SL g300 ( .A(n_179), .B(n_11), .Y(n_300) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_214), .B(n_121), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_179), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_204), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_291), .A2(n_196), .B(n_224), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_239), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_239), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_280), .A2(n_227), .B(n_204), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_235), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_237), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_302), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_241), .B(n_204), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_242), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_247), .B(n_232), .Y(n_314) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_276), .B(n_224), .Y(n_315) );
AND2x6_ASAP7_75t_L g316 ( .A(n_251), .B(n_204), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_302), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
BUFx10_ASAP7_75t_L g319 ( .A(n_276), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_268), .B(n_181), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
O2A1O1Ixp5_ASAP7_75t_L g323 ( .A1(n_264), .A2(n_224), .B(n_225), .C(n_214), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_258), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_296), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_269), .B(n_224), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_246), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_265), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_294), .A2(n_215), .B(n_216), .Y(n_329) );
CKINVDCx14_ASAP7_75t_R g330 ( .A(n_263), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_283), .A2(n_215), .B(n_216), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_272), .A2(n_189), .B1(n_186), .B2(n_181), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_247), .B(n_186), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_289), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_258), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_246), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_237), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_266), .B(n_189), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_288), .A2(n_218), .B(n_225), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_271), .A2(n_218), .B(n_225), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_255), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_270), .B(n_181), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_270), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_274), .A2(n_225), .B(n_227), .Y(n_346) );
INVx3_ASAP7_75t_SL g347 ( .A(n_287), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_268), .B(n_107), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_293), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_247), .A2(n_101), .B1(n_121), .B2(n_200), .C(n_206), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_240), .B(n_11), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_238), .A2(n_200), .B1(n_191), .B2(n_206), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_245), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_259), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_259), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_307), .A2(n_279), .B(n_253), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_351), .B(n_295), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_307), .A2(n_228), .B(n_220), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_315), .A2(n_287), .B1(n_298), .B2(n_254), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_304), .A2(n_297), .B(n_281), .Y(n_362) );
CKINVDCx12_ASAP7_75t_R g363 ( .A(n_349), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_306), .B(n_238), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_262), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_305), .A2(n_273), .B1(n_248), .B2(n_295), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_323), .A2(n_228), .B(n_211), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_330), .A2(n_300), .B1(n_290), .B2(n_244), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_349), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_314), .A2(n_261), .B1(n_244), .B2(n_278), .C(n_250), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_322), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_275), .B1(n_295), .B2(n_278), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_342), .B(n_346), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_315), .A2(n_298), .B1(n_254), .B2(n_299), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_351), .A2(n_275), .B1(n_252), .B2(n_299), .Y(n_378) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_322), .A2(n_149), .A3(n_127), .B(n_128), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_354), .B(n_252), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_308), .B(n_303), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_354), .B(n_275), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_325), .A2(n_228), .B(n_220), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_310), .Y(n_385) );
NAND3xp33_ASAP7_75t_SL g386 ( .A(n_332), .B(n_261), .C(n_243), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_348), .A2(n_260), .B1(n_292), .B2(n_298), .C(n_264), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_308), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_347), .A2(n_256), .B1(n_260), .B2(n_236), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_370), .A2(n_332), .B1(n_319), .B2(n_333), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_372), .A2(n_387), .B(n_362), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_361), .A2(n_319), .B1(n_309), .B2(n_339), .Y(n_392) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_360), .B(n_380), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_386), .A2(n_319), .B1(n_309), .B2(n_339), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_360), .B(n_340), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_358), .A2(n_317), .B1(n_311), .B2(n_350), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_389), .A2(n_314), .B(n_334), .C(n_348), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_382), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_358), .A2(n_317), .B1(n_311), .B2(n_336), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_360), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_375), .A2(n_321), .B1(n_281), .B2(n_336), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_375), .A2(n_321), .B1(n_335), .B2(n_326), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_383), .A2(n_321), .B1(n_335), .B2(n_334), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_378), .A2(n_352), .B1(n_313), .B2(n_328), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_365), .B(n_312), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_357), .B(n_301), .C(n_221), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_365), .B(n_312), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_367), .A2(n_256), .B1(n_328), .B2(n_345), .C(n_331), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_358), .A2(n_313), .B1(n_308), .B2(n_310), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_363), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_358), .A2(n_313), .B1(n_308), .B2(n_310), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_310), .B1(n_324), .B2(n_320), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_383), .B(n_312), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_364), .A2(n_345), .B1(n_316), .B2(n_337), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_366), .B(n_286), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_398), .A2(n_381), .B(n_369), .C(n_373), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_396), .B(n_366), .Y(n_422) );
NOR2x1_ASAP7_75t_SL g423 ( .A(n_399), .B(n_374), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_374), .B1(n_371), .B2(n_357), .C1(n_301), .C2(n_363), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_396), .B(n_388), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_393), .A2(n_359), .B(n_376), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_286), .B1(n_329), .B2(n_388), .C(n_373), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_406), .A2(n_373), .B1(n_388), .B2(n_316), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_400), .A2(n_373), .B1(n_388), .B2(n_382), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_417), .B(n_385), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_344), .B1(n_385), .B2(n_337), .C(n_320), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_382), .B1(n_385), .B2(n_353), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g433 ( .A1(n_394), .A2(n_385), .B1(n_316), .B2(n_310), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_405), .A2(n_126), .A3(n_149), .B1(n_128), .B2(n_127), .B3(n_220), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_385), .B1(n_337), .B2(n_320), .C(n_149), .Y(n_435) );
AOI31xp33_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_327), .A3(n_338), .B(n_343), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_417), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_359), .B(n_376), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_408), .A2(n_126), .B1(n_128), .B2(n_127), .C(n_324), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_316), .B1(n_327), .B2(n_338), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_399), .B(n_379), .Y(n_442) );
OAI33xp33_ASAP7_75t_L g443 ( .A1(n_414), .A2(n_211), .A3(n_210), .B1(n_191), .B2(n_208), .B3(n_233), .Y(n_443) );
NAND2xp33_ASAP7_75t_R g444 ( .A(n_394), .B(n_12), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_411), .B(n_353), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_412), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_418), .B(n_379), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_393), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_418), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_415), .B(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
NOR5xp2_ASAP7_75t_SL g454 ( .A(n_397), .B(n_13), .C(n_15), .D(n_16), .E(n_17), .Y(n_454) );
OAI221xp5_ASAP7_75t_SL g455 ( .A1(n_424), .A2(n_397), .B1(n_392), .B2(n_395), .C(n_416), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_449), .Y(n_456) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_426), .A2(n_368), .B(n_384), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_451), .A2(n_316), .B1(n_353), .B2(n_355), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_449), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_439), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_448), .B(n_439), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_448), .B(n_379), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_437), .B(n_379), .Y(n_464) );
OAI33xp33_ASAP7_75t_L g465 ( .A1(n_437), .A2(n_13), .A3(n_15), .B1(n_17), .B2(n_18), .B3(n_19), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_447), .B(n_379), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_451), .A2(n_316), .B1(n_353), .B2(n_356), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_422), .B(n_420), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_450), .B(n_379), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_447), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_368), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_384), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_442), .B(n_211), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_421), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_422), .A2(n_324), .B1(n_356), .B2(n_343), .C(n_355), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_450), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_442), .B(n_18), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_431), .A2(n_353), .B1(n_324), .B2(n_303), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_452), .B(n_19), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_452), .B(n_20), .Y(n_482) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_453), .B(n_324), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_21), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_419), .A2(n_227), .B(n_233), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_438), .B(n_22), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_425), .B(n_22), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_444), .B(n_23), .C(n_24), .D(n_227), .Y(n_489) );
OAI211xp5_ASAP7_75t_SL g490 ( .A1(n_446), .A2(n_208), .B(n_210), .C(n_233), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_453), .B(n_24), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_423), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_432), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_429), .B(n_222), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_445), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_428), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_433), .B(n_222), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_443), .B(n_26), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_434), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_435), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_454), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_427), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_441), .A2(n_267), .B1(n_222), .B2(n_221), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_454), .B(n_222), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_462), .B(n_222), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_487), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_462), .B(n_222), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_470), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_487), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_470), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_463), .B(n_28), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_489), .B(n_40), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_463), .B(n_42), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
NAND2xp33_ASAP7_75t_R g519 ( .A(n_479), .B(n_45), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_492), .B(n_267), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_489), .B(n_47), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_492), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_496), .A2(n_285), .B1(n_282), .B2(n_257), .Y(n_523) );
NAND2xp33_ASAP7_75t_SL g524 ( .A(n_479), .B(n_50), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_463), .B(n_52), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_478), .B(n_54), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_477), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_468), .B(n_55), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_478), .B(n_58), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_479), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_477), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_471), .B(n_59), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g535 ( .A1(n_502), .A2(n_203), .B1(n_202), .B2(n_194), .C(n_190), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_481), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_464), .B(n_60), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_456), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_456), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_475), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_464), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_484), .B(n_65), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_471), .B(n_66), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_466), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_471), .B(n_69), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_466), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_481), .Y(n_547) );
NAND4xp25_ASAP7_75t_SL g548 ( .A(n_481), .B(n_71), .C(n_72), .D(n_75), .Y(n_548) );
NOR4xp25_ASAP7_75t_SL g549 ( .A(n_455), .B(n_76), .C(n_183), .D(n_285), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_474), .Y(n_550) );
NAND2xp33_ASAP7_75t_R g551 ( .A(n_482), .B(n_173), .Y(n_551) );
NAND2xp33_ASAP7_75t_SL g552 ( .A(n_482), .B(n_285), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_484), .B(n_173), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_465), .A2(n_173), .B1(n_203), .B2(n_184), .C(n_190), .Y(n_554) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_483), .B(n_285), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_484), .B(n_202), .Y(n_556) );
NAND2xp33_ASAP7_75t_SL g557 ( .A(n_482), .B(n_282), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_502), .B(n_257), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_459), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_466), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_486), .B(n_202), .Y(n_561) );
INVx4_ASAP7_75t_L g562 ( .A(n_483), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_516), .B(n_502), .C(n_486), .Y(n_563) );
AOI21xp33_ASAP7_75t_L g564 ( .A1(n_519), .A2(n_491), .B(n_505), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_532), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_546), .B(n_473), .Y(n_566) );
OAI221xp5_ASAP7_75t_SL g567 ( .A1(n_542), .A2(n_496), .B1(n_488), .B2(n_497), .C(n_503), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_521), .B(n_505), .C(n_497), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_544), .B(n_503), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_560), .B(n_473), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_540), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_538), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_541), .B(n_491), .Y(n_573) );
AOI322xp5_ASAP7_75t_L g574 ( .A1(n_547), .A2(n_530), .A3(n_524), .B1(n_536), .B2(n_552), .C1(n_557), .C2(n_515), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_547), .A2(n_483), .B1(n_495), .B2(n_488), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_558), .A2(n_504), .B(n_490), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_538), .A2(n_465), .B1(n_455), .B2(n_501), .C(n_493), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_551), .A2(n_490), .B1(n_501), .B2(n_499), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_527), .B(n_531), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_542), .A2(n_467), .B1(n_458), .B2(n_480), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_522), .A2(n_495), .B1(n_469), .B2(n_476), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_515), .B(n_474), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_522), .A2(n_493), .B(n_469), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_548), .A2(n_506), .B1(n_500), .B2(n_476), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_508), .B(n_474), .Y(n_588) );
OAI32xp33_ASAP7_75t_L g589 ( .A1(n_517), .A2(n_494), .A3(n_498), .B1(n_504), .B2(n_500), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_513), .Y(n_590) );
AND3x2_ASAP7_75t_L g591 ( .A(n_513), .B(n_498), .C(n_473), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_550), .B(n_474), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_517), .A2(n_498), .B(n_494), .C(n_506), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g594 ( .A(n_520), .B(n_457), .Y(n_594) );
OR3x1_ASAP7_75t_L g595 ( .A(n_512), .B(n_485), .C(n_472), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_550), .B(n_460), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_500), .B1(n_485), .B2(n_460), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_507), .B(n_472), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_534), .A2(n_460), .B1(n_472), .B2(n_457), .Y(n_600) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_562), .A2(n_457), .B(n_184), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_534), .B(n_457), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_525), .A2(n_457), .B1(n_282), .B2(n_257), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
NAND2xp33_ASAP7_75t_R g606 ( .A(n_591), .B(n_549), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_590), .B(n_562), .Y(n_607) );
XNOR2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_520), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_573), .B(n_539), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_569), .B(n_539), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
AOI22xp5_ASAP7_75t_SL g612 ( .A1(n_583), .A2(n_588), .B1(n_562), .B2(n_582), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_574), .B(n_555), .Y(n_613) );
XNOR2x2_ASAP7_75t_L g614 ( .A(n_568), .B(n_526), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_588), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_575), .A2(n_564), .B1(n_593), .B2(n_577), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_566), .Y(n_617) );
NAND2xp33_ASAP7_75t_L g618 ( .A(n_584), .B(n_526), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
NOR3xp33_ASAP7_75t_SL g620 ( .A(n_567), .B(n_528), .C(n_535), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_601), .B(n_555), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_570), .B(n_572), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_575), .B(n_549), .C(n_537), .Y(n_623) );
NOR3x1_ASAP7_75t_L g624 ( .A(n_598), .B(n_537), .C(n_556), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_605), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_603), .B(n_555), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_579), .A2(n_562), .B1(n_545), .B2(n_543), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_578), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_581), .B(n_556), .Y(n_630) );
AOI221x1_ASAP7_75t_SL g631 ( .A1(n_599), .A2(n_518), .B1(n_511), .B2(n_510), .C(n_559), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_615), .B(n_602), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_616), .A2(n_595), .B1(n_587), .B2(n_592), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_613), .A2(n_576), .B1(n_594), .B2(n_600), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_617), .B(n_596), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_613), .A2(n_587), .B1(n_603), .B2(n_594), .C(n_597), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_609), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_607), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_622), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_612), .B(n_591), .C(n_553), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_631), .A2(n_589), .B1(n_553), .B2(n_561), .C(n_586), .Y(n_641) );
OAI22xp5_ASAP7_75t_SL g642 ( .A1(n_630), .A2(n_523), .B1(n_518), .B2(n_511), .Y(n_642) );
INVx8_ASAP7_75t_L g643 ( .A(n_608), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_626), .B(n_604), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_623), .B(n_529), .C(n_509), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_630), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_621), .A2(n_529), .B(n_597), .Y(n_647) );
AOI322xp5_ASAP7_75t_L g648 ( .A1(n_618), .A2(n_604), .A3(n_565), .B1(n_585), .B2(n_586), .C1(n_510), .C2(n_554), .Y(n_648) );
NAND3x1_ASAP7_75t_SL g649 ( .A(n_614), .B(n_585), .C(n_183), .Y(n_649) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_634), .B(n_621), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_640), .B(n_611), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_633), .A2(n_628), .B1(n_627), .B2(n_620), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_636), .B(n_627), .Y(n_653) );
INVxp33_ASAP7_75t_L g654 ( .A(n_645), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_643), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_643), .A2(n_618), .B(n_610), .Y(n_656) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_643), .B(n_625), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_637), .A2(n_629), .B1(n_619), .B2(n_624), .C(n_606), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_644), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_647), .A2(n_606), .B1(n_619), .B2(n_190), .C(n_194), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g661 ( .A(n_648), .B(n_183), .C(n_249), .D(n_282), .E(n_641), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_638), .A2(n_183), .B1(n_249), .B2(n_642), .C(n_632), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_639), .A2(n_249), .B1(n_635), .B2(n_649), .Y(n_663) );
AOI221xp5_ASAP7_75t_SL g664 ( .A1(n_634), .A2(n_646), .B1(n_636), .B2(n_613), .C(n_637), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_655), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_650), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_659), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_652), .A2(n_654), .B(n_663), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_665), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_666), .B(n_664), .Y(n_670) );
AND3x1_ASAP7_75t_L g671 ( .A(n_667), .B(n_653), .C(n_657), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_669), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_670), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_672), .A2(n_665), .B1(n_671), .B2(n_668), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
AOI22xp5_ASAP7_75t_SL g676 ( .A1(n_674), .A2(n_661), .B1(n_656), .B2(n_651), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_675), .B1(n_658), .B2(n_662), .C(n_660), .Y(n_677) );
endmodule