module fake_ariane_209_n_1731 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1731);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1731;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g157 ( 
.A(n_10),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_48),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_32),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_48),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_77),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_51),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_40),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_39),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_97),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_32),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_46),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_20),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_55),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_1),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_15),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_72),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_50),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_37),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_78),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_53),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_87),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_56),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_46),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_74),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_136),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_130),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_17),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_29),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_58),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_57),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_49),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_95),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_24),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_16),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_143),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_79),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_47),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_36),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_85),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_102),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_73),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_20),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_76),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_88),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_13),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_119),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_121),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_26),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_132),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_135),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_55),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_62),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_104),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_122),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_139),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_148),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_28),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_19),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_53),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_12),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_45),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_67),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_51),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_43),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_134),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_21),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_115),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_150),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_112),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_127),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_126),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_75),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_111),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_40),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_30),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_68),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_128),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_19),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_21),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_84),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_129),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_42),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_52),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_2),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_144),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_56),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_54),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_146),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_35),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_63),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_96),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_110),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_162),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_3),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_174),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_162),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_203),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_163),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_200),
.B(n_213),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_180),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_191),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_199),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_203),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_184),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_223),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_226),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_184),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_179),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_231),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_158),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_165),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_206),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_232),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_217),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_160),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_161),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_262),
.Y(n_345)
);

NAND2xp33_ASAP7_75t_R g346 ( 
.A(n_200),
.B(n_59),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_166),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_167),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_272),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_195),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_169),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_196),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_263),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_176),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_171),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_196),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_204),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_213),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_173),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_203),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_178),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_193),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_293),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_203),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_293),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_R g368 ( 
.A(n_168),
.B(n_106),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_245),
.B(n_3),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_202),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_204),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_4),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_218),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_304),
.B(n_7),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_211),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_293),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_221),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_212),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_224),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_293),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_215),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_216),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_216),
.B(n_228),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_228),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_179),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_241),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_236),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_227),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_322),
.A2(n_243),
.B(n_241),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_346),
.B(n_314),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_326),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_210),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_335),
.B(n_194),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_386),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_308),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_243),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_337),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_340),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_248),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_341),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_321),
.B(n_248),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_258),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g422 ( 
.A1(n_331),
.A2(n_249),
.B(n_258),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_343),
.B(n_170),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_327),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_344),
.B(n_313),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_338),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_335),
.B(n_194),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_329),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_332),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_336),
.Y(n_435)
);

BUFx8_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_360),
.A2(n_276),
.B1(n_157),
.B2(n_251),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_271),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_359),
.B(n_271),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_359),
.B(n_285),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_339),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_348),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_349),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_342),
.B(n_172),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_354),
.A2(n_175),
.B1(n_182),
.B2(n_309),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_376),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_352),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_345),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_356),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_407),
.A2(n_369),
.B1(n_358),
.B2(n_375),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_395),
.B(n_317),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_403),
.B(n_317),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_411),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_442),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_412),
.B(n_400),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_397),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_401),
.B(n_318),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_285),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_398),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_415),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_418),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_433),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_403),
.B(n_384),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_408),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_418),
.Y(n_493)
);

NOR2x1p5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_361),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_433),
.B(n_363),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_399),
.B(n_364),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_286),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_429),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_405),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

INVx6_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_370),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_427),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_433),
.B(n_373),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_457),
.B(n_388),
.C(n_381),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_402),
.B(n_384),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_453),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_453),
.B(n_286),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_405),
.A2(n_385),
.B1(n_387),
.B2(n_390),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_442),
.B(n_385),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_434),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_453),
.B(n_291),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_466),
.B(n_291),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_461),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_404),
.A2(n_460),
.B1(n_372),
.B2(n_375),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_448),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_401),
.B(n_318),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_442),
.B(n_387),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_461),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_421),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_430),
.B(n_316),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_423),
.B(n_389),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_461),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_462),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_462),
.B(n_297),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_462),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_462),
.B(n_297),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_438),
.B(n_390),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_462),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_430),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_458),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_416),
.B(n_392),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_443),
.B(n_319),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_443),
.B(n_391),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_430),
.B(n_372),
.Y(n_554)
);

INVx6_ASAP7_75t_L g555 ( 
.A(n_430),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_455),
.B(n_176),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_394),
.A2(n_383),
.B1(n_377),
.B2(n_365),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_394),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_447),
.B(n_333),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_464),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_463),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_465),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_465),
.B(n_367),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_394),
.A2(n_265),
.B1(n_311),
.B2(n_310),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_426),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_259),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_432),
.B(n_305),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_424),
.B(n_368),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_432),
.B(n_305),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_413),
.B(n_159),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_454),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_439),
.B(n_159),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_428),
.B(n_177),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_455),
.B(n_454),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_413),
.B(n_229),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_417),
.A2(n_270),
.B1(n_233),
.B2(n_234),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_459),
.B(n_177),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_444),
.B(n_183),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_409),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_444),
.B(n_186),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_450),
.B(n_188),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_450),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_394),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_451),
.B(n_188),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_451),
.B(n_219),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_417),
.B(n_254),
.Y(n_596)
);

NOR2x1p5_ASAP7_75t_L g597 ( 
.A(n_436),
.B(n_181),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_451),
.B(n_189),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_419),
.B(n_445),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_456),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_456),
.B(n_192),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_419),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_456),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_459),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_409),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_459),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_445),
.B(n_197),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_446),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_446),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_396),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_409),
.B(n_256),
.Y(n_611)
);

AND2x4_ASAP7_75t_SL g612 ( 
.A(n_436),
.B(n_350),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_396),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_422),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_480),
.B(n_437),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_559),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_599),
.B(n_436),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_608),
.B(n_436),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_469),
.B(n_499),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_260),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_491),
.B(n_422),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_264),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_556),
.A2(n_488),
.B1(n_481),
.B2(n_484),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_547),
.B(n_210),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_533),
.B(n_210),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_545),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_602),
.B(n_265),
.Y(n_629)
);

BUFx5_ASAP7_75t_L g630 ( 
.A(n_497),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_492),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_478),
.B(n_437),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_565),
.B(n_409),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_496),
.B(n_266),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_565),
.B(n_219),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_571),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_210),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_181),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_596),
.B(n_185),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_498),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_483),
.B(n_185),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_483),
.B(n_187),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_483),
.B(n_187),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_524),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_579),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_502),
.B(n_268),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_473),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_565),
.B(n_238),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_476),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_547),
.B(n_269),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_190),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_483),
.B(n_491),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_483),
.B(n_190),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_574),
.B(n_497),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_547),
.B(n_238),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_SL g660 ( 
.A(n_494),
.B(n_273),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_481),
.A2(n_220),
.B1(n_235),
.B2(n_311),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_586),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_506),
.B(n_274),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_568),
.B(n_275),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_501),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_475),
.B(n_205),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_467),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_576),
.B(n_205),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_516),
.A2(n_279),
.B(n_214),
.C(n_220),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_607),
.B(n_207),
.Y(n_674)
);

OAI22x1_ASAP7_75t_L g675 ( 
.A1(n_582),
.A2(n_298),
.B1(n_294),
.B2(n_299),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_485),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_524),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_551),
.B(n_207),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_471),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_484),
.B(n_503),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_560),
.B(n_302),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_532),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_503),
.B(n_267),
.C(n_214),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_531),
.B(n_235),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_486),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_493),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_487),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_531),
.B(n_505),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_509),
.B(n_240),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_471),
.B(n_306),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_523),
.B(n_240),
.Y(n_692)
);

AOI21x1_ASAP7_75t_L g693 ( 
.A1(n_585),
.A2(n_414),
.B(n_410),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_476),
.B(n_255),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_537),
.B(n_242),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_476),
.B(n_255),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_606),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_548),
.B(n_242),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_570),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_549),
.A2(n_307),
.B1(n_279),
.B2(n_247),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_550),
.B(n_247),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_581),
.A2(n_278),
.B1(n_201),
.B2(n_208),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_476),
.B(n_277),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_557),
.B(n_267),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_508),
.B(n_517),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_577),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_612),
.A2(n_521),
.B1(n_515),
.B2(n_517),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_500),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_591),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_501),
.B(n_295),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_555),
.B(n_300),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_581),
.B(n_198),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_559),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_567),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_572),
.B(n_300),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_592),
.Y(n_716)
);

AOI22x1_ASAP7_75t_SL g717 ( 
.A1(n_544),
.A2(n_307),
.B1(n_303),
.B2(n_310),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_510),
.B(n_303),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_612),
.B(n_203),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_487),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_482),
.A2(n_209),
.B1(n_222),
.B2(n_230),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_600),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_529),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_515),
.B(n_237),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_482),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_468),
.B(n_239),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_515),
.B(n_244),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_487),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_497),
.B(n_257),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_535),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_535),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_603),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_527),
.A2(n_249),
.B(n_277),
.C(n_292),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_500),
.B(n_292),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_541),
.B(n_246),
.Y(n_736)
);

AO22x1_ASAP7_75t_L g737 ( 
.A1(n_497),
.A2(n_236),
.B1(n_261),
.B2(n_282),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_555),
.B(n_250),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_555),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_611),
.B(n_252),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_578),
.B(n_261),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_497),
.B(n_253),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_604),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_472),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_558),
.B(n_257),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_500),
.B(n_249),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_497),
.B(n_257),
.Y(n_747)
);

INVxp67_ASAP7_75t_SL g748 ( 
.A(n_593),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_468),
.B(n_296),
.Y(n_749)
);

BUFx8_ASAP7_75t_L g750 ( 
.A(n_519),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_614),
.A2(n_593),
.B(n_513),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_SL g752 ( 
.A(n_584),
.B(n_280),
.C(n_281),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_495),
.B(n_8),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_500),
.B(n_249),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_519),
.A2(n_257),
.B1(n_283),
.B2(n_425),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_597),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_495),
.B(n_312),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_504),
.B(n_9),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_482),
.A2(n_287),
.B1(n_284),
.B2(n_257),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_504),
.A2(n_573),
.B(n_575),
.C(n_587),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_569),
.A2(n_257),
.B1(n_283),
.B2(n_425),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_535),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_482),
.B(n_525),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_512),
.B(n_283),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_525),
.A2(n_425),
.B1(n_283),
.B2(n_410),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_525),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_525),
.B(n_425),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_554),
.B(n_414),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_554),
.B(n_10),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_554),
.B(n_588),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_554),
.B(n_414),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_588),
.B(n_410),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_511),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_588),
.B(n_406),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_512),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_589),
.A2(n_598),
.B1(n_601),
.B2(n_540),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_618),
.B(n_605),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_774),
.A2(n_605),
.B(n_563),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_772),
.A2(n_751),
.B(n_760),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_634),
.B(n_514),
.C(n_540),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_620),
.B(n_605),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_628),
.B(n_474),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_620),
.B(n_625),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_617),
.A2(n_563),
.B(n_477),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_669),
.B(n_679),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_637),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_634),
.B(n_477),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_639),
.A2(n_580),
.B(n_514),
.C(n_536),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_649),
.B(n_477),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_713),
.A2(n_563),
.B(n_546),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_748),
.A2(n_522),
.B(n_539),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_616),
.A2(n_595),
.B1(n_594),
.B2(n_590),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_724),
.A2(n_546),
.B(n_526),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_753),
.A2(n_534),
.B(n_539),
.C(n_561),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_653),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_776),
.A2(n_534),
.B(n_507),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_623),
.A2(n_513),
.B(n_522),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_753),
.A2(n_507),
.B(n_564),
.C(n_526),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_650),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_613),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_627),
.B(n_511),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_633),
.A2(n_561),
.B(n_564),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_622),
.B(n_489),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_638),
.B(n_538),
.Y(n_804)
);

NAND2x1_ASAP7_75t_L g805 ( 
.A(n_653),
.B(n_512),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_633),
.A2(n_610),
.B(n_538),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_623),
.A2(n_595),
.B(n_594),
.Y(n_807)
);

OAI21xp33_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_536),
.B(n_518),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_624),
.B(n_490),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_624),
.B(n_490),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_689),
.A2(n_562),
.B1(n_552),
.B2(n_520),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_658),
.A2(n_610),
.B(n_562),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_681),
.B(n_528),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_740),
.A2(n_652),
.B(n_635),
.Y(n_814)
);

O2A1O1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_672),
.A2(n_518),
.B(n_590),
.C(n_585),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_635),
.A2(n_542),
.B(n_530),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_652),
.A2(n_542),
.B(n_530),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_654),
.B(n_542),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_758),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_654),
.B(n_542),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_667),
.A2(n_528),
.B1(n_520),
.B2(n_512),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_766),
.B(n_528),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_659),
.A2(n_770),
.B(n_744),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_670),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_676),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_744),
.A2(n_520),
.B(n_406),
.Y(n_826)
);

NOR2x1_ASAP7_75t_L g827 ( 
.A(n_669),
.B(n_406),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_615),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_659),
.A2(n_406),
.B(n_81),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_705),
.B(n_406),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_667),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_831)
);

OAI321xp33_ASAP7_75t_L g832 ( 
.A1(n_671),
.A2(n_31),
.A3(n_34),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_688),
.A2(n_99),
.B(n_153),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_710),
.B(n_711),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_769),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_44),
.C(n_45),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_688),
.A2(n_105),
.B(n_152),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_711),
.B(n_47),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_721),
.A2(n_109),
.B(n_149),
.Y(n_839)
);

INVx11_ASAP7_75t_L g840 ( 
.A(n_750),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_686),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_721),
.A2(n_731),
.B(n_729),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_729),
.A2(n_98),
.B(n_147),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_731),
.A2(n_93),
.B(n_145),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_769),
.A2(n_50),
.B(n_54),
.C(n_61),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_656),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_621),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_687),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_680),
.B(n_83),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_732),
.A2(n_117),
.B(n_120),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_679),
.B(n_124),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_631),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_732),
.A2(n_155),
.B(n_762),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_694),
.A2(n_735),
.B(n_703),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_714),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_743),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_668),
.A2(n_736),
.B1(n_674),
.B2(n_762),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_SL g859 ( 
.A(n_684),
.B(n_682),
.C(n_722),
.Y(n_859)
);

O2A1O1Ixp5_ASAP7_75t_L g860 ( 
.A1(n_734),
.A2(n_746),
.B(n_754),
.C(n_757),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_629),
.B(n_691),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_630),
.B(n_683),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_699),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_773),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_706),
.A2(n_709),
.B(n_733),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_691),
.B(n_685),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_745),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_630),
.B(n_750),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_678),
.B(n_763),
.Y(n_869)
);

OAI321xp33_ASAP7_75t_L g870 ( 
.A1(n_632),
.A2(n_755),
.A3(n_752),
.B1(n_700),
.B2(n_728),
.C(n_725),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_642),
.B(n_756),
.Y(n_871)
);

AOI22x1_ASAP7_75t_L g872 ( 
.A1(n_706),
.A2(n_716),
.B1(n_733),
.B2(n_723),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_630),
.B(n_707),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_716),
.A2(n_723),
.B(n_651),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_626),
.B(n_663),
.C(n_660),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_718),
.B(n_739),
.Y(n_876)
);

AO22x1_ASAP7_75t_L g877 ( 
.A1(n_720),
.A2(n_719),
.B1(n_677),
.B2(n_632),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_643),
.A2(n_655),
.B(n_645),
.C(n_646),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_657),
.B(n_698),
.Y(n_879)
);

INVx5_ASAP7_75t_L g880 ( 
.A(n_641),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_759),
.A2(n_726),
.B1(n_632),
.B2(n_630),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_647),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_690),
.B(n_692),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_653),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_730),
.A2(n_747),
.B(n_673),
.C(n_636),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_636),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_630),
.B(n_738),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_726),
.A2(n_630),
.B1(n_749),
.B2(n_727),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_695),
.B(n_701),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_704),
.B(n_726),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_644),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_767),
.A2(n_675),
.B1(n_702),
.B2(n_712),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_641),
.B(n_648),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_746),
.A2(n_754),
.B(n_648),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_662),
.A2(n_697),
.B(n_665),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_653),
.B(n_708),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_662),
.A2(n_664),
.B(n_742),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_664),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_768),
.B(n_771),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_641),
.B(n_761),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_737),
.B(n_775),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_696),
.A2(n_735),
.B(n_703),
.Y(n_902)
);

OR2x6_ASAP7_75t_SL g903 ( 
.A(n_677),
.B(n_765),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_708),
.A2(n_775),
.B1(n_696),
.B2(n_764),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_708),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_741),
.A2(n_649),
.B1(n_634),
.B2(n_618),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_775),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_717),
.A2(n_760),
.B(n_724),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_634),
.A2(n_649),
.B(n_620),
.C(n_753),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_634),
.A2(n_649),
.B1(n_618),
.B2(n_599),
.Y(n_910)
);

OAI321xp33_ASAP7_75t_L g911 ( 
.A1(n_634),
.A2(n_649),
.A3(n_407),
.B1(n_661),
.B2(n_625),
.C(n_640),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_634),
.A2(n_649),
.B(n_620),
.C(n_753),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_653),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_637),
.Y(n_915)
);

BUFx8_ASAP7_75t_L g916 ( 
.A(n_677),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_620),
.B(n_608),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_753),
.A2(n_758),
.B(n_649),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_631),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_760),
.A2(n_724),
.B(n_776),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_637),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_637),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_774),
.A2(n_693),
.B(n_772),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_618),
.B(n_620),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_618),
.B(n_620),
.Y(n_926)
);

AND2x4_ASAP7_75t_SL g927 ( 
.A(n_647),
.B(n_524),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_616),
.B(n_492),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_760),
.A2(n_724),
.B(n_776),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_637),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_615),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_637),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_681),
.B(n_481),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_620),
.B(n_608),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_620),
.B(n_608),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_634),
.A2(n_649),
.B1(n_618),
.B2(n_599),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_637),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_620),
.B(n_608),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_628),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_774),
.A2(n_614),
.B(n_772),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_639),
.A2(n_640),
.B(n_407),
.C(n_608),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_620),
.B(n_608),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_620),
.B(n_608),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_773),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_910),
.A2(n_939),
.B1(n_906),
.B2(n_926),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_928),
.B(n_927),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_834),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_942),
.Y(n_951)
);

O2A1O1Ixp5_ASAP7_75t_L g952 ( 
.A1(n_918),
.A2(n_909),
.B(n_913),
.C(n_783),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_925),
.A2(n_926),
.B1(n_946),
.B2(n_945),
.Y(n_953)
);

OAI21x1_ASAP7_75t_SL g954 ( 
.A1(n_908),
.A2(n_929),
.B(n_920),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_786),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_925),
.A2(n_911),
.B(n_944),
.C(n_777),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_852),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_779),
.A2(n_924),
.B(n_912),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_942),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_828),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_787),
.A2(n_789),
.B(n_781),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_919),
.B(n_782),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_919),
.B(n_917),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_930),
.A2(n_933),
.B(n_931),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_943),
.A2(n_872),
.B(n_897),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_937),
.B(n_938),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_796),
.A2(n_874),
.B(n_823),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_854),
.A2(n_902),
.B(n_865),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_880),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_814),
.A2(n_887),
.B(n_820),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_880),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_880),
.B(n_871),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_941),
.B(n_866),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_916),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_859),
.A2(n_936),
.B1(n_804),
.B2(n_801),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_944),
.A2(n_777),
.B(n_861),
.C(n_801),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_802),
.A2(n_793),
.B(n_812),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_880),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_890),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_798),
.A2(n_860),
.B(n_778),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_916),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_877),
.B(n_869),
.Y(n_982)
);

AO31x2_ASAP7_75t_L g983 ( 
.A1(n_899),
.A2(n_857),
.A3(n_878),
.B(n_800),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_799),
.Y(n_984)
);

AND2x6_ASAP7_75t_L g985 ( 
.A(n_851),
.B(n_881),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_824),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_899),
.A2(n_800),
.A3(n_885),
.B(n_867),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_826),
.A2(n_895),
.B(n_791),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_901),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_903),
.Y(n_990)
);

AO31x2_ASAP7_75t_L g991 ( 
.A1(n_809),
.A2(n_810),
.A3(n_803),
.B(n_858),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_894),
.A2(n_853),
.B(n_806),
.Y(n_992)
);

AOI21x1_ASAP7_75t_SL g993 ( 
.A1(n_838),
.A2(n_818),
.B(n_889),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_816),
.A2(n_817),
.B(n_790),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_883),
.A2(n_842),
.B(n_784),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_879),
.B(n_863),
.Y(n_996)
);

AOI221xp5_ASAP7_75t_L g997 ( 
.A1(n_832),
.A2(n_819),
.B1(n_859),
.B2(n_836),
.C(n_835),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_905),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_860),
.A2(n_904),
.B(n_827),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_825),
.B(n_932),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_841),
.B(n_855),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_805),
.A2(n_896),
.B(n_829),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_785),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_840),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_780),
.A2(n_819),
.B(n_870),
.C(n_788),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_830),
.A2(n_873),
.B1(n_813),
.B2(n_875),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_833),
.A2(n_837),
.B(n_843),
.Y(n_1007)
);

BUFx4_ASAP7_75t_R g1008 ( 
.A(n_847),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_788),
.A2(n_808),
.B(n_815),
.C(n_892),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_848),
.B(n_922),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_915),
.B(n_921),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_935),
.B(n_940),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_839),
.A2(n_850),
.B(n_844),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_785),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_875),
.A2(n_822),
.B1(n_851),
.B2(n_888),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_811),
.A2(n_886),
.B(n_898),
.Y(n_1016)
);

BUFx4_ASAP7_75t_SL g1017 ( 
.A(n_856),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_868),
.B(n_864),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_876),
.B(n_891),
.Y(n_1019)
);

BUFx5_ASAP7_75t_L g1020 ( 
.A(n_907),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_795),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_862),
.A2(n_815),
.B(n_884),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_900),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_795),
.A2(n_914),
.B(n_884),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_849),
.A2(n_934),
.B(n_846),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_821),
.A2(n_893),
.B(n_947),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_822),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_845),
.A2(n_792),
.B(n_831),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_795),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_914),
.A2(n_939),
.B(n_910),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_910),
.A2(n_939),
.B(n_913),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_786),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_909),
.A2(n_913),
.B(n_939),
.C(n_910),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_880),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_779),
.A2(n_923),
.B(n_814),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_880),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_925),
.B(n_926),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_786),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_828),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_882),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_925),
.B(n_926),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_909),
.A2(n_913),
.B(n_779),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_906),
.B(n_911),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_911),
.B(n_625),
.C(n_634),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_787),
.A2(n_789),
.B(n_910),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_787),
.A2(n_789),
.B(n_910),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_925),
.B(n_926),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1051)
);

BUFx8_ASAP7_75t_L g1052 ( 
.A(n_882),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_787),
.A2(n_789),
.B(n_910),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_786),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_927),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_925),
.B(n_926),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_928),
.B(n_400),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_918),
.A2(n_779),
.A3(n_798),
.B(n_794),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_925),
.B(n_926),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_909),
.A2(n_913),
.B1(n_939),
.B2(n_910),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_925),
.B(n_926),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_787),
.A2(n_789),
.B(n_910),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_918),
.A2(n_779),
.A3(n_798),
.B(n_794),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_925),
.B(n_926),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_880),
.B(n_669),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_909),
.A2(n_913),
.B(n_939),
.C(n_910),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_906),
.B(n_911),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_779),
.A2(n_923),
.B(n_814),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_786),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_910),
.A2(n_939),
.B1(n_649),
.B2(n_634),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_786),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_925),
.B(n_926),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_925),
.B(n_926),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_910),
.A2(n_939),
.B1(n_649),
.B2(n_634),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_786),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_909),
.A2(n_913),
.B(n_779),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_910),
.A2(n_939),
.B(n_913),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_925),
.B(n_926),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_797),
.A2(n_807),
.B(n_923),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_925),
.B(n_926),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1075),
.A2(n_1081),
.B(n_1032),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1052),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1047),
.B(n_1062),
.C(n_997),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_951),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_1034),
.A2(n_1071),
.B(n_1085),
.C(n_1032),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1000),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1039),
.B(n_1043),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_972),
.B(n_1003),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1039),
.B(n_1043),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1085),
.A2(n_1062),
.B(n_1049),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1000),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1001),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_948),
.A2(n_956),
.B(n_997),
.C(n_1056),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1048),
.A2(n_1067),
.B(n_1053),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_972),
.B(n_1014),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1050),
.B(n_1056),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1001),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1008),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1059),
.B(n_963),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1050),
.A2(n_1088),
.B1(n_1086),
.B2(n_1079),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1010),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_962),
.B(n_1061),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_961),
.A2(n_1045),
.B(n_1083),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1010),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1061),
.A2(n_1088),
.B(n_1064),
.C(n_1069),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1052),
.Y(n_1114)
);

CKINVDCx8_ASAP7_75t_R g1115 ( 
.A(n_990),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1064),
.A2(n_1079),
.B1(n_1086),
.B2(n_1069),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1046),
.A2(n_1072),
.B1(n_1078),
.B2(n_953),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1078),
.B(n_953),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_959),
.B(n_982),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1041),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1038),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_949),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_950),
.B(n_973),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1017),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1004),
.B(n_985),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_974),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_973),
.B(n_966),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1027),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_981),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_985),
.A2(n_1028),
.B1(n_954),
.B2(n_989),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1045),
.A2(n_1083),
.B(n_958),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_966),
.A2(n_975),
.B1(n_976),
.B2(n_1028),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_985),
.B(n_971),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_1070),
.B(n_957),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_996),
.B(n_1019),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_SL g1136 ( 
.A(n_1018),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1042),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_985),
.A2(n_1015),
.B1(n_1055),
.B2(n_1006),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_996),
.B(n_1019),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_955),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1011),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1023),
.B(n_1011),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_952),
.A2(n_1005),
.B(n_1009),
.C(n_1030),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1012),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1018),
.B(n_998),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1023),
.B(n_1012),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_989),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_984),
.B(n_986),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1033),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_R g1151 ( 
.A(n_969),
.B(n_1035),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1040),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1054),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_979),
.B(n_983),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1021),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1074),
.A2(n_1082),
.B(n_1077),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_979),
.B(n_983),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_1021),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_995),
.A2(n_964),
.B(n_980),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_980),
.A2(n_1013),
.B(n_1007),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1021),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_1024),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1029),
.B(n_1020),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1029),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1020),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1024),
.B(n_1026),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_994),
.A2(n_992),
.B(n_1036),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1020),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_L g1169 ( 
.A(n_1025),
.B(n_970),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1016),
.B(n_999),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_987),
.B(n_1002),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1020),
.A2(n_987),
.B1(n_965),
.B2(n_968),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_993),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_991),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_967),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1031),
.A2(n_1087),
.B(n_1065),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1044),
.A2(n_1084),
.B(n_1063),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1051),
.A2(n_1080),
.B(n_1058),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1060),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1037),
.A2(n_1073),
.B1(n_1060),
.B2(n_1068),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1068),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_991),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_988),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1057),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1066),
.A2(n_1076),
.B(n_977),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_960),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1059),
.B(n_628),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1047),
.A2(n_582),
.B1(n_649),
.B2(n_634),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1039),
.B(n_1056),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1000),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1032),
.A2(n_1085),
.B(n_1062),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1000),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1047),
.A2(n_649),
.B1(n_634),
.B2(n_910),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_974),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_951),
.B(n_928),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_978),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1032),
.A2(n_1085),
.B(n_1062),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1039),
.B(n_481),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_1081),
.B(n_1032),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1059),
.B(n_628),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1032),
.A2(n_1085),
.B(n_1062),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1017),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_985),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_974),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1000),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_954),
.A2(n_918),
.B(n_1075),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1039),
.B(n_1056),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1052),
.Y(n_1208)
);

BUFx4f_ASAP7_75t_L g1209 ( 
.A(n_974),
.Y(n_1209)
);

INVx3_ASAP7_75t_SL g1210 ( 
.A(n_981),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1003),
.B(n_880),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1059),
.B(n_628),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1075),
.A2(n_632),
.B1(n_647),
.B2(n_544),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1000),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1047),
.A2(n_582),
.B1(n_649),
.B2(n_634),
.Y(n_1215)
);

BUFx5_ASAP7_75t_L g1216 ( 
.A(n_985),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1017),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_972),
.B(n_880),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_972),
.B(n_880),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1047),
.A2(n_649),
.B1(n_634),
.B2(n_910),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1039),
.B(n_481),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1052),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_972),
.B(n_880),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1213),
.A2(n_1108),
.B1(n_1203),
.B2(n_1217),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1149),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1097),
.B(n_1116),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1195),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1102),
.A2(n_1160),
.B(n_1159),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1188),
.A2(n_1215),
.B1(n_1091),
.B2(n_1221),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1140),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1107),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1089),
.B(n_1199),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1158),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1193),
.A2(n_1117),
.B1(n_1101),
.B2(n_1118),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1089),
.A2(n_1199),
.B(n_1144),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1152),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1179),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1118),
.B(n_1110),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1185),
.A2(n_1178),
.B(n_1177),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1153),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_SL g1242 ( 
.A(n_1090),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1203),
.B(n_1133),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1203),
.A2(n_1216),
.B1(n_1132),
.B2(n_1116),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1150),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1216),
.A2(n_1132),
.B1(n_1222),
.B2(n_1198),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1171),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1191),
.A2(n_1197),
.B(n_1201),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1104),
.B(n_1189),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1216),
.A2(n_1130),
.B1(n_1138),
.B2(n_1187),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1216),
.A2(n_1200),
.B1(n_1212),
.B2(n_1123),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1125),
.A2(n_1207),
.B1(n_1189),
.B2(n_1104),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1154),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1154),
.B(n_1157),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1165),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1185),
.A2(n_1167),
.B(n_1177),
.Y(n_1256)
);

CKINVDCx14_ASAP7_75t_R g1257 ( 
.A(n_1194),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1094),
.B(n_1099),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1157),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1181),
.Y(n_1260)
);

BUFx4f_ASAP7_75t_SL g1261 ( 
.A(n_1204),
.Y(n_1261)
);

BUFx8_ASAP7_75t_SL g1262 ( 
.A(n_1209),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1128),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1223),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1216),
.A2(n_1123),
.B1(n_1119),
.B2(n_1148),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1171),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1100),
.B(n_1105),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1156),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1142),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1148),
.A2(n_1136),
.B1(n_1186),
.B2(n_1120),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1129),
.Y(n_1271)
);

BUFx4f_ASAP7_75t_SL g1272 ( 
.A(n_1126),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1142),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1114),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_R g1276 ( 
.A1(n_1124),
.A2(n_1202),
.B1(n_1218),
.B2(n_1106),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1207),
.A2(n_1106),
.B1(n_1127),
.B2(n_1139),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1092),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1102),
.A2(n_1098),
.B(n_1111),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1137),
.Y(n_1280)
);

BUFx2_ASAP7_75t_SL g1281 ( 
.A(n_1136),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1113),
.A2(n_1197),
.B1(n_1191),
.B2(n_1201),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1168),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1127),
.A2(n_1131),
.B1(n_1098),
.B2(n_1095),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1135),
.A2(n_1139),
.B1(n_1147),
.B2(n_1190),
.Y(n_1285)
);

BUFx2_ASAP7_75t_R g1286 ( 
.A(n_1208),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1147),
.B(n_1135),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1131),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1206),
.A2(n_1145),
.B1(n_1141),
.B2(n_1214),
.Y(n_1289)
);

AO21x1_ASAP7_75t_SL g1290 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1093),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1192),
.B(n_1205),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1166),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1146),
.B(n_1163),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1122),
.A2(n_1115),
.B1(n_1210),
.B2(n_1134),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1166),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1143),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1096),
.A2(n_1103),
.B1(n_1173),
.B2(n_1224),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1175),
.A2(n_1180),
.B(n_1172),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1155),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1219),
.A2(n_1220),
.B1(n_1151),
.B2(n_1211),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1170),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1176),
.A2(n_1170),
.B(n_1162),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1170),
.Y(n_1303)
);

AO22x1_ASAP7_75t_L g1304 ( 
.A1(n_1168),
.A2(n_1161),
.B1(n_1196),
.B2(n_1121),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1164),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1121),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1149),
.Y(n_1308)
);

INVx4_ASAP7_75t_SL g1309 ( 
.A(n_1133),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1102),
.A2(n_1160),
.B(n_1159),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1149),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1203),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1165),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1154),
.B(n_1157),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1158),
.Y(n_1315)
);

INVx3_ASAP7_75t_SL g1316 ( 
.A(n_1129),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_SL g1317 ( 
.A1(n_1089),
.A2(n_1199),
.B(n_954),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1128),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1169),
.A2(n_1182),
.B(n_1174),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1149),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1149),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1149),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1149),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1149),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1223),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1128),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1160),
.A2(n_1185),
.B(n_1167),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1193),
.A2(n_1072),
.B(n_1046),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1247),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1254),
.B(n_1314),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1233),
.B(n_1239),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1264),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1260),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1247),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1302),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1233),
.B(n_1239),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1302),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1260),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1325),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1227),
.B(n_1249),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1325),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1288),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1266),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1254),
.B(n_1314),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1288),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1263),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1253),
.Y(n_1347)
);

BUFx2_ASAP7_75t_SL g1348 ( 
.A(n_1328),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1259),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1304),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1318),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1234),
.B(n_1315),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1259),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1326),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1296),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1264),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1236),
.B(n_1292),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1278),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1292),
.B(n_1295),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1280),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1295),
.B(n_1258),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1235),
.A2(n_1317),
.B1(n_1312),
.B2(n_1281),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1319),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1256),
.A2(n_1327),
.B(n_1279),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1258),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1267),
.B(n_1274),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1304),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1301),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1274),
.B(n_1226),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1283),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1301),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1283),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1303),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1303),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1299),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1248),
.A2(n_1282),
.B(n_1317),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1298),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1229),
.A2(n_1310),
.B(n_1284),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1283),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1230),
.A2(n_1289),
.B(n_1252),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1308),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1245),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1268),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1291),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1311),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1238),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1238),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1287),
.B(n_1285),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1255),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1231),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1237),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1324),
.Y(n_1395)
);

INVx4_ASAP7_75t_SL g1396 ( 
.A(n_1243),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1241),
.Y(n_1397)
);

INVx4_ASAP7_75t_SL g1398 ( 
.A(n_1243),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1305),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1269),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1273),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1298),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1229),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1240),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1331),
.B(n_1229),
.Y(n_1405)
);

OAI222xp33_ASAP7_75t_L g1406 ( 
.A1(n_1390),
.A2(n_1225),
.B1(n_1246),
.B2(n_1277),
.C1(n_1244),
.C2(n_1250),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1331),
.B(n_1310),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1348),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1340),
.B(n_1228),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1336),
.B(n_1310),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1333),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1336),
.B(n_1366),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1384),
.B(n_1265),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1329),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_SL g1415 ( 
.A(n_1362),
.B(n_1251),
.C(n_1297),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1366),
.B(n_1290),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1378),
.B(n_1290),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1365),
.B(n_1232),
.Y(n_1418)
);

OAI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1381),
.A2(n_1306),
.B(n_1257),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1369),
.B(n_1293),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1333),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1381),
.B(n_1294),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1378),
.B(n_1293),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1384),
.B(n_1385),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1385),
.B(n_1255),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1403),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1338),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1377),
.B(n_1255),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1348),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1338),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1383),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1342),
.B(n_1313),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1330),
.B(n_1344),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1330),
.B(n_1234),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1396),
.B(n_1309),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1346),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1351),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1345),
.B(n_1307),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1347),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1361),
.B(n_1315),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1354),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1355),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1376),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1419),
.B(n_1350),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1446)
);

OAI221xp5_ASAP7_75t_L g1447 ( 
.A1(n_1422),
.A2(n_1419),
.B1(n_1413),
.B2(n_1415),
.C(n_1402),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1422),
.B(n_1358),
.C(n_1360),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1406),
.A2(n_1257),
.B(n_1417),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1435),
.A2(n_1341),
.B1(n_1339),
.B2(n_1343),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1413),
.A2(n_1402),
.B1(n_1367),
.B2(n_1400),
.C(n_1401),
.Y(n_1451)
);

NOR3xp33_ASAP7_75t_L g1452 ( 
.A(n_1406),
.B(n_1391),
.C(n_1352),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1417),
.A2(n_1379),
.B(n_1300),
.Y(n_1453)
);

OAI21xp33_ASAP7_75t_L g1454 ( 
.A1(n_1426),
.A2(n_1382),
.B(n_1395),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1444),
.B(n_1370),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1408),
.A2(n_1364),
.B(n_1404),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1415),
.A2(n_1400),
.B1(n_1401),
.B2(n_1374),
.C(n_1368),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1409),
.A2(n_1375),
.B1(n_1372),
.B2(n_1368),
.C(n_1374),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1409),
.A2(n_1386),
.B1(n_1270),
.B2(n_1375),
.C(n_1372),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1442),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1437),
.B(n_1404),
.C(n_1373),
.D(n_1371),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1412),
.B(n_1334),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1408),
.A2(n_1357),
.B1(n_1392),
.B2(n_1388),
.C(n_1344),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1437),
.B(n_1388),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1405),
.B(n_1410),
.Y(n_1465)
);

NAND4xp25_ASAP7_75t_L g1466 ( 
.A(n_1438),
.B(n_1371),
.C(n_1380),
.D(n_1373),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_L g1467 ( 
.A(n_1430),
.B(n_1349),
.C(n_1353),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1423),
.A2(n_1276),
.B1(n_1387),
.B2(n_1389),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1417),
.A2(n_1379),
.B(n_1332),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1405),
.B(n_1410),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1423),
.B(n_1343),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1423),
.B(n_1359),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_SL g1474 ( 
.A1(n_1429),
.A2(n_1335),
.B(n_1337),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1399),
.C(n_1363),
.Y(n_1475)
);

OAI21xp33_ASAP7_75t_L g1476 ( 
.A1(n_1407),
.A2(n_1433),
.B(n_1439),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1441),
.B(n_1359),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1411),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_1359),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1435),
.A2(n_1418),
.B1(n_1420),
.B2(n_1434),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1424),
.A2(n_1393),
.B1(n_1397),
.B2(n_1394),
.C(n_1418),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_R g1483 ( 
.A(n_1418),
.B(n_1356),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1445),
.B(n_1425),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1456),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1465),
.B(n_1425),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1478),
.B(n_1411),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1478),
.B(n_1421),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1456),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1456),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1476),
.B(n_1407),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1446),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1456),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1471),
.B(n_1416),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1476),
.B(n_1421),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1482),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1481),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1448),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1467),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1467),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1480),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1448),
.B(n_1431),
.C(n_1424),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1455),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1425),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1464),
.B(n_1431),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1454),
.B(n_1440),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1451),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1483),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1461),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1475),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1503),
.B(n_1480),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1503),
.B(n_1462),
.Y(n_1518)
);

OAI21xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1500),
.A2(n_1466),
.B(n_1462),
.Y(n_1519)
);

AND2x2_ASAP7_75t_SL g1520 ( 
.A(n_1511),
.B(n_1425),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1488),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1503),
.B(n_1472),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1496),
.B(n_1469),
.Y(n_1524)
);

NAND2xp33_ASAP7_75t_R g1525 ( 
.A(n_1510),
.B(n_1436),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1501),
.B(n_1458),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1502),
.B(n_1457),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1472),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1507),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1503),
.B(n_1470),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1507),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1432),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1486),
.B(n_1474),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1504),
.A2(n_1449),
.B(n_1447),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1499),
.B(n_1463),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1490),
.Y(n_1538)
);

NOR2x1p5_ASAP7_75t_SL g1539 ( 
.A(n_1485),
.B(n_1427),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1486),
.B(n_1477),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1497),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1512),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1477),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1485),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1485),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1490),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1489),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1486),
.B(n_1479),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1510),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1316),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1534),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1511),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1509),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1520),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1523),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1551),
.B(n_1316),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1536),
.A2(n_1509),
.B(n_1511),
.C(n_1504),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1520),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1550),
.B(n_1486),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1515),
.B(n_1527),
.Y(n_1562)
);

NOR2x1_ASAP7_75t_L g1563 ( 
.A(n_1550),
.B(n_1490),
.Y(n_1563)
);

NOR2x1p5_ASAP7_75t_SL g1564 ( 
.A(n_1526),
.B(n_1493),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_1498),
.Y(n_1565)
);

OAI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1542),
.A2(n_1498),
.B(n_1490),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1486),
.Y(n_1567)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1568 ( 
.A1(n_1536),
.A2(n_1495),
.B(n_1450),
.C(n_1459),
.D(n_1508),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1523),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1530),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1526),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1506),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1535),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1549),
.B(n_1506),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1508),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1549),
.B(n_1506),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1532),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1542),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1534),
.B(n_1492),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1541),
.B(n_1492),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1531),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_L g1585 ( 
.A(n_1531),
.B(n_1490),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1535),
.B(n_1506),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1505),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1513),
.B(n_1506),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1533),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1494),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1514),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1537),
.A2(n_1489),
.B1(n_1493),
.B2(n_1484),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1580),
.B(n_1537),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1562),
.B(n_1543),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1556),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1543),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1261),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1556),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1559),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1565),
.B(n_1514),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1577),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1577),
.B(n_1524),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1518),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1559),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1554),
.A2(n_1524),
.B1(n_1452),
.B2(n_1519),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1584),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1552),
.B(n_1516),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1559),
.B(n_1518),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1574),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1569),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1584),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1554),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1522),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1560),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.B(n_1522),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1566),
.C(n_1593),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1555),
.B(n_1529),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1575),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1569),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1560),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1574),
.B(n_1529),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1568),
.B(n_1519),
.C(n_1517),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1561),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1553),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1570),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1619),
.A2(n_1563),
.B(n_1566),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1599),
.A2(n_1585),
.B(n_1563),
.Y(n_1632)
);

AOI222xp33_ASAP7_75t_L g1633 ( 
.A1(n_1626),
.A2(n_1564),
.B1(n_1539),
.B2(n_1553),
.C1(n_1589),
.C2(n_1591),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_R g1634 ( 
.A1(n_1598),
.A2(n_1595),
.B1(n_1629),
.B2(n_1614),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1595),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1604),
.Y(n_1636)
);

OAI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1599),
.A2(n_1575),
.B(n_1585),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1575),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_SL g1639 ( 
.A(n_1600),
.B(n_1286),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1573),
.C(n_1571),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1609),
.B(n_1575),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1644)
);

INVxp33_ASAP7_75t_L g1645 ( 
.A(n_1621),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1621),
.A2(n_1547),
.B(n_1538),
.Y(n_1646)
);

O2A1O1Ixp5_ASAP7_75t_L g1647 ( 
.A1(n_1602),
.A2(n_1573),
.B(n_1571),
.C(n_1579),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1576),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1606),
.A2(n_1591),
.B1(n_1592),
.B2(n_1579),
.C(n_1583),
.Y(n_1649)
);

AOI32xp33_ASAP7_75t_L g1650 ( 
.A1(n_1605),
.A2(n_1489),
.A3(n_1493),
.B1(n_1547),
.B2(n_1538),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1597),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1601),
.A2(n_1489),
.B1(n_1548),
.B2(n_1546),
.C(n_1544),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1607),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1623),
.B(n_1581),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1601),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1607),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1634),
.A2(n_1628),
.B1(n_1612),
.B2(n_1620),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1641),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1633),
.A2(n_1612),
.B1(n_1628),
.B2(n_1276),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1643),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1651),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1649),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1638),
.B(n_1616),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1655),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1635),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1272),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1647),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1644),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1603),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1653),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1643),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1654),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1616),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1637),
.B1(n_1632),
.B2(n_1652),
.C(n_1650),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1657),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1668),
.A2(n_1564),
.B(n_1539),
.C(n_1645),
.Y(n_1679)
);

AOI222xp33_ASAP7_75t_L g1680 ( 
.A1(n_1676),
.A2(n_1645),
.B1(n_1646),
.B2(n_1630),
.C1(n_1627),
.C2(n_1613),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1668),
.A2(n_1630),
.B1(n_1627),
.B2(n_1613),
.C(n_1622),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1673),
.B(n_1663),
.C(n_1658),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_L g1683 ( 
.A(n_1661),
.B(n_1602),
.C(n_1622),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1666),
.B(n_1602),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1672),
.B(n_1618),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1660),
.A2(n_1612),
.B(n_1611),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1671),
.B(n_1625),
.C(n_1603),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1685),
.Y(n_1688)
);

NAND5xp2_ASAP7_75t_L g1689 ( 
.A(n_1677),
.B(n_1672),
.C(n_1670),
.D(n_1671),
.E(n_1664),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_SL g1690 ( 
.A(n_1678),
.B(n_1271),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1682),
.A2(n_1669),
.B1(n_1667),
.B2(n_1674),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1680),
.B(n_1675),
.Y(n_1692)
);

NOR4xp75_ASAP7_75t_L g1693 ( 
.A(n_1684),
.B(n_1606),
.C(n_1611),
.D(n_1618),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1665),
.B(n_1659),
.C(n_1662),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1687),
.B(n_1659),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1683),
.Y(n_1696)
);

NAND5xp2_ASAP7_75t_L g1697 ( 
.A(n_1681),
.B(n_1665),
.C(n_1624),
.D(n_1588),
.E(n_1576),
.Y(n_1697)
);

NAND5xp2_ASAP7_75t_L g1698 ( 
.A(n_1691),
.B(n_1686),
.C(n_1624),
.D(n_1262),
.E(n_1588),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1689),
.B(n_1572),
.C(n_1561),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1688),
.B(n_1620),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1692),
.B(n_1625),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1690),
.A2(n_1620),
.B(n_1592),
.C(n_1262),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1695),
.B(n_1583),
.Y(n_1703)
);

NOR2xp67_ASAP7_75t_L g1704 ( 
.A(n_1696),
.B(n_1697),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1703),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1701),
.B(n_1690),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1698),
.B(n_1271),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1704),
.B(n_1694),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1699),
.A2(n_1594),
.B1(n_1582),
.B2(n_1572),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1700),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1706),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1710),
.Y(n_1713)
);

NAND2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1708),
.B(n_1275),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1705),
.Y(n_1715)
);

NOR2xp67_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1711),
.Y(n_1716)
);

XOR2xp5_ASAP7_75t_L g1717 ( 
.A(n_1714),
.B(n_1712),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1715),
.B(n_1709),
.C(n_1242),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1713),
.B(n_1716),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1719),
.Y(n_1720)
);

OAI211xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1720),
.A2(n_1718),
.B(n_1717),
.C(n_1693),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1594),
.B1(n_1582),
.B2(n_1561),
.Y(n_1722)
);

OR3x2_ASAP7_75t_L g1723 ( 
.A(n_1721),
.B(n_1275),
.C(n_1242),
.Y(n_1723)
);

OA22x2_ASAP7_75t_L g1724 ( 
.A1(n_1722),
.A2(n_1594),
.B1(n_1582),
.B2(n_1572),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1723),
.A2(n_1548),
.B(n_1546),
.Y(n_1725)
);

AOI21xp33_ASAP7_75t_SL g1726 ( 
.A1(n_1724),
.A2(n_1242),
.B(n_1546),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1548),
.B1(n_1587),
.B2(n_1525),
.Y(n_1727)
);

AOI32xp33_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1590),
.A3(n_1578),
.B1(n_1567),
.B2(n_1517),
.Y(n_1728)
);

AOI322xp5_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1727),
.A3(n_1521),
.B1(n_1468),
.B2(n_1590),
.C1(n_1578),
.C2(n_1567),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1521),
.B1(n_1545),
.B2(n_1281),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1545),
.B(n_1491),
.C(n_1453),
.Y(n_1731)
);


endmodule