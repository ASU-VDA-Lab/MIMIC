module fake_netlist_1_7033_n_730 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_730);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_730;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_638;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp33_ASAP7_75t_L g82 ( .A(n_34), .B(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_44), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_54), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_21), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_39), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_72), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_23), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_57), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_51), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_78), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_2), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_73), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
XOR2xp5_ASAP7_75t_L g107 ( .A(n_80), .B(n_61), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_35), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_38), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_77), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_30), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_24), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_3), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_26), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_17), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_56), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_18), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_52), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_37), .Y(n_123) );
BUFx5_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_42), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_69), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_19), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_43), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_17), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_20), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
OR2x6_ASAP7_75t_L g133 ( .A(n_105), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_84), .B(n_36), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_124), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_88), .B(n_0), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_118), .B(n_1), .Y(n_140) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_102), .A2(n_45), .B(n_79), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_95), .B(n_2), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_90), .B(n_3), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
XNOR2xp5_ASAP7_75t_L g147 ( .A(n_131), .B(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
INVx6_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_102), .A2(n_46), .B(n_76), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_91), .B(n_5), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_108), .B(n_5), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_95), .B(n_6), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_104), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_121), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_115), .B(n_7), .Y(n_158) );
INVxp67_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_115), .B(n_8), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_94), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_126), .B(n_9), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
AOI22xp5_ASAP7_75t_SL g165 ( .A1(n_121), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_93), .Y(n_166) );
INVxp67_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_96), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_86), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_130), .A2(n_103), .B1(n_86), .B2(n_129), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_85), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_129), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_85), .B(n_15), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_98), .B(n_59), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_131), .A2(n_16), .B1(n_19), .B2(n_21), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_127), .B1(n_125), .B2(n_100), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_146), .B(n_111), .C(n_101), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_156), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_172), .B(n_112), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_144), .B(n_109), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_133), .A2(n_112), .B1(n_123), .B2(n_113), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_172), .B(n_113), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_135), .B(n_123), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_110), .B(n_122), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_156), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
OR2x6_ASAP7_75t_L g193 ( .A(n_133), .B(n_107), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_135), .B(n_119), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_143), .B(n_117), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_143), .B(n_120), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
BUFx10_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_158), .A2(n_120), .B1(n_99), .B2(n_97), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_155), .B(n_94), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_146), .B(n_124), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_174), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_148), .B(n_124), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_159), .B(n_124), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_148), .B(n_82), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_133), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_163), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_149), .B(n_16), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
BUFx10_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_161), .A2(n_28), .B1(n_29), .B2(n_40), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_149), .B(n_49), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
INVx8_ASAP7_75t_L g222 ( .A(n_133), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_132), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_171), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_150), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_174), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_150), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_160), .B(n_50), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_162), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_167), .B(n_160), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_166), .B(n_53), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_141), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_134), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_166), .B(n_58), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_162), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_168), .B(n_60), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_168), .B(n_62), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_175), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_134), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_154), .B(n_66), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_175), .A2(n_68), .B1(n_70), .B2(n_71), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_183), .B(n_163), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_204), .A2(n_139), .B1(n_140), .B2(n_173), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_209), .B(n_153), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_228), .B(n_152), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_228), .B(n_137), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_232), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_232), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_180), .B(n_136), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_222), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_234), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_188), .B(n_151), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_211), .B(n_147), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_231), .A2(n_136), .B(n_141), .C(n_151), .Y(n_259) );
AND2x2_ASAP7_75t_SL g260 ( .A(n_226), .B(n_170), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_226), .B(n_206), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_222), .A2(n_151), .B1(n_141), .B2(n_176), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_222), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_235), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_193), .A2(n_165), .B1(n_157), .B2(n_147), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_185), .B(n_141), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_201), .B(n_151), .C(n_162), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_206), .B(n_162), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_186), .B(n_81), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_200), .B(n_162), .Y(n_271) );
AO22x1_ASAP7_75t_L g272 ( .A1(n_179), .A2(n_164), .B1(n_191), .B2(n_222), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_194), .B(n_164), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_241), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_200), .B(n_164), .Y(n_275) );
INVx8_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_241), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_188), .B(n_164), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_200), .B(n_164), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_187), .Y(n_280) );
INVx8_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_196), .B(n_182), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_217), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_187), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_217), .B(n_190), .Y(n_285) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_202), .B(n_190), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_182), .B(n_177), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_182), .A2(n_188), .B1(n_197), .B2(n_184), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_184), .B(n_190), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_217), .Y(n_290) );
NOR2x2_ASAP7_75t_L g291 ( .A(n_193), .B(n_224), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_208), .B(n_212), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_187), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_210), .B(n_212), .Y(n_294) );
NOR2xp33_ASAP7_75t_SL g295 ( .A(n_234), .B(n_227), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_202), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_210), .B(n_212), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_SL g298 ( .A1(n_229), .A2(n_233), .B(n_238), .C(n_210), .Y(n_298) );
INVx8_ASAP7_75t_L g299 ( .A(n_202), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_202), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_224), .A2(n_179), .B1(n_191), .B2(n_193), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_189), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_192), .B(n_207), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_214), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_203), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_193), .B(n_178), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_227), .B(n_225), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_192), .B(n_207), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_227), .B(n_178), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_242), .B(n_219), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_189), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_240), .A2(n_243), .B1(n_199), .B2(n_195), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_287), .A2(n_218), .B1(n_236), .B2(n_239), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_256), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_283), .B(n_199), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_246), .B(n_225), .Y(n_320) );
OAI22xp5_ASAP7_75t_SL g321 ( .A1(n_265), .A2(n_215), .B1(n_220), .B2(n_213), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_282), .B(n_215), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_244), .A2(n_195), .B(n_213), .C(n_220), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_305), .B(n_230), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_257), .A2(n_221), .B(n_223), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_261), .B(n_230), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_261), .B(n_230), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_257), .A2(n_221), .B(n_223), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_264), .B(n_230), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_245), .A2(n_230), .B1(n_237), .B2(n_216), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g332 ( .A1(n_253), .A2(n_237), .B(n_198), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g333 ( .A(n_265), .B(n_230), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_292), .A2(n_181), .B(n_198), .C(n_216), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_307), .A2(n_216), .B1(n_181), .B2(n_198), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_262), .B(n_181), .C(n_198), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_276), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_254), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_255), .B(n_181), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_293), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_307), .A2(n_216), .B1(n_181), .B2(n_198), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_301), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_263), .B(n_216), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_266), .A2(n_298), .B(n_259), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_288), .A2(n_294), .B1(n_247), .B2(n_277), .C(n_274), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_267), .B(n_309), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_258), .B(n_260), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_276), .B(n_281), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_314), .A2(n_304), .B1(n_309), .B2(n_283), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_280), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_302), .B(n_290), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_247), .B(n_249), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_256), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_268), .A2(n_278), .B(n_295), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_284), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_312), .A2(n_256), .B1(n_306), .B2(n_301), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_291), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_300), .B(n_295), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_248), .B(n_250), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_281), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_289), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_300), .B(n_296), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_278), .A2(n_269), .B(n_249), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_L g366 ( .A1(n_310), .A2(n_285), .B(n_273), .C(n_251), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_303), .A2(n_313), .B1(n_252), .B2(n_281), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_272), .B(n_270), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_311), .B(n_286), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_299), .B(n_300), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
AO31x2_ASAP7_75t_L g372 ( .A1(n_345), .A2(n_308), .A3(n_311), .B(n_279), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_348), .A2(n_311), .B(n_275), .Y(n_373) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_356), .A2(n_271), .A3(n_299), .B(n_351), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_299), .B1(n_333), .B2(n_347), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_356), .A2(n_336), .B(n_347), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_354), .A2(n_319), .B1(n_363), .B2(n_321), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_365), .A2(n_323), .B(n_324), .C(n_368), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_365), .A2(n_316), .B(n_329), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_326), .A2(n_325), .B(n_361), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_325), .A2(n_361), .B(n_330), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g383 ( .A1(n_366), .A2(n_353), .B(n_357), .C(n_334), .Y(n_383) );
NAND3xp33_ASAP7_75t_SL g384 ( .A(n_359), .B(n_349), .C(n_369), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_327), .B(n_328), .Y(n_385) );
OAI22x1_ASAP7_75t_L g386 ( .A1(n_318), .A2(n_369), .B1(n_341), .B2(n_320), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_355), .B(n_358), .Y(n_387) );
AO21x1_ASAP7_75t_L g388 ( .A1(n_331), .A2(n_360), .B(n_330), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_340), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_322), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_338), .B(n_337), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_332), .A2(n_317), .B(n_343), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_335), .A2(n_367), .B(n_364), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_342), .B(n_344), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_339), .A2(n_343), .B(n_355), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_342), .A2(n_362), .B1(n_350), .B2(n_370), .C(n_344), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_339), .A2(n_347), .B(n_244), .C(n_282), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_350), .A2(n_345), .B(n_365), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_355), .A2(n_346), .B1(n_348), .B2(n_347), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_346), .A2(n_348), .B1(n_347), .B2(n_351), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_346), .B(n_204), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_346), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_345), .A2(n_329), .B(n_326), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_380), .B(n_379), .C(n_400), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_402), .A2(n_401), .B(n_375), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_378), .A2(n_384), .B1(n_385), .B2(n_377), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_371), .B(n_404), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_377), .B(n_403), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_405), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_389), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_382), .B(n_399), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_390), .B(n_398), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_386), .B1(n_373), .B2(n_383), .Y(n_416) );
INVx8_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_379), .A2(n_381), .B(n_383), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_391), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_376), .A2(n_388), .B(n_387), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_392), .B(n_395), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_395), .B(n_374), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_374), .B(n_372), .Y(n_424) );
BUFx12f_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_374), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_387), .A2(n_394), .B1(n_393), .B2(n_372), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_394), .A2(n_345), .B(n_380), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_372), .B(n_377), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_372), .B(n_346), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_380), .A2(n_345), .B(n_405), .Y(n_433) );
CKINVDCx11_ASAP7_75t_R g434 ( .A(n_390), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_399), .A2(n_333), .B(n_346), .C(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_432), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_412), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_432), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_431), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_425), .A2(n_408), .B1(n_410), .B2(n_422), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_435), .A2(n_407), .B(n_406), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_425), .A2(n_410), .B1(n_422), .B2(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_431), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_423), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_410), .A2(n_413), .B1(n_425), .B2(n_416), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_417), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_409), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_418), .A2(n_420), .B(n_430), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_411), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_416), .A2(n_414), .B(n_418), .C(n_428), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_409), .B(n_419), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_411), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_424), .B(n_428), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_424), .B(n_406), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
AOI211xp5_ASAP7_75t_SL g460 ( .A1(n_423), .A2(n_415), .B(n_414), .C(n_422), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_417), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_434), .B(n_422), .Y(n_463) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_420), .A2(n_430), .B(n_429), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_424), .B(n_426), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_433), .Y(n_467) );
AOI21xp5_ASAP7_75t_SL g468 ( .A1(n_415), .A2(n_426), .B(n_427), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_426), .A2(n_427), .B1(n_433), .B2(n_421), .C(n_417), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_427), .B(n_421), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_439), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_459), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_462), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_446), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_436), .B(n_433), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_447), .B(n_433), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_448), .A2(n_415), .B1(n_417), .B2(n_421), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_459), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_436), .B(n_415), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_448), .A2(n_417), .B1(n_444), .B2(n_442), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_440), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_463), .B(n_450), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_438), .B(n_440), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_447), .B(n_445), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
NOR2x1_ASAP7_75t_SL g490 ( .A(n_451), .B(n_449), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_467), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_454), .A2(n_443), .B(n_467), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_466), .B(n_458), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_445), .B(n_455), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_466), .Y(n_495) );
OAI222xp33_ASAP7_75t_L g496 ( .A1(n_450), .A2(n_469), .B1(n_465), .B2(n_455), .C1(n_456), .C2(n_453), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_466), .B(n_458), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_457), .B(n_458), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_458), .B(n_457), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_462), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_457), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_437), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_458), .B(n_457), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_443), .A2(n_470), .B(n_469), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_460), .B(n_471), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_470), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_460), .B(n_471), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_441), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_471), .B(n_452), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_441), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_451), .A2(n_449), .B1(n_462), .B2(n_471), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_461), .B(n_456), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_452), .B(n_464), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_449), .A2(n_451), .B1(n_462), .B2(n_453), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_452), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_495), .B(n_486), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_489), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_496), .B(n_468), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_493), .B(n_452), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_495), .B(n_452), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_493), .B(n_464), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_487), .B(n_464), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_487), .B(n_464), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_497), .B(n_464), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_479), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_497), .B(n_499), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_475), .B(n_477), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_499), .B(n_503), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_503), .B(n_476), .Y(n_535) );
INVx4_ASAP7_75t_L g536 ( .A(n_474), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_485), .B(n_494), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_476), .B(n_501), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_507), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_501), .B(n_504), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_504), .B(n_486), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_498), .B(n_510), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_494), .B(n_488), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_488), .B(n_491), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_475), .B(n_477), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_515), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_510), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_472), .B(n_484), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_498), .B(n_508), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_472), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_474), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_498), .B(n_512), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_491), .B(n_484), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_508), .B(n_505), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_478), .B(n_509), .Y(n_558) );
INVx3_ASAP7_75t_L g559 ( .A(n_507), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_474), .B(n_500), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_506), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_506), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_505), .B(n_478), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_516), .B(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_509), .Y(n_566) );
OR2x6_ASAP7_75t_L g567 ( .A(n_492), .B(n_512), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_502), .B(n_511), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_515), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_490), .B(n_482), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_482), .B(n_511), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_516), .B(n_507), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_560), .B(n_496), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_525), .B(n_535), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_507), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_551), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_537), .B(n_520), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_535), .B(n_520), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_565), .B(n_515), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_564), .B(n_513), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_564), .B(n_517), .Y(n_582) );
BUFx3_ASAP7_75t_L g583 ( .A(n_554), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_542), .B(n_480), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_542), .B(n_480), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_521), .B(n_519), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_538), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_517), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_533), .B(n_518), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_547), .B(n_519), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_538), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_565), .B(n_483), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_521), .B(n_514), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_544), .B(n_490), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_545), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_550), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_527), .B(n_474), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_474), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_544), .B(n_474), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_547), .B(n_474), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_500), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_522), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_556), .B(n_500), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_571), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_539), .B(n_500), .Y(n_609) );
NOR4xp25_ASAP7_75t_SL g610 ( .A(n_553), .B(n_500), .C(n_560), .D(n_566), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_567), .A2(n_500), .B1(n_523), .B2(n_553), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_554), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_568), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_571), .B(n_500), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_561), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_539), .B(n_546), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_562), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_523), .A2(n_572), .B(n_557), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_530), .B(n_532), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_546), .B(n_532), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_572), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_541), .B(n_531), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_534), .B(n_555), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_522), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_562), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_622), .B(n_567), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_613), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_606), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_577), .B(n_526), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_573), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_584), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_605), .B(n_531), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_578), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_588), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_611), .A2(n_570), .B1(n_536), .B2(n_567), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_592), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_621), .B(n_526), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_595), .Y(n_639) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_574), .B(n_536), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_622), .B(n_567), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_608), .B(n_541), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_606), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_598), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_575), .B(n_567), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_583), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_625), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_593), .B(n_552), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_625), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_593), .A2(n_555), .B1(n_557), .B2(n_552), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_587), .B(n_543), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_575), .B(n_555), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_615), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_617), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_620), .B(n_555), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_616), .B(n_549), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_583), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_579), .B(n_549), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_612), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_620), .B(n_543), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_611), .A2(n_536), .B1(n_548), .B2(n_558), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_580), .B(n_536), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_634), .B(n_624), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_628), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_629), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_661), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_647), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_652), .A2(n_619), .B1(n_585), .B2(n_586), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_631), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_631), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_SL g674 ( .A1(n_659), .A2(n_596), .B(n_609), .C(n_614), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_640), .A2(n_610), .B(n_601), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_638), .B(n_576), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_636), .A2(n_614), .B1(n_602), .B2(n_591), .Y(n_677) );
AOI211x1_ASAP7_75t_SL g678 ( .A1(n_664), .A2(n_607), .B(n_623), .C(n_558), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_665), .B(n_602), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_632), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_646), .B(n_654), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_629), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_632), .Y(n_683) );
INVxp33_ASAP7_75t_L g684 ( .A(n_665), .Y(n_684) );
AOI322xp5_ASAP7_75t_L g685 ( .A1(n_650), .A2(n_576), .A3(n_624), .B1(n_579), .B2(n_580), .C1(n_599), .C2(n_600), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_635), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_630), .B(n_581), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_638), .B(n_594), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_633), .A2(n_627), .B1(n_641), .B2(n_653), .C1(n_646), .C2(n_658), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_670), .A2(n_591), .B(n_627), .C(n_641), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_678), .B(n_662), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_667), .B(n_662), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_677), .A2(n_665), .B1(n_599), .B2(n_600), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_669), .B(n_657), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_677), .A2(n_663), .B1(n_645), .B2(n_655), .C(n_656), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_672), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_671), .A2(n_642), .B(n_630), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_685), .B(n_675), .C(n_689), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_674), .A2(n_660), .B(n_559), .C(n_540), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_684), .B(n_657), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_674), .A2(n_639), .B1(n_649), .B2(n_637), .C(n_635), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_673), .B(n_637), .C(n_639), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_688), .A2(n_679), .B1(n_666), .B2(n_676), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_680), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_697), .B(n_666), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_698), .A2(n_679), .B1(n_686), .B2(n_683), .C1(n_644), .C2(n_649), .Y(n_706) );
OAI21xp33_ASAP7_75t_SL g707 ( .A1(n_703), .A2(n_681), .B(n_654), .Y(n_707) );
AOI221x1_ASAP7_75t_L g708 ( .A1(n_691), .A2(n_644), .B1(n_682), .B2(n_668), .C(n_540), .Y(n_708) );
AOI221x1_ASAP7_75t_L g709 ( .A1(n_702), .A2(n_682), .B1(n_559), .B2(n_540), .C(n_626), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_701), .B(n_559), .C(n_540), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_694), .A2(n_687), .B(n_589), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_690), .A2(n_603), .B1(n_559), .B2(n_643), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g713 ( .A1(n_699), .A2(n_589), .B(n_581), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_710), .A2(n_695), .B1(n_693), .B2(n_696), .C(n_704), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_706), .A2(n_695), .B(n_700), .C(n_692), .Y(n_715) );
NOR4xp25_ASAP7_75t_L g716 ( .A(n_707), .B(n_651), .C(n_648), .D(n_643), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_708), .B(n_603), .C(n_529), .D(n_528), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g718 ( .A(n_705), .B(n_528), .C(n_529), .D(n_548), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_715), .Y(n_719) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_716), .B(n_712), .Y(n_720) );
NOR3xp33_ASAP7_75t_SL g721 ( .A(n_717), .B(n_711), .C(n_713), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_720), .Y(n_722) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_719), .A2(n_714), .B1(n_709), .B2(n_718), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_722), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_723), .B(n_721), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_721), .B1(n_651), .B2(n_648), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_726), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_727), .Y(n_728) );
OA22x2_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_724), .B1(n_569), .B2(n_563), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_582), .B1(n_566), .B2(n_590), .Y(n_730) );
endmodule