module fake_jpeg_30532_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_79),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_77),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_51),
.B1(n_53),
.B2(n_60),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_76),
.C(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_49),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_53),
.B1(n_50),
.B2(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_8),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_53),
.B1(n_55),
.B2(n_48),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_45),
.B1(n_4),
.B2(n_6),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_95),
.B1(n_9),
.B2(n_11),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_96),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_3),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_28),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_15),
.B(n_21),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_29),
.C(n_41),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.C(n_108),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_25),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_30),
.C(n_40),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_12),
.B1(n_43),
.B2(n_16),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_31),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_12),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_32),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_34),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_105),
.CI(n_110),
.CON(n_122),
.SN(n_122)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_23),
.C(n_14),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_133),
.B(n_115),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_103),
.B1(n_120),
.B2(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_22),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_137),
.B1(n_132),
.B2(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_129),
.B(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_122),
.C(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_124),
.B1(n_127),
.B2(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_136),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_142),
.B(n_124),
.Y(n_148)
);


endmodule