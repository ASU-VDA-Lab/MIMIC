module fake_jpeg_26073_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_34),
.Y(n_52)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_8),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_15),
.B1(n_28),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_39),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_15),
.B1(n_29),
.B2(n_16),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_36),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_29),
.B1(n_23),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_38),
.C(n_31),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_25),
.B(n_19),
.C(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_56),
.B1(n_64),
.B2(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_56),
.B1(n_44),
.B2(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_18),
.B1(n_17),
.B2(n_2),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_66),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_71),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_46),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_96),
.B(n_98),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_56),
.B1(n_58),
.B2(n_47),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_59),
.B(n_62),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_73),
.B1(n_70),
.B2(n_68),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_65),
.B1(n_18),
.B2(n_17),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_36),
.C(n_57),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_79),
.C(n_83),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_51),
.B1(n_61),
.B2(n_57),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_105),
.B1(n_81),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_62),
.B1(n_63),
.B2(n_18),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_81),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_90),
.C(n_95),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_83),
.B(n_81),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_122),
.B(n_126),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_88),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_115),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_66),
.B1(n_71),
.B2(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_97),
.B1(n_103),
.B2(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_11),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_139),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_108),
.B1(n_91),
.B2(n_21),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_90),
.A3(n_99),
.B1(n_95),
.B2(n_96),
.C1(n_103),
.C2(n_104),
.Y(n_135)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_117),
.A3(n_115),
.B1(n_119),
.B2(n_108),
.C1(n_110),
.C2(n_21),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_91),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_92),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_20),
.C(n_1),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_145),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_141),
.C(n_133),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_159),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_155),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_21),
.B1(n_20),
.B2(n_0),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_158),
.B1(n_163),
.B2(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_20),
.B1(n_0),
.B2(n_4),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_2),
.B(n_4),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_138),
.B(n_137),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_148),
.B1(n_144),
.B2(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_148),
.B1(n_146),
.B2(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_166),
.B1(n_153),
.B2(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

OAI31xp33_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_181),
.A3(n_137),
.B(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_151),
.C(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_183),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_136),
.C(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_155),
.C(n_157),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_193),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_181),
.B(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_129),
.C(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_167),
.B1(n_169),
.B2(n_158),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_191),
.B1(n_152),
.B2(n_177),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_128),
.B(n_179),
.C(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_199),
.B1(n_195),
.B2(n_202),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_202),
.B(n_188),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_198),
.B(n_10),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_182),
.C(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_190),
.B1(n_10),
.B2(n_11),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.Y(n_213)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_194),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_213),
.B1(n_214),
.B2(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_212),
.B(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_10),
.C(n_12),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_218),
.C(n_12),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_215),
.B(n_12),
.C(n_14),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_5),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_219),
.A2(n_221),
.B(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_14),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);


endmodule