module real_aes_16525_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_0), .A2(n_71), .B1(n_962), .B2(n_967), .Y(n_966) );
INVxp33_ASAP7_75t_SL g995 ( .A(n_0), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_1), .A2(n_5), .B1(n_1085), .B2(n_1088), .Y(n_1084) );
INVx1_ASAP7_75t_L g861 ( .A(n_2), .Y(n_861) );
INVx1_ASAP7_75t_L g774 ( .A(n_3), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_3), .A2(n_126), .B1(n_678), .B2(n_789), .C(n_796), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_4), .A2(n_186), .B1(n_442), .B2(n_913), .C(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g941 ( .A(n_4), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_6), .Y(n_1428) );
INVx1_ASAP7_75t_L g300 ( .A(n_7), .Y(n_300) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_7), .A2(n_87), .B1(n_392), .B2(n_393), .C(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g915 ( .A(n_8), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g943 ( .A1(n_8), .A2(n_132), .B1(n_567), .B2(n_695), .C(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g466 ( .A(n_9), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_9), .A2(n_103), .B1(n_298), .B2(n_516), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g878 ( .A1(n_10), .A2(n_606), .B(n_612), .Y(n_878) );
INVx1_ASAP7_75t_L g900 ( .A(n_10), .Y(n_900) );
INVxp67_ASAP7_75t_SL g1328 ( .A(n_11), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_11), .A2(n_25), .B1(n_345), .B2(n_1337), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_12), .A2(n_199), .B1(n_392), .B2(n_393), .C(n_414), .Y(n_455) );
OA222x2_ASAP7_75t_L g531 ( .A1(n_12), .A2(n_51), .B1(n_203), .B2(n_532), .C1(n_536), .C2(n_540), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_13), .A2(n_225), .B1(n_327), .B2(n_817), .C(n_819), .Y(n_816) );
INVx1_ASAP7_75t_L g838 ( .A(n_13), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_14), .Y(n_1381) );
INVx1_ASAP7_75t_L g259 ( .A(n_15), .Y(n_259) );
AND2x2_ASAP7_75t_L g302 ( .A(n_15), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g314 ( .A(n_15), .B(n_208), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_15), .B(n_269), .Y(n_494) );
INVx1_ASAP7_75t_L g573 ( .A(n_16), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_16), .A2(n_234), .B1(n_591), .B2(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g719 ( .A(n_17), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_17), .A2(n_36), .B1(n_679), .B2(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_18), .A2(n_108), .B1(n_637), .B2(n_639), .Y(n_636) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_18), .Y(n_687) );
INVx2_ASAP7_75t_L g1081 ( .A(n_19), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_19), .B(n_100), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_19), .B(n_1087), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_20), .A2(n_213), .B1(n_637), .B2(n_639), .Y(n_758) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_20), .Y(n_799) );
XNOR2x2_ASAP7_75t_L g907 ( .A(n_21), .B(n_908), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_21), .A2(n_216), .B1(n_1085), .B2(n_1088), .Y(n_1106) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_22), .Y(n_1389) );
INVx1_ASAP7_75t_L g652 ( .A(n_23), .Y(n_652) );
INVx1_ASAP7_75t_L g869 ( .A(n_24), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_24), .A2(n_127), .B1(n_306), .B2(n_569), .Y(n_895) );
INVxp67_ASAP7_75t_SL g1316 ( .A(n_25), .Y(n_1316) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_26), .A2(n_238), .B1(n_261), .B2(n_1413), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g1433 ( .A1(n_26), .A2(n_238), .B1(n_1363), .B2(n_1434), .Y(n_1433) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_27), .A2(n_78), .B1(n_604), .B2(n_608), .C(n_880), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_27), .A2(n_29), .B1(n_308), .B2(n_569), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g1038 ( .A(n_28), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g961 ( .A1(n_29), .A2(n_119), .B1(n_762), .B2(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g1290 ( .A(n_30), .Y(n_1290) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_31), .Y(n_1393) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_32), .A2(n_158), .B1(n_196), .B2(n_443), .C1(n_476), .C2(n_612), .Y(n_664) );
INVx1_ASAP7_75t_L g698 ( .A(n_32), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_33), .A2(n_241), .B1(n_1078), .B2(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g556 ( .A(n_34), .Y(n_556) );
INVx1_ASAP7_75t_L g972 ( .A(n_35), .Y(n_972) );
OA222x2_ASAP7_75t_L g985 ( .A1(n_35), .A2(n_148), .B1(n_245), .B2(n_532), .C1(n_540), .C2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g728 ( .A(n_36), .Y(n_728) );
INVx1_ASAP7_75t_L g725 ( .A(n_37), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_37), .A2(n_155), .B1(n_567), .B2(n_679), .Y(n_745) );
INVx1_ASAP7_75t_L g916 ( .A(n_38), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_38), .A2(n_75), .B1(n_937), .B2(n_938), .C(n_940), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_39), .A2(n_185), .B1(n_606), .B2(n_964), .C(n_965), .Y(n_963) );
INVx1_ASAP7_75t_L g1001 ( .A(n_39), .Y(n_1001) );
INVx1_ASAP7_75t_L g749 ( .A(n_40), .Y(n_749) );
INVx1_ASAP7_75t_L g823 ( .A(n_41), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_42), .A2(n_65), .B1(n_594), .B2(n_598), .C(n_635), .Y(n_926) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_42), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_43), .A2(n_224), .B1(n_1085), .B2(n_1088), .Y(n_1099) );
OAI21xp33_ASAP7_75t_L g558 ( .A1(n_44), .A2(n_532), .B(n_559), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_44), .A2(n_54), .B1(n_615), .B2(n_616), .C(n_618), .Y(n_614) );
AO22x1_ASAP7_75t_L g1103 ( .A1(n_45), .A2(n_59), .B1(n_1078), .B2(n_1082), .Y(n_1103) );
OAI211xp5_ASAP7_75t_SL g857 ( .A1(n_46), .A2(n_621), .B(n_858), .C(n_862), .Y(n_857) );
INVx1_ASAP7_75t_L g885 ( .A(n_46), .Y(n_885) );
INVx1_ASAP7_75t_L g1319 ( .A(n_47), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_47), .A2(n_117), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
XNOR2xp5_ASAP7_75t_L g1374 ( .A(n_48), .B(n_1375), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_49), .A2(n_106), .B1(n_761), .B2(n_763), .C(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g791 ( .A(n_49), .Y(n_791) );
INVx1_ASAP7_75t_L g360 ( .A(n_50), .Y(n_360) );
INVx1_ASAP7_75t_L g381 ( .A(n_50), .Y(n_381) );
INVx1_ASAP7_75t_L g453 ( .A(n_51), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_52), .A2(n_135), .B1(n_308), .B2(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g412 ( .A(n_52), .Y(n_412) );
INVx1_ASAP7_75t_L g576 ( .A(n_53), .Y(n_576) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_54), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_55), .A2(n_94), .B1(n_484), .B2(n_772), .C(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g798 ( .A(n_55), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_56), .A2(n_101), .B1(n_637), .B2(n_639), .C(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_56), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_57), .A2(n_140), .B1(n_643), .B2(n_645), .C(n_647), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_57), .A2(n_202), .B1(n_692), .B2(n_694), .C(n_696), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_58), .A2(n_228), .B1(n_594), .B2(n_598), .C(n_635), .Y(n_634) );
OAI21xp33_ASAP7_75t_SL g675 ( .A1(n_58), .A2(n_518), .B(n_540), .Y(n_675) );
INVx1_ASAP7_75t_L g253 ( .A(n_60), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_61), .A2(n_192), .B1(n_637), .B2(n_639), .Y(n_925) );
INVx1_ASAP7_75t_L g935 ( .A(n_61), .Y(n_935) );
INVx2_ASAP7_75t_L g367 ( .A(n_62), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g1390 ( .A(n_63), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_64), .A2(n_168), .B1(n_654), .B2(n_657), .Y(n_911) );
INVx1_ASAP7_75t_L g933 ( .A(n_64), .Y(n_933) );
INVx1_ASAP7_75t_L g952 ( .A(n_65), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_66), .A2(n_137), .B1(n_1301), .B2(n_1302), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_66), .A2(n_137), .B1(n_1360), .B2(n_1363), .Y(n_1359) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_67), .Y(n_807) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_67), .A2(n_598), .B(n_621), .C(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g1289 ( .A(n_68), .Y(n_1289) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_69), .A2(n_73), .B1(n_654), .B2(n_657), .Y(n_653) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_69), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_70), .A2(n_161), .B1(n_1078), .B2(n_1082), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g1002 ( .A(n_71), .Y(n_1002) );
AO221x2_ASAP7_75t_L g1170 ( .A1(n_72), .A2(n_198), .B1(n_1085), .B2(n_1088), .C(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g674 ( .A(n_73), .Y(n_674) );
INVx1_ASAP7_75t_L g775 ( .A(n_74), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_75), .A2(n_187), .B1(n_442), .B2(n_918), .C(n_920), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_76), .A2(n_162), .B1(n_327), .B2(n_333), .C(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g413 ( .A(n_76), .Y(n_413) );
INVx1_ASAP7_75t_L g633 ( .A(n_77), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_77), .A2(n_536), .B(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g991 ( .A1(n_78), .A2(n_185), .B1(n_333), .B2(n_992), .C(n_993), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_79), .Y(n_460) );
INVx1_ASAP7_75t_L g809 ( .A(n_80), .Y(n_809) );
INVx1_ASAP7_75t_L g470 ( .A(n_81), .Y(n_470) );
AOI221x1_ASAP7_75t_SL g495 ( .A1(n_81), .A2(n_93), .B1(n_327), .B2(n_337), .C(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_82), .A2(n_231), .B1(n_1415), .B2(n_1418), .Y(n_1414) );
OAI22xp33_ASAP7_75t_L g1441 ( .A1(n_82), .A2(n_231), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
INVx1_ASAP7_75t_L g979 ( .A(n_83), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_83), .B(n_706), .Y(n_983) );
INVx1_ASAP7_75t_L g726 ( .A(n_84), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_84), .A2(n_210), .B1(n_308), .B2(n_337), .Y(n_742) );
INVx1_ASAP7_75t_L g882 ( .A(n_85), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_86), .A2(n_123), .B1(n_608), .B2(n_871), .C(n_872), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_86), .A2(n_174), .B1(n_306), .B2(n_345), .Y(n_903) );
INVx1_ASAP7_75t_L g319 ( .A(n_87), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_88), .Y(n_715) );
INVx1_ASAP7_75t_L g448 ( .A(n_89), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_89), .A2(n_199), .B1(n_524), .B2(n_529), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_90), .A2(n_217), .B1(n_582), .B2(n_583), .Y(n_811) );
AOI21xp33_ASAP7_75t_L g841 ( .A1(n_90), .A2(n_484), .B(n_606), .Y(n_841) );
INVx1_ASAP7_75t_L g980 ( .A(n_91), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_91), .A2(n_165), .B1(n_526), .B2(n_575), .Y(n_1004) );
OAI221xp5_ASAP7_75t_L g284 ( .A1(n_92), .A2(n_247), .B1(n_285), .B2(n_287), .C(n_292), .Y(n_284) );
INVx1_ASAP7_75t_L g351 ( .A(n_92), .Y(n_351) );
INVx1_ASAP7_75t_L g486 ( .A(n_93), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_94), .A2(n_170), .B1(n_678), .B2(n_789), .C(n_790), .Y(n_788) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_95), .Y(n_255) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_95), .B(n_253), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_96), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_97), .A2(n_141), .B1(n_880), .B2(n_1033), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_97), .A2(n_98), .B1(n_306), .B2(n_569), .Y(n_1062) );
INVx1_ASAP7_75t_L g1044 ( .A(n_98), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_99), .A2(n_164), .B1(n_329), .B2(n_567), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_99), .A2(n_149), .B1(n_604), .B2(n_605), .C(n_606), .Y(n_603) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_100), .B(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1087 ( .A(n_100), .Y(n_1087) );
INVx1_ASAP7_75t_L g748 ( .A(n_101), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_102), .A2(n_1008), .B1(n_1009), .B2(n_1068), .Y(n_1007) );
INVx1_ASAP7_75t_L g1068 ( .A(n_102), .Y(n_1068) );
INVx1_ASAP7_75t_L g477 ( .A(n_103), .Y(n_477) );
INVx1_ASAP7_75t_L g311 ( .A(n_104), .Y(n_311) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_104), .A2(n_385), .B(n_389), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_105), .A2(n_139), .B1(n_654), .B2(n_657), .Y(n_770) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_105), .Y(n_801) );
INVx1_ASAP7_75t_L g797 ( .A(n_106), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_107), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g404 ( .A(n_107), .Y(n_404) );
INVx1_ASAP7_75t_L g432 ( .A(n_107), .Y(n_432) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_108), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_109), .A2(n_193), .B1(n_1078), .B2(n_1082), .Y(n_1077) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_110), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_110), .A2(n_123), .B1(n_890), .B2(n_892), .Y(n_889) );
XOR2xp5_ASAP7_75t_L g433 ( .A(n_111), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g1293 ( .A(n_112), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_113), .A2(n_279), .B1(n_280), .B2(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_113), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_114), .A2(n_235), .B1(n_343), .B2(n_569), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_114), .A2(n_191), .B1(n_390), .B2(n_604), .C(n_608), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_115), .Y(n_473) );
INVx1_ASAP7_75t_L g729 ( .A(n_116), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_116), .A2(n_167), .B1(n_293), .B2(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_SL g1311 ( .A(n_117), .Y(n_1311) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_118), .A2(n_173), .B1(n_594), .B2(n_598), .C(n_635), .Y(n_757) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_118), .A2(n_518), .B(n_540), .Y(n_784) );
INVxp67_ASAP7_75t_SL g994 ( .A(n_119), .Y(n_994) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_120), .A2(n_125), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g549 ( .A(n_120), .Y(n_549) );
INVx1_ASAP7_75t_L g924 ( .A(n_121), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_122), .A2(n_169), .B1(n_343), .B2(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g426 ( .A(n_122), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_124), .A2(n_855), .B1(n_905), .B2(n_906), .Y(n_854) );
INVx1_ASAP7_75t_L g906 ( .A(n_124), .Y(n_906) );
INVx1_ASAP7_75t_L g545 ( .A(n_125), .Y(n_545) );
INVx1_ASAP7_75t_L g767 ( .A(n_126), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_127), .A2(n_174), .B1(n_602), .B2(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g820 ( .A(n_128), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_128), .A2(n_201), .B1(n_602), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g863 ( .A(n_129), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_129), .A2(n_172), .B1(n_529), .B2(n_786), .C(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_130), .A2(n_190), .B1(n_343), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_130), .A2(n_235), .B1(n_390), .B2(n_602), .Y(n_601) );
AOI221xp5_ASAP7_75t_SL g326 ( .A1(n_131), .A2(n_150), .B1(n_327), .B2(n_333), .C(n_334), .Y(n_326) );
INVx1_ASAP7_75t_L g416 ( .A(n_131), .Y(n_416) );
INVx1_ASAP7_75t_L g921 ( .A(n_132), .Y(n_921) );
AO22x1_ASAP7_75t_L g1104 ( .A1(n_133), .A2(n_212), .B1(n_1085), .B2(n_1088), .Y(n_1104) );
BUFx3_ASAP7_75t_L g357 ( .A(n_134), .Y(n_357) );
INVx1_ASAP7_75t_L g428 ( .A(n_135), .Y(n_428) );
INVx1_ASAP7_75t_L g864 ( .A(n_136), .Y(n_864) );
INVx1_ASAP7_75t_L g756 ( .A(n_138), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_139), .A2(n_173), .B1(n_529), .B2(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_140), .B(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g1057 ( .A1(n_141), .A2(n_220), .B1(n_344), .B2(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g649 ( .A(n_142), .Y(n_649) );
INVx1_ASAP7_75t_L g825 ( .A(n_143), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_144), .A2(n_153), .B1(n_1085), .B2(n_1088), .Y(n_1131) );
INVx1_ASAP7_75t_L g1312 ( .A(n_145), .Y(n_1312) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_146), .Y(n_266) );
INVx1_ASAP7_75t_L g560 ( .A(n_147), .Y(n_560) );
INVx1_ASAP7_75t_L g982 ( .A(n_148), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_149), .A2(n_191), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g425 ( .A(n_150), .Y(n_425) );
INVx1_ASAP7_75t_L g1327 ( .A(n_151), .Y(n_1327) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_152), .Y(n_324) );
INVx1_ASAP7_75t_L g808 ( .A(n_154), .Y(n_808) );
INVx1_ASAP7_75t_L g718 ( .A(n_155), .Y(n_718) );
INVx1_ASAP7_75t_L g1281 ( .A(n_156), .Y(n_1281) );
INVx1_ASAP7_75t_L g1430 ( .A(n_157), .Y(n_1430) );
OAI211xp5_ASAP7_75t_L g1436 ( .A1(n_157), .A2(n_1357), .B(n_1437), .C(n_1439), .Y(n_1436) );
INVx1_ASAP7_75t_L g683 ( .A(n_158), .Y(n_683) );
INVx1_ASAP7_75t_L g1284 ( .A(n_159), .Y(n_1284) );
INVx1_ASAP7_75t_L g1025 ( .A(n_160), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_160), .A2(n_503), .B1(n_540), .B2(n_1060), .C(n_1063), .Y(n_1059) );
INVx1_ASAP7_75t_L g429 ( .A(n_162), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_163), .A2(n_226), .B1(n_1078), .B2(n_1082), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_164), .A2(n_190), .B1(n_602), .B2(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g971 ( .A(n_165), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_166), .Y(n_1382) );
INVx1_ASAP7_75t_L g722 ( .A(n_167), .Y(n_722) );
INVxp67_ASAP7_75t_SL g950 ( .A(n_168), .Y(n_950) );
INVx1_ASAP7_75t_L g422 ( .A(n_169), .Y(n_422) );
INVx1_ASAP7_75t_L g769 ( .A(n_170), .Y(n_769) );
INVx1_ASAP7_75t_L g1320 ( .A(n_171), .Y(n_1320) );
INVx1_ASAP7_75t_L g883 ( .A(n_172), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_175), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_176), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_177), .A2(n_222), .B1(n_1078), .B2(n_1082), .Y(n_1130) );
INVx1_ASAP7_75t_L g711 ( .A(n_178), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_178), .A2(n_180), .B1(n_526), .B2(n_575), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_179), .A2(n_1297), .B(n_1423), .C(n_1426), .Y(n_1422) );
INVx1_ASAP7_75t_L g1440 ( .A(n_179), .Y(n_1440) );
INVx1_ASAP7_75t_L g714 ( .A(n_180), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_181), .Y(n_463) );
XNOR2x1_ASAP7_75t_L g752 ( .A(n_182), .B(n_753), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g1395 ( .A(n_183), .Y(n_1395) );
INVx1_ASAP7_75t_L g1314 ( .A(n_184), .Y(n_1314) );
INVx1_ASAP7_75t_L g945 ( .A(n_186), .Y(n_945) );
INVx1_ASAP7_75t_L g947 ( .A(n_187), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_188), .Y(n_1387) );
AO22x1_ASAP7_75t_L g1120 ( .A1(n_189), .A2(n_218), .B1(n_1078), .B2(n_1121), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_192), .Y(n_929) );
CKINVDCx16_ASAP7_75t_R g1172 ( .A(n_194), .Y(n_1172) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_195), .A2(n_781), .B(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_195), .A2(n_214), .B1(n_637), .B2(n_639), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_196), .A2(n_297), .B(n_686), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_197), .A2(n_598), .B(n_623), .C(n_713), .Y(n_712) );
INVxp33_ASAP7_75t_SL g737 ( .A(n_197), .Y(n_737) );
INVx1_ASAP7_75t_L g804 ( .A(n_200), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_201), .A2(n_233), .B1(n_337), .B2(n_516), .Y(n_812) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_202), .A2(n_660), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g444 ( .A(n_203), .Y(n_444) );
INVx1_ASAP7_75t_L g1011 ( .A(n_204), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1017 ( .A(n_205), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_205), .A2(n_598), .B1(n_637), .B2(n_1035), .C(n_1042), .Y(n_1034) );
INVx1_ASAP7_75t_L g847 ( .A(n_206), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_207), .A2(n_230), .B1(n_1085), .B2(n_1088), .Y(n_1093) );
BUFx3_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
INVx1_ASAP7_75t_L g303 ( .A(n_208), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_209), .Y(n_1384) );
INVx1_ASAP7_75t_L g721 ( .A(n_210), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g1174 ( .A(n_211), .Y(n_1174) );
AOI222xp33_ASAP7_75t_L g1274 ( .A1(n_211), .A2(n_1275), .B1(n_1370), .B2(n_1373), .C1(n_1444), .C2(n_1446), .Y(n_1274) );
INVx1_ASAP7_75t_L g1005 ( .A(n_212), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_213), .Y(n_779) );
INVxp33_ASAP7_75t_L g827 ( .A(n_214), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_215), .A2(n_606), .B(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1055 ( .A(n_215), .Y(n_1055) );
INVx1_ASAP7_75t_L g834 ( .A(n_217), .Y(n_834) );
INVx1_ASAP7_75t_L g859 ( .A(n_219), .Y(n_859) );
INVx1_ASAP7_75t_L g1041 ( .A(n_220), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g1022 ( .A(n_221), .Y(n_1022) );
INVx2_ASAP7_75t_L g348 ( .A(n_223), .Y(n_348) );
INVx1_ASAP7_75t_L g365 ( .A(n_223), .Y(n_365) );
INVx1_ASAP7_75t_L g400 ( .A(n_223), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_225), .A2(n_233), .B1(n_353), .B2(n_608), .C(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g922 ( .A(n_227), .Y(n_922) );
INVx1_ASAP7_75t_L g673 ( .A(n_228), .Y(n_673) );
AO22x1_ASAP7_75t_L g1122 ( .A1(n_229), .A2(n_242), .B1(n_1085), .B2(n_1088), .Y(n_1122) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_230), .B(n_630), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_232), .Y(n_1027) );
INVx1_ASAP7_75t_L g561 ( .A(n_234), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g1064 ( .A(n_236), .B(n_1065), .Y(n_1064) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_237), .Y(n_481) );
OAI21xp33_ASAP7_75t_SL g705 ( .A1(n_239), .A2(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_239), .Y(n_710) );
INVx1_ASAP7_75t_L g867 ( .A(n_240), .Y(n_867) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_243), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_244), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_245), .A2(n_248), .B1(n_478), .B2(n_977), .C(n_978), .Y(n_976) );
INVx1_ASAP7_75t_L g1024 ( .A(n_246), .Y(n_1024) );
INVx1_ASAP7_75t_L g369 ( .A(n_247), .Y(n_369) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_248), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1069), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1372 ( .A(n_251), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1445 ( .A(n_252), .B(n_255), .Y(n_1445) );
INVx1_ASAP7_75t_L g1447 ( .A(n_252), .Y(n_1447) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1449 ( .A(n_255), .B(n_1447), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g1306 ( .A(n_258), .B(n_1307), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1371 ( .A(n_258), .B(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g335 ( .A(n_259), .B(n_268), .Y(n_335) );
AND2x4_ASAP7_75t_L g341 ( .A(n_259), .B(n_269), .Y(n_341) );
INVx1_ASAP7_75t_L g1301 ( .A(n_260), .Y(n_1301) );
AND2x4_ASAP7_75t_SL g1370 ( .A(n_260), .B(n_1371), .Y(n_1370) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_262), .Y(n_682) );
INVxp67_ASAP7_75t_L g793 ( .A(n_262), .Y(n_793) );
INVx1_ASAP7_75t_L g822 ( .A(n_262), .Y(n_822) );
OR2x6_ASAP7_75t_L g1417 ( .A(n_262), .B(n_1304), .Y(n_1417) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx4f_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
INVx3_ASAP7_75t_L g498 ( .A(n_263), .Y(n_498) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g291 ( .A(n_265), .Y(n_291) );
INVx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
AND2x2_ASAP7_75t_L g299 ( .A(n_265), .B(n_266), .Y(n_299) );
INVx1_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
AND2x2_ASAP7_75t_L g331 ( .A(n_265), .B(n_332), .Y(n_331) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_265), .B(n_266), .Y(n_501) );
OR2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
BUFx2_ASAP7_75t_L g318 ( .A(n_266), .Y(n_318) );
INVx2_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_266), .B(n_295), .Y(n_514) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g1299 ( .A(n_268), .Y(n_1299) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_269), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_269), .B(n_322), .Y(n_1296) );
XNOR2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_701), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
XNOR2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_550), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
XNOR2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_433), .Y(n_277) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_349), .Y(n_281) );
AOI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_325), .B(n_346), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_301), .B(n_304), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_285), .A2(n_510), .B1(n_994), .B2(n_995), .Y(n_993) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx4_ASAP7_75t_L g942 ( .A(n_286), .Y(n_942) );
BUFx6f_ASAP7_75t_L g1400 ( .A(n_286), .Y(n_1400) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g899 ( .A(n_288), .Y(n_899) );
INVx4_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g509 ( .A(n_290), .Y(n_509) );
BUFx3_ASAP7_75t_L g1000 ( .A(n_290), .Y(n_1000) );
INVx2_ASAP7_75t_L g1054 ( .A(n_290), .Y(n_1054) );
AND2x2_ASAP7_75t_L g309 ( .A(n_291), .B(n_310), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_297), .B2(n_300), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
BUFx3_ASAP7_75t_L g569 ( .A(n_294), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_296), .A2(n_390), .B(n_391), .C(n_398), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_297), .A2(n_306), .B(n_311), .C(n_312), .Y(n_305) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
BUFx3_ASAP7_75t_L g567 ( .A(n_298), .Y(n_567) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_298), .Y(n_693) );
BUFx3_ASAP7_75t_L g741 ( .A(n_298), .Y(n_741) );
INVx1_ASAP7_75t_L g818 ( .A(n_298), .Y(n_818) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_298), .B(n_1299), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g585 ( .A(n_299), .Y(n_585) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_302), .B(n_400), .Y(n_539) );
AND2x2_ASAP7_75t_L g544 ( .A(n_302), .B(n_309), .Y(n_544) );
AND2x2_ASAP7_75t_L g547 ( .A(n_302), .B(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_303), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_315), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_307), .Y(n_1333) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_308), .B(n_1283), .Y(n_1282) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g517 ( .A(n_309), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_309), .B(n_314), .Y(n_535) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_314), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_314), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_314), .B(n_348), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_319), .B1(n_320), .B2(n_324), .Y(n_315) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g528 ( .A(n_318), .Y(n_528) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_318), .B(n_1283), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_318), .B(n_1283), .Y(n_1427) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g529 ( .A(n_321), .B(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g575 ( .A(n_321), .B(n_530), .Y(n_575) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_324), .A2(n_369), .B1(n_370), .B2(n_376), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_336), .B1(n_339), .B2(n_342), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g582 ( .A(n_328), .Y(n_582) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g992 ( .A(n_330), .Y(n_992) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_331), .Y(n_548) );
BUFx3_ASAP7_75t_L g695 ( .A(n_331), .Y(n_695) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_331), .B(n_1304), .Y(n_1303) );
AOI222xp33_ASAP7_75t_L g1288 ( .A1(n_333), .A2(n_1289), .B1(n_1290), .B2(n_1291), .C1(n_1293), .C2(n_1294), .Y(n_1288) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g537 ( .A(n_337), .B(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g504 ( .A(n_341), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_341), .B(n_505), .Y(n_894) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g580 ( .A(n_345), .Y(n_580) );
HB1xp67_ASAP7_75t_L g1334 ( .A(n_345), .Y(n_1334) );
INVx1_ASAP7_75t_L g490 ( .A(n_346), .Y(n_490) );
BUFx2_ASAP7_75t_L g777 ( .A(n_346), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_346), .B(n_640), .Y(n_1067) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g430 ( .A(n_347), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g493 ( .A(n_347), .B(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g587 ( .A(n_348), .Y(n_587) );
NAND3xp33_ASAP7_75t_SL g349 ( .A(n_350), .B(n_368), .C(n_383), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_361), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx8_ASAP7_75t_L g390 ( .A(n_354), .Y(n_390) );
INVx3_ASAP7_75t_L g454 ( .A(n_354), .Y(n_454) );
INVx2_ASAP7_75t_L g913 ( .A(n_354), .Y(n_913) );
INVx8_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_355), .B(n_401), .Y(n_623) );
BUFx3_ASAP7_75t_L g651 ( .A(n_355), .Y(n_651) );
AND2x2_ASAP7_75t_L g655 ( .A(n_355), .B(n_656), .Y(n_655) );
BUFx3_ASAP7_75t_L g874 ( .A(n_355), .Y(n_874) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
AND2x4_ASAP7_75t_L g373 ( .A(n_356), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_357), .B(n_381), .Y(n_388) );
OR2x2_ASAP7_75t_L g411 ( .A(n_357), .B(n_359), .Y(n_411) );
AND2x4_ASAP7_75t_L g447 ( .A(n_357), .B(n_396), .Y(n_447) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g375 ( .A(n_362), .Y(n_375) );
OR2x2_ASAP7_75t_L g377 ( .A(n_362), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g385 ( .A(n_362), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .Y(n_362) );
OR2x2_ASAP7_75t_L g407 ( .A(n_363), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g506 ( .A(n_363), .Y(n_506) );
HB1xp67_ASAP7_75t_L g1369 ( .A(n_363), .Y(n_1369) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g530 ( .A(n_364), .Y(n_530) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g440 ( .A(n_366), .Y(n_440) );
INVx1_ASAP7_75t_L g656 ( .A(n_366), .Y(n_656) );
INVx3_ASAP7_75t_L g402 ( .A(n_367), .Y(n_402) );
NAND2xp33_ASAP7_75t_SL g408 ( .A(n_367), .B(n_404), .Y(n_408) );
BUFx3_ASAP7_75t_L g488 ( .A(n_367), .Y(n_488) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVx2_ASAP7_75t_L g424 ( .A(n_371), .Y(n_424) );
INVx2_ASAP7_75t_L g833 ( .A(n_371), .Y(n_833) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_SL g637 ( .A(n_372), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_373), .Y(n_485) );
BUFx8_ASAP7_75t_L g612 ( .A(n_373), .Y(n_612) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_378), .Y(n_414) );
INVx4_ASAP7_75t_L g468 ( .A(n_378), .Y(n_468) );
INVx3_ASAP7_75t_L g766 ( .A(n_378), .Y(n_766) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_378), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g397 ( .A(n_379), .Y(n_397) );
BUFx2_ASAP7_75t_L g599 ( .A(n_379), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_380), .Y(n_1347) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g396 ( .A(n_381), .Y(n_396) );
INVx2_ASAP7_75t_L g392 ( .A(n_382), .Y(n_392) );
AND2x4_ASAP7_75t_L g443 ( .A(n_382), .B(n_395), .Y(n_443) );
BUFx2_ASAP7_75t_L g1344 ( .A(n_382), .Y(n_1344) );
NOR2xp33_ASAP7_75t_SL g383 ( .A(n_384), .B(n_405), .Y(n_383) );
INVx1_ASAP7_75t_L g731 ( .A(n_386), .Y(n_731) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_387), .Y(n_617) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g421 ( .A(n_388), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_390), .A2(n_964), .B1(n_1016), .B2(n_1022), .Y(n_1021) );
INVx3_ASAP7_75t_L g596 ( .A(n_392), .Y(n_596) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g593 ( .A(n_394), .B(n_401), .Y(n_593) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_410), .B1(n_428), .B2(n_429), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g914 ( .A1(n_397), .A2(n_451), .B1(n_487), .B2(n_915), .C(n_916), .Y(n_914) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_397), .A2(n_410), .B1(n_471), .B2(n_921), .C(n_922), .Y(n_920) );
INVx2_ASAP7_75t_L g1037 ( .A(n_397), .Y(n_1037) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
OR2x2_ASAP7_75t_L g534 ( .A(n_399), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g689 ( .A(n_399), .Y(n_689) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g1325 ( .A(n_400), .Y(n_1325) );
INVx1_ASAP7_75t_L g457 ( .A(n_401), .Y(n_457) );
AND2x6_ASAP7_75t_L g595 ( .A(n_401), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_402), .B(n_432), .Y(n_431) );
NAND3x1_ASAP7_75t_L g1324 ( .A(n_402), .B(n_432), .C(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1354 ( .A(n_402), .Y(n_1354) );
OR2x6_ASAP7_75t_L g1356 ( .A(n_402), .B(n_421), .Y(n_1356) );
AND2x4_ASAP7_75t_L g1358 ( .A(n_402), .B(n_447), .Y(n_1358) );
OR2x4_ASAP7_75t_L g1362 ( .A(n_402), .B(n_411), .Y(n_1362) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g487 ( .A(n_404), .B(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_404), .Y(n_1367) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .A3(n_415), .B1(n_423), .B2(n_427), .B3(n_430), .Y(n_405) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_406), .Y(n_1317) );
BUFx4f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx8_ASAP7_75t_L g1379 ( .A(n_407), .Y(n_1379) );
BUFx2_ASAP7_75t_L g606 ( .A(n_408), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g1040 ( .A(n_410), .Y(n_1040) );
BUFx4f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
BUFx3_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
INVx2_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
OR2x4_ASAP7_75t_L g1353 ( .A(n_411), .B(n_1354), .Y(n_1353) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_414), .A2(n_487), .B1(n_611), .B2(n_718), .C(n_719), .Y(n_717) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_414), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_419), .B2(n_422), .Y(n_415) );
INVx8_ASAP7_75t_L g605 ( .A(n_417), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_417), .A2(n_867), .B1(n_868), .B2(n_869), .C(n_870), .Y(n_866) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g451 ( .A(n_418), .Y(n_451) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
INVx2_ASAP7_75t_SL g968 ( .A(n_418), .Y(n_968) );
INVx3_ASAP7_75t_L g977 ( .A(n_418), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_419), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g1388 ( .A1(n_424), .A2(n_464), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
INVx3_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
NAND4xp75_ASAP7_75t_L g434 ( .A(n_435), .B(n_491), .C(n_531), .D(n_541), .Y(n_434) );
OAI21x1_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_458), .B(n_489), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_441), .B(n_452), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_438), .A2(n_560), .B1(n_614), .B2(n_620), .Y(n_613) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g975 ( .A(n_439), .Y(n_975) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g638 ( .A(n_440), .Y(n_638) );
AND2x4_ASAP7_75t_L g640 ( .A(n_440), .B(n_443), .Y(n_640) );
AOI221xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_444), .B1(n_445), .B2(n_448), .C(n_449), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx12f_ASAP7_75t_L g602 ( .A(n_443), .Y(n_602) );
INVx5_ASAP7_75t_L g648 ( .A(n_443), .Y(n_648) );
BUFx2_ASAP7_75t_L g962 ( .A(n_443), .Y(n_962) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g836 ( .A(n_446), .Y(n_836) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g604 ( .A(n_447), .Y(n_604) );
BUFx2_ASAP7_75t_L g619 ( .A(n_447), .Y(n_619) );
AND2x2_ASAP7_75t_L g658 ( .A(n_447), .B(n_656), .Y(n_658) );
BUFx2_ASAP7_75t_L g871 ( .A(n_447), .Y(n_871) );
BUFx2_ASAP7_75t_L g964 ( .A(n_447), .Y(n_964) );
BUFx2_ASAP7_75t_L g981 ( .A(n_447), .Y(n_981) );
BUFx2_ASAP7_75t_L g1350 ( .A(n_447), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_450), .A2(n_471), .B1(n_482), .B2(n_725), .C(n_726), .Y(n_724) );
INVx2_ASAP7_75t_L g965 ( .A(n_451), .Y(n_965) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_455), .C(n_456), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_454), .A2(n_556), .B1(n_576), .B2(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x6_ASAP7_75t_L g598 ( .A(n_457), .B(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_465), .B1(n_472), .B2(n_480), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_463), .B2(n_464), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_460), .A2(n_473), .B1(n_497), .B2(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_463), .A2(n_481), .B1(n_508), .B2(n_510), .C(n_515), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_464), .A2(n_1314), .B1(n_1315), .B2(n_1316), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_469), .B2(n_470), .C(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g482 ( .A(n_468), .Y(n_482) );
INVx2_ASAP7_75t_L g646 ( .A(n_468), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_469), .A2(n_471), .B1(n_765), .B2(n_774), .C(n_775), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g1310 ( .A1(n_469), .A2(n_1036), .B1(n_1311), .B2(n_1312), .Y(n_1310) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_469), .A2(n_1319), .B1(n_1320), .B2(n_1321), .Y(n_1318) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_469), .A2(n_1036), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_469), .A2(n_1393), .B1(n_1394), .B2(n_1395), .Y(n_1392) );
INVx3_ASAP7_75t_L g608 ( .A(n_471), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_471), .B(n_664), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_471), .A2(n_1036), .B1(n_1038), .B2(n_1039), .C(n_1041), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_477), .B2(n_478), .Y(n_472) );
BUFx4f_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_475), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_720) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_483), .B2(n_486), .C(n_487), .Y(n_480) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g615 ( .A(n_485), .Y(n_615) );
INVx1_ASAP7_75t_L g644 ( .A(n_485), .Y(n_644) );
INVx2_ASAP7_75t_L g1315 ( .A(n_485), .Y(n_1315) );
AND2x4_ASAP7_75t_L g1364 ( .A(n_485), .B(n_1354), .Y(n_1364) );
BUFx6f_ASAP7_75t_L g1386 ( .A(n_485), .Y(n_1386) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_487), .A2(n_648), .B1(n_649), .B2(n_650), .C(n_652), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_487), .A2(n_765), .B1(n_767), .B2(n_768), .C(n_769), .Y(n_764) );
INVx3_ASAP7_75t_L g1343 ( .A(n_488), .Y(n_1343) );
OAI31xp33_ASAP7_75t_L g829 ( .A1(n_489), .A2(n_830), .A3(n_831), .B(n_845), .Y(n_829) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI211x1_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B(n_502), .C(n_523), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_492), .A2(n_504), .B1(n_688), .B2(n_788), .C1(n_795), .C2(n_799), .Y(n_787) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI31xp33_ASAP7_75t_L g565 ( .A1(n_493), .A2(n_566), .A3(n_568), .B(n_570), .Y(n_565) );
INVx2_ASAP7_75t_L g686 ( .A(n_493), .Y(n_686) );
INVx4_ASAP7_75t_L g744 ( .A(n_493), .Y(n_744) );
INVx2_ASAP7_75t_L g815 ( .A(n_493), .Y(n_815) );
AOI222xp33_ASAP7_75t_L g934 ( .A1(n_493), .A2(n_504), .B1(n_688), .B2(n_935), .C1(n_936), .C2(n_943), .Y(n_934) );
INVx1_ASAP7_75t_L g1397 ( .A(n_493), .Y(n_1397) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g697 ( .A(n_498), .Y(n_697) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g540 ( .A(n_500), .B(n_539), .Y(n_540) );
OR2x2_ASAP7_75t_L g563 ( .A(n_500), .B(n_539), .Y(n_563) );
INVx2_ASAP7_75t_SL g1406 ( .A(n_500), .Y(n_1406) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_501), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_507), .B(n_518), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_503), .A2(n_814), .B1(n_1330), .B2(n_1335), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_504), .B(n_578), .C(n_581), .Y(n_577) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_504), .A2(n_677), .A3(n_680), .B1(n_685), .B2(n_687), .C1(n_688), .C2(n_691), .Y(n_676) );
AOI332xp33_ASAP7_75t_L g739 ( .A1(n_504), .A2(n_688), .A3(n_740), .B1(n_742), .B2(n_743), .B3(n_745), .C1(n_746), .C2(n_748), .Y(n_739) );
AOI322xp5_ASAP7_75t_L g810 ( .A1(n_504), .A2(n_562), .A3(n_811), .B1(n_812), .B2(n_813), .C1(n_816), .C2(n_825), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g990 ( .A1(n_504), .A2(n_991), .B(n_996), .C(n_1004), .Y(n_990) );
INVx2_ASAP7_75t_L g1407 ( .A(n_504), .Y(n_1407) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_510), .A2(n_1381), .B1(n_1393), .B2(n_1399), .Y(n_1398) );
INVx6_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g684 ( .A(n_511), .Y(n_684) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g699 ( .A(n_512), .Y(n_699) );
INVx4_ASAP7_75t_L g824 ( .A(n_512), .Y(n_824) );
INVx2_ASAP7_75t_SL g948 ( .A(n_512), .Y(n_948) );
INVx1_ASAP7_75t_L g1410 ( .A(n_512), .Y(n_1410) );
INVx8_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g794 ( .A(n_513), .Y(n_794) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_513), .B(n_1283), .Y(n_1287) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g747 ( .A(n_517), .Y(n_747) );
INVx2_ASAP7_75t_L g1058 ( .A(n_517), .Y(n_1058) );
INVx2_ASAP7_75t_L g1337 ( .A(n_517), .Y(n_1337) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_518), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_518), .A2(n_897), .B(n_898), .Y(n_896) );
OAI21xp5_ASAP7_75t_L g996 ( .A1(n_518), .A2(n_814), .B(n_997), .Y(n_996) );
OAI21xp5_ASAP7_75t_SL g1049 ( .A1(n_518), .A2(n_1050), .B(n_1052), .Y(n_1049) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx4_ASAP7_75t_L g902 ( .A(n_519), .Y(n_902) );
BUFx4f_ASAP7_75t_L g1056 ( .A(n_519), .Y(n_1056) );
BUFx4f_ASAP7_75t_L g1061 ( .A(n_519), .Y(n_1061) );
BUFx4f_ASAP7_75t_L g1425 ( .A(n_519), .Y(n_1425) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2x2_ASAP7_75t_L g526 ( .A(n_521), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_526), .Y(n_786) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g543 ( .A(n_530), .Y(n_543) );
INVxp67_ASAP7_75t_L g1014 ( .A(n_530), .Y(n_1014) );
INVx1_ASAP7_75t_L g1307 ( .A(n_530), .Y(n_1307) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_534), .B(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g690 ( .A(n_535), .Y(n_690) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_537), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_537), .A2(n_737), .B(n_738), .Y(n_736) );
AOI211xp5_ASAP7_75t_L g783 ( .A1(n_537), .A2(n_756), .B(n_784), .C(n_785), .Y(n_783) );
AOI222xp33_ASAP7_75t_L g806 ( .A1(n_537), .A2(n_572), .B1(n_574), .B2(n_807), .C1(n_808), .C2(n_809), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g884 ( .A1(n_537), .A2(n_562), .B1(n_688), .B2(n_861), .C1(n_864), .C2(n_885), .Y(n_884) );
AOI222xp33_ASAP7_75t_L g931 ( .A1(n_537), .A2(n_572), .B1(n_574), .B2(n_924), .C1(n_932), .C2(n_933), .Y(n_931) );
INVxp67_ASAP7_75t_L g986 ( .A(n_537), .Y(n_986) );
INVx1_ASAP7_75t_L g1015 ( .A(n_537), .Y(n_1015) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_545), .B1(n_546), .B2(n_549), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_542), .B(n_556), .Y(n_555) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_542), .A2(n_670), .B(n_671), .C(n_675), .Y(n_669) );
INVx3_ASAP7_75t_L g706 ( .A(n_542), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_542), .B(n_801), .Y(n_800) );
AOI211x1_ASAP7_75t_L g803 ( .A1(n_542), .A2(n_804), .B(n_805), .C(n_828), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_542), .A2(n_780), .B1(n_859), .B2(n_882), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_542), .B(n_950), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_542), .A2(n_546), .B1(n_1011), .B2(n_1012), .C1(n_1016), .C2(n_1017), .Y(n_1010) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x4_ASAP7_75t_L g546 ( .A(n_543), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g625 ( .A(n_546), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_546), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_546), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g781 ( .A(n_546), .Y(n_781) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_546), .Y(n_989) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_548), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_628), .B1(n_629), .B2(n_700), .Y(n_550) );
INVx1_ASAP7_75t_L g700 ( .A(n_551), .Y(n_700) );
OAI21x1_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_553), .B(n_627), .Y(n_551) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_552), .B(n_555), .C(n_557), .D(n_586), .Y(n_627) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .C(n_586), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_562), .A2(n_570), .B(n_715), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_562), .A2(n_570), .B(n_952), .Y(n_951) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_565), .B(n_571), .C(n_577), .Y(n_564) );
AOI21xp33_ASAP7_75t_L g826 ( .A1(n_570), .A2(n_688), .B(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_573), .B1(n_574), .B2(n_576), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_572), .A2(n_574), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_572), .A2(n_574), .B1(n_1022), .B2(n_1024), .Y(n_1063) );
INVx2_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g789 ( .A(n_584), .Y(n_789) );
INVx1_ASAP7_75t_L g892 ( .A(n_584), .Y(n_892) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B1(n_624), .B2(n_626), .Y(n_586) );
INVx2_ASAP7_75t_SL g665 ( .A(n_587), .Y(n_665) );
OAI31xp33_ASAP7_75t_SL g707 ( .A1(n_587), .A2(n_708), .A3(n_712), .B(n_716), .Y(n_707) );
INVx1_ASAP7_75t_L g1047 ( .A(n_587), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .C(n_613), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_597), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g635 ( .A(n_593), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_593), .A2(n_595), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_593), .A2(n_595), .B1(n_808), .B2(n_825), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_593), .A2(n_595), .B1(n_597), .B2(n_863), .C(n_864), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_593), .A2(n_595), .B1(n_597), .B2(n_971), .C(n_972), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_593), .A2(n_595), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
INVx4_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g840 ( .A(n_599), .Y(n_840) );
INVx1_ASAP7_75t_L g1438 ( .A(n_599), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B1(n_607), .B2(n_609), .Y(n_600) );
BUFx2_ASAP7_75t_L g763 ( .A(n_602), .Y(n_763) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_611), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g768 ( .A(n_612), .Y(n_768) );
INVx2_ASAP7_75t_SL g919 ( .A(n_612), .Y(n_919) );
INVx3_ASAP7_75t_L g1031 ( .A(n_612), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_616), .A2(n_823), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_616), .A2(n_768), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_616), .A2(n_1384), .B1(n_1385), .B2(n_1387), .Y(n_1383) );
CKINVDCx8_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g723 ( .A(n_617), .Y(n_723) );
INVx3_ASAP7_75t_L g868 ( .A(n_617), .Y(n_868) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI211xp5_ASAP7_75t_SL g632 ( .A1(n_622), .A2(n_633), .B(n_634), .C(n_636), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g755 ( .A1(n_622), .A2(n_756), .B(n_757), .C(n_758), .Y(n_755) );
AOI211xp5_ASAP7_75t_SL g923 ( .A1(n_622), .A2(n_924), .B(n_925), .C(n_926), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_622), .A2(n_974), .B1(n_976), .B2(n_982), .Y(n_973) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_623), .B(n_1014), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_624), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_668), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_641), .B(n_665), .C(n_666), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_637), .Y(n_860) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_640), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_858) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_642), .B(n_653), .C(n_659), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_644), .A2(n_868), .B1(n_1327), .B2(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_R g772 ( .A(n_648), .Y(n_772) );
INVx1_ASAP7_75t_L g1033 ( .A(n_648), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_649), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g762 ( .A(n_650), .Y(n_762) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
BUFx3_ASAP7_75t_L g843 ( .A(n_651), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_652), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_655), .A2(n_658), .B1(n_710), .B2(n_711), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_655), .A2(n_658), .B1(n_804), .B2(n_809), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_655), .A2(n_658), .B1(n_882), .B2(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_676), .Y(n_668) );
BUFx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_682), .A2(n_794), .B1(n_797), .B2(n_798), .Y(n_796) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g891 ( .A(n_695), .Y(n_891) );
INVx1_ASAP7_75t_L g939 ( .A(n_695), .Y(n_939) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_850), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_750), .B1(n_848), .B2(n_849), .Y(n_702) );
INVx1_ASAP7_75t_L g849 ( .A(n_703), .Y(n_849) );
XOR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_749), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_732), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .B1(n_724), .B2(n_727), .Y(n_716) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND4xp25_ASAP7_75t_SL g732 ( .A(n_733), .B(n_734), .C(n_736), .D(n_739), .Y(n_732) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_743), .Y(n_1051) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g848 ( .A(n_750), .Y(n_848) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
XOR2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_802), .Y(n_751) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_782), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_SL g754 ( .A1(n_755), .A2(n_759), .B(n_776), .C(n_778), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_770), .C(n_771), .Y(n_759) );
BUFx2_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g877 ( .A(n_766), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g790 ( .A1(n_775), .A2(n_791), .B1(n_792), .B2(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_777), .A2(n_857), .B(n_865), .Y(n_856) );
INVx2_ASAP7_75t_L g927 ( .A(n_777), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_777), .A2(n_959), .B(n_983), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .C(n_800), .Y(n_782) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
XOR2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_847), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .C(n_826), .Y(n_805) );
INVx1_ASAP7_75t_L g897 ( .A(n_813), .Y(n_897) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g937 ( .A(n_818), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_821), .B1(n_823), .B2(n_824), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g946 ( .A(n_822), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_824), .A2(n_922), .B1(n_941), .B2(n_942), .Y(n_940) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_837), .C(n_844), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B(n_841), .C(n_842), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_953), .B2(n_954), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
XOR2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_907), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g905 ( .A(n_855), .Y(n_905) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_856), .B(n_884), .C(n_886), .D(n_904), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_875), .C(n_881), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_867), .A2(n_899), .B1(n_900), .B2(n_901), .C(n_903), .Y(n_898) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx2_ASAP7_75t_L g880 ( .A(n_874), .Y(n_880) );
OAI211xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_877), .B(n_878), .C(n_879), .Y(n_875) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_877), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_896), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_893), .C(n_895), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
OAI221xp5_ASAP7_75t_L g1060 ( .A1(n_899), .A2(n_1027), .B1(n_1038), .B2(n_1061), .C(n_1062), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_901), .A2(n_998), .B1(n_1001), .B2(n_1002), .C(n_1003), .Y(n_997) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OR2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_930), .Y(n_908) );
A2O1A1Ixp33_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_923), .B(n_927), .C(n_928), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .C(n_917), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_913), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND4xp25_ASAP7_75t_L g930 ( .A(n_931), .B(n_934), .C(n_949), .D(n_951), .Y(n_930) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_944) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_955), .Y(n_954) );
XNOR2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_1007), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_1005), .B(n_1006), .Y(n_956) );
AND3x1_ASAP7_75t_L g957 ( .A(n_958), .B(n_984), .C(n_990), .Y(n_957) );
AOI31xp33_ASAP7_75t_L g1006 ( .A1(n_958), .A2(n_984), .A3(n_990), .B(n_1005), .Y(n_1006) );
NAND3xp33_ASAP7_75t_SL g959 ( .A(n_960), .B(n_970), .C(n_973), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_963), .B1(n_966), .B2(n_969), .Y(n_960) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_974), .Y(n_1020) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AND2x2_ASAP7_75t_L g984 ( .A(n_985), .B(n_987), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .Y(n_987) );
INVx3_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1018), .C(n_1048), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1015), .Y(n_1012) );
OAI21xp33_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1034), .B(n_1045), .Y(n_1018) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B(n_1023), .C(n_1026), .Y(n_1019) );
OAI211xp5_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B(n_1029), .C(n_1032), .Y(n_1026) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_1043), .A2(n_1053), .B1(n_1055), .B2(n_1056), .C(n_1057), .Y(n_1052) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
NOR3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1059), .C(n_1064), .Y(n_1048) );
INVxp67_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_1053), .A2(n_1056), .B1(n_1384), .B2(n_1389), .Y(n_1401) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1053), .Y(n_1404) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx2_ASAP7_75t_L g1331 ( .A(n_1054), .Y(n_1331) );
OAI221xp5_ASAP7_75t_SL g1330 ( .A1(n_1056), .A2(n_1314), .B1(n_1327), .B2(n_1331), .C(n_1332), .Y(n_1330) );
OAI221xp5_ASAP7_75t_SL g1335 ( .A1(n_1056), .A2(n_1312), .B1(n_1320), .B2(n_1331), .C(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI21xp33_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1270), .B(n_1274), .Y(n_1069) );
NOR2xp67_ASAP7_75t_SL g1070 ( .A(n_1071), .B(n_1221), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1168), .B(n_1176), .Y(n_1071) );
NOR4xp25_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1135), .C(n_1147), .D(n_1163), .Y(n_1072) );
OAI211xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1090), .B(n_1108), .C(n_1123), .Y(n_1073) );
CKINVDCx14_ASAP7_75t_R g1074 ( .A(n_1075), .Y(n_1074) );
OAI322xp33_ASAP7_75t_L g1147 ( .A1(n_1075), .A2(n_1092), .A3(n_1148), .B1(n_1149), .B2(n_1154), .C1(n_1159), .C2(n_1161), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_1075), .A2(n_1101), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
INVx3_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1076), .B(n_1118), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1076), .B(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1076), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1076), .B(n_1137), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1076), .B(n_1129), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1076), .B(n_1119), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1076), .B(n_1118), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1076), .B(n_1129), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1076), .B(n_1119), .Y(n_1260) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1084), .Y(n_1076) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1078), .Y(n_1173) );
AND2x6_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1080), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1079), .B(n_1083), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_1079), .B(n_1086), .Y(n_1085) );
AND2x6_ASAP7_75t_L g1088 ( .A(n_1079), .B(n_1089), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1079), .B(n_1083), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1079), .B(n_1083), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1081), .B(n_1087), .Y(n_1086) );
INVxp67_ASAP7_75t_L g1175 ( .A(n_1082), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1273 ( .A(n_1082), .Y(n_1273) );
OAI21xp5_ASAP7_75t_L g1446 ( .A1(n_1083), .A2(n_1447), .B(n_1448), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1096), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1091), .B(n_1105), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1091), .B(n_1144), .Y(n_1143) );
AND3x1_ASAP7_75t_L g1196 ( .A(n_1091), .B(n_1105), .C(n_1115), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1091), .B(n_1115), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1091), .B(n_1097), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1091), .B(n_1235), .Y(n_1234) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_1092), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1092), .B(n_1144), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1092), .B(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1092), .B(n_1101), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1092), .B(n_1235), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1101), .Y(n_1096) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1097), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1097), .B(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1097), .B(n_1144), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1097), .B(n_1152), .Y(n_1230) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1098), .B(n_1110), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1098), .B(n_1129), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1098), .B(n_1129), .Y(n_1137) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1098), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1098), .B(n_1119), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1098), .B(n_1113), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1098), .B(n_1128), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1098), .B(n_1138), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1098), .B(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1100), .Y(n_1098) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1101), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1101), .B(n_1214), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .Y(n_1101) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1102), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1102), .B(n_1145), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1102), .B(n_1113), .Y(n_1262) );
NAND3xp33_ASAP7_75t_L g1263 ( .A(n_1102), .B(n_1170), .C(n_1225), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1105), .B(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1105), .Y(n_1145) );
OAI211xp5_ASAP7_75t_L g1187 ( .A1(n_1105), .A2(n_1133), .B(n_1188), .C(n_1192), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_1105), .B(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1112), .B(n_1116), .Y(n_1108) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1111), .B(n_1126), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1242 ( .A1(n_1111), .A2(n_1166), .B1(n_1197), .B2(n_1243), .C(n_1244), .Y(n_1242) );
AOI21xp33_ASAP7_75t_L g1247 ( .A1(n_1111), .A2(n_1133), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1112), .B(n_1142), .Y(n_1182) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1112), .B(n_1143), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1113), .B(n_1115), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1113), .B(n_1115), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1114), .B(n_1144), .Y(n_1148) );
NAND3xp33_ASAP7_75t_L g1154 ( .A(n_1114), .B(n_1155), .C(n_1158), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1114), .B(n_1214), .Y(n_1213) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_1115), .A2(n_1143), .B1(n_1184), .B2(n_1185), .C(n_1187), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1115), .B(n_1145), .Y(n_1235) );
AOI21xp5_ASAP7_75t_L g1244 ( .A1(n_1116), .A2(n_1245), .B(n_1247), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1116), .B(n_1182), .Y(n_1249) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_1118), .B(n_1133), .Y(n_1132) );
NOR2xp33_ASAP7_75t_SL g1150 ( .A(n_1118), .B(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1118), .B(n_1128), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1118), .B(n_1170), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1118), .B(n_1190), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1118), .B(n_1152), .Y(n_1254) );
CKINVDCx6p67_ASAP7_75t_R g1118 ( .A(n_1119), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_1119), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1119), .B(n_1165), .Y(n_1164) );
OR2x6_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1122), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1120), .B(n_1122), .Y(n_1158) );
OAI21xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1132), .B(n_1134), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
CKINVDCx6p67_ASAP7_75t_R g1165 ( .A(n_1127), .Y(n_1165) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1128), .Y(n_1157) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1129), .B(n_1153), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1131), .Y(n_1129) );
CKINVDCx14_ASAP7_75t_R g1210 ( .A(n_1134), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1134), .B(n_1230), .Y(n_1229) );
O2A1O1Ixp33_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1138), .B(n_1139), .C(n_1146), .Y(n_1135) );
AOI21xp33_ASAP7_75t_L g1267 ( .A1(n_1136), .A2(n_1268), .B(n_1269), .Y(n_1267) );
CKINVDCx14_ASAP7_75t_R g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1143), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1141), .B(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1141), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1141), .B(n_1190), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1141), .B(n_1234), .Y(n_1233) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1143), .B(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1143), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1144), .B(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1144), .Y(n_1248) );
O2A1O1Ixp33_ASAP7_75t_L g1238 ( .A1(n_1146), .A2(n_1159), .B(n_1239), .C(n_1241), .Y(n_1238) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
AOI21xp33_ASAP7_75t_L g1231 ( .A1(n_1151), .A2(n_1232), .B(n_1233), .Y(n_1231) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1152), .B(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1155), .B(n_1160), .Y(n_1266) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1157), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1157), .B(n_1160), .Y(n_1237) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI21xp5_ASAP7_75t_SL g1202 ( .A1(n_1160), .A2(n_1203), .B(n_1205), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_1161), .A2(n_1165), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1165), .A2(n_1260), .B1(n_1261), .B2(n_1263), .Y(n_1259) );
OAI31xp33_ASAP7_75t_SL g1236 ( .A1(n_1168), .A2(n_1237), .A3(n_1238), .B(n_1242), .Y(n_1236) );
INVx3_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
INVx2_ASAP7_75t_SL g1169 ( .A(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_1170), .Y(n_1211) );
OAI22xp5_ASAP7_75t_SL g1171 ( .A1(n_1172), .A2(n_1173), .B1(n_1174), .B2(n_1175), .Y(n_1171) );
XOR2x2_ASAP7_75t_L g1276 ( .A(n_1174), .B(n_1277), .Y(n_1276) );
AOI211xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1179), .B(n_1193), .C(n_1208), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OAI21xp5_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1181), .B(n_1183), .Y(n_1179) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1180), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1180), .B(n_1198), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1180), .B(n_1218), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVxp67_ASAP7_75t_SL g1209 ( .A(n_1184), .Y(n_1209) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
OAI321xp33_ASAP7_75t_L g1208 ( .A1(n_1191), .A2(n_1209), .A3(n_1210), .B1(n_1211), .B2(n_1212), .C(n_1215), .Y(n_1208) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1197), .B1(n_1199), .B2(n_1201), .C(n_1202), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1198), .B(n_1225), .Y(n_1243) );
OAI21xp5_ASAP7_75t_L g1264 ( .A1(n_1198), .A2(n_1265), .B(n_1267), .Y(n_1264) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVxp67_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1217), .Y(n_1215) );
AOI211xp5_ASAP7_75t_L g1222 ( .A1(n_1216), .A2(n_1223), .B(n_1226), .C(n_1231), .Y(n_1222) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1216), .Y(n_1232) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND5xp2_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1236), .C(n_1249), .D(n_1250), .E(n_1264), .Y(n_1221) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
OAI21xp5_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1228), .B(n_1229), .Y(n_1226) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1234), .Y(n_1241) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
NOR3xp33_ASAP7_75t_SL g1250 ( .A(n_1251), .B(n_1255), .C(n_1259), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .Y(n_1252) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1253), .Y(n_1269) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVxp67_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
CKINVDCx20_ASAP7_75t_R g1270 ( .A(n_1271), .Y(n_1270) );
CKINVDCx20_ASAP7_75t_R g1271 ( .A(n_1272), .Y(n_1271) );
INVx4_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
HB1xp67_ASAP7_75t_SL g1275 ( .A(n_1276), .Y(n_1275) );
NAND3x1_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1308), .C(n_1338), .Y(n_1277) );
OAI21xp5_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1300), .B(n_1305), .Y(n_1278) );
NAND3xp33_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1288), .C(n_1297), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1282), .B1(n_1284), .B2(n_1285), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_1281), .A2(n_1284), .B1(n_1352), .B2(n_1355), .Y(n_1351) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_1286), .Y(n_1285) );
BUFx2_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1287), .Y(n_1421) );
AOI222xp33_ASAP7_75t_L g1340 ( .A1(n_1289), .A2(n_1290), .B1(n_1293), .B2(n_1341), .C1(n_1345), .C2(n_1348), .Y(n_1340) );
BUFx3_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1295), .Y(n_1429) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx3_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx3_ASAP7_75t_SL g1302 ( .A(n_1303), .Y(n_1302) );
INVx4_ASAP7_75t_L g1413 ( .A(n_1303), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
BUFx3_ASAP7_75t_L g1431 ( .A(n_1306), .Y(n_1431) );
NOR2x1_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1329), .Y(n_1308) );
OAI33xp33_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1313), .A3(n_1317), .B1(n_1318), .B2(n_1322), .B3(n_1326), .Y(n_1309) );
CKINVDCx5p33_ASAP7_75t_R g1322 ( .A(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1323), .Y(n_1391) );
INVx3_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI21xp33_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1359), .B(n_1365), .Y(n_1338) );
NAND3xp33_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1351), .C(n_1357), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_1341), .A2(n_1345), .B1(n_1428), .B2(n_1440), .Y(n_1439) );
BUFx3_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1344), .Y(n_1342) );
AND2x4_ASAP7_75t_L g1346 ( .A(n_1343), .B(n_1347), .Y(n_1346) );
BUFx6f_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_SL g1352 ( .A(n_1353), .Y(n_1352) );
BUFx2_ASAP7_75t_L g1442 ( .A(n_1353), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1355), .Y(n_1443) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
CKINVDCx8_ASAP7_75t_R g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx2_ASAP7_75t_SL g1435 ( .A(n_1362), .Y(n_1435) );
INVx2_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OAI31xp33_ASAP7_75t_L g1432 ( .A1(n_1365), .A2(n_1433), .A3(n_1436), .B(n_1441), .Y(n_1432) );
AND2x2_ASAP7_75t_SL g1365 ( .A(n_1366), .B(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_SL g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVxp67_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
AND3x1_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1411), .C(n_1432), .Y(n_1376) );
NOR2xp33_ASAP7_75t_SL g1377 ( .A(n_1378), .B(n_1396), .Y(n_1377) );
OAI33xp33_ASAP7_75t_L g1378 ( .A1(n_1379), .A2(n_1380), .A3(n_1383), .B1(n_1388), .B2(n_1391), .B3(n_1392), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1382), .A2(n_1395), .B1(n_1403), .B2(n_1405), .Y(n_1402) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_1387), .A2(n_1390), .B1(n_1399), .B2(n_1409), .Y(n_1408) );
OAI33xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1398), .A3(n_1401), .B1(n_1402), .B2(n_1407), .B3(n_1408), .Y(n_1396) );
INVx2_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx5_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
BUFx3_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
OAI31xp33_ASAP7_75t_L g1411 ( .A1(n_1412), .A2(n_1414), .A3(n_1422), .B(n_1431), .Y(n_1411) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx2_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx2_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1428), .B1(n_1429), .B2(n_1430), .Y(n_1426) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVxp67_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
HB1xp67_ASAP7_75t_SL g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
endmodule