module fake_ibex_491_n_1051 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1051);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1051;

wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_580;
wire n_483;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_200;
wire n_564;
wire n_506;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_1033;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_947;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_890;
wire n_874;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_202;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_67),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_150),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_171),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_107),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_130),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_57),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_40),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_21),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_38),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_52),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_27),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_17),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_45),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_152),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_116),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_20),
.B(n_14),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_92),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_71),
.B(n_17),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_72),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_42),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_76),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_159),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_185),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_112),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_74),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_73),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_91),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_79),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_58),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_125),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_114),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_4),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_62),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_170),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_160),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_109),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_127),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_102),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_33),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_65),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_161),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_84),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_86),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_53),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_184),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_68),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_69),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_88),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_75),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_98),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_131),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_138),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_135),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_81),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_165),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_77),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_153),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_136),
.B(n_101),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_15),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_167),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_80),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_28),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_35),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_103),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_2),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_32),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_99),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_16),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_27),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_113),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_143),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_154),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_15),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_14),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_221),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_200),
.B(n_0),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_247),
.B(n_0),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_200),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_231),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_199),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_1),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g340 ( 
.A(n_264),
.B(n_2),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_221),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_275),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_201),
.A2(n_106),
.B(n_196),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_221),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_223),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_203),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_287),
.B(n_3),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_256),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_223),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_206),
.Y(n_358)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_227),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_213),
.B(n_7),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_239),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_209),
.A2(n_110),
.B(n_192),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_268),
.B(n_9),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_257),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_214),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_257),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_257),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_216),
.A2(n_108),
.B(n_190),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_267),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_254),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_219),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_246),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g380 ( 
.A1(n_265),
.A2(n_104),
.B(n_188),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_285),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_298),
.B(n_11),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_228),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_232),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_266),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_267),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_282),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_235),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_237),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_204),
.B(n_12),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_290),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_282),
.Y(n_396)
);

BUFx8_ASAP7_75t_L g397 ( 
.A(n_282),
.Y(n_397)
);

CKINVDCx8_ASAP7_75t_R g398 ( 
.A(n_269),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_280),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_282),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_299),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_335),
.B(n_299),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_238),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_295),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_326),
.B(n_229),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_236),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_357),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

AO21x2_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_242),
.B(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

BUFx6f_ASAP7_75t_SL g433 ( 
.A(n_352),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_338),
.B(n_250),
.Y(n_436)
);

AOI21x1_ASAP7_75t_L g437 ( 
.A1(n_380),
.A2(n_258),
.B(n_244),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_328),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_272),
.Y(n_439)
);

CKINVDCx6p67_ASAP7_75t_R g440 ( 
.A(n_343),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_338),
.B(n_319),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_338),
.B(n_319),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_350),
.B(n_207),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_328),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_327),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_210),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_328),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_333),
.A2(n_262),
.B(n_259),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_336),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_374),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_328),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_336),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_328),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_332),
.B(n_311),
.C(n_283),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_339),
.B(n_314),
.C(n_245),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_337),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_343),
.B(n_312),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_336),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_330),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

BUFx6f_ASAP7_75t_SL g473 ( 
.A(n_337),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_330),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_330),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_330),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_327),
.B(n_212),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_330),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_342),
.Y(n_483)
);

AND2x4_ASAP7_75t_SL g484 ( 
.A(n_361),
.B(n_211),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_342),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_342),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_345),
.B(n_215),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_342),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_342),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_342),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_398),
.B(n_217),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_377),
.B(n_399),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_398),
.B(n_218),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_346),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_359),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_359),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_358),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_399),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_359),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_402),
.B(n_220),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_454),
.Y(n_502)
);

BUFx6f_ASAP7_75t_SL g503 ( 
.A(n_450),
.Y(n_503)
);

OR2x6_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_341),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_498),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_402),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_368),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_368),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_465),
.B(n_368),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_454),
.Y(n_511)
);

NOR2x1p5_ASAP7_75t_L g512 ( 
.A(n_440),
.B(n_391),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_351),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_351),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_356),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_409),
.B(n_369),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_409),
.B(n_378),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_392),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_415),
.A2(n_386),
.B(n_387),
.C(n_393),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_427),
.B(n_391),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_411),
.B(n_383),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_495),
.B(n_222),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_499),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_415),
.B(n_383),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_461),
.B(n_224),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_391),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_447),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_457),
.B(n_436),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_442),
.B(n_383),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_499),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_416),
.B(n_395),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_424),
.B(n_395),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_445),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_391),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_473),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_473),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_459),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_464),
.A2(n_362),
.B1(n_208),
.B2(n_302),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_433),
.A2(n_340),
.B1(n_358),
.B2(n_382),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_459),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_473),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_419),
.B(n_230),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_425),
.B(n_234),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_439),
.B(n_243),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_481),
.B(n_360),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_491),
.B(n_340),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_404),
.B(n_360),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

AND2x4_ASAP7_75t_SL g555 ( 
.A(n_484),
.B(n_225),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_433),
.A2(n_382),
.B1(n_397),
.B2(n_389),
.Y(n_556)
);

BUFx5_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_249),
.B1(n_226),
.B2(n_233),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_406),
.B(n_263),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_406),
.A2(n_397),
.B1(n_389),
.B2(n_241),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_469),
.B(n_389),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_452),
.B(n_397),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_248),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_251),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g567 ( 
.A(n_422),
.B(n_271),
.C(n_270),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_446),
.B(n_252),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_403),
.Y(n_570)
);

AND2x4_ASAP7_75t_SL g571 ( 
.A(n_438),
.B(n_288),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_407),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_407),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_403),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_437),
.A2(n_412),
.B(n_405),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_466),
.B(n_253),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_412),
.B(n_255),
.Y(n_577)
);

NOR3xp33_ASAP7_75t_L g578 ( 
.A(n_420),
.B(n_292),
.C(n_291),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_413),
.A2(n_294),
.B(n_301),
.C(n_304),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_413),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_414),
.A2(n_397),
.B1(n_310),
.B2(n_293),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_261),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_418),
.A2(n_305),
.B1(n_321),
.B2(n_322),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_431),
.B(n_202),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_414),
.B(n_273),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_408),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_417),
.Y(n_587)
);

CKINVDCx14_ASAP7_75t_R g588 ( 
.A(n_408),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_532),
.B(n_449),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_538),
.B(n_417),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_519),
.A2(n_431),
.B(n_460),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_519),
.A2(n_431),
.B(n_421),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_516),
.B(n_438),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_L g595 ( 
.A1(n_517),
.A2(n_430),
.B(n_428),
.Y(n_595)
);

NOR2x1_ASAP7_75t_L g596 ( 
.A(n_526),
.B(n_430),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_527),
.A2(n_363),
.B(n_344),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_575),
.A2(n_363),
.B(n_344),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_527),
.A2(n_536),
.B(n_564),
.Y(n_599)
);

AND3x2_ASAP7_75t_L g600 ( 
.A(n_525),
.B(n_16),
.C(n_18),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_515),
.A2(n_363),
.B(n_344),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_520),
.A2(n_373),
.B(n_458),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_514),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_508),
.A2(n_479),
.B(n_467),
.C(n_462),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_535),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_408),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_512),
.B(n_18),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_580),
.A2(n_474),
.B(n_472),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_567),
.A2(n_584),
.B1(n_518),
.B2(n_528),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_534),
.A2(n_474),
.B(n_472),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_279),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_553),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_559),
.B(n_19),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_553),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_505),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_281),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_SL g619 ( 
.A(n_559),
.B(n_286),
.C(n_284),
.Y(n_619)
);

AND2x4_ASAP7_75t_SL g620 ( 
.A(n_540),
.B(n_295),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_523),
.B(n_289),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_555),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_506),
.B(n_296),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_562),
.A2(n_475),
.B(n_471),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_571),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_521),
.A2(n_480),
.B(n_479),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_529),
.A2(n_565),
.B(n_566),
.C(n_572),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_522),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_587),
.A2(n_306),
.B1(n_316),
.B2(n_297),
.Y(n_630)
);

OAI321xp33_ASAP7_75t_L g631 ( 
.A1(n_561),
.A2(n_376),
.A3(n_401),
.B1(n_375),
.B2(n_346),
.C(n_348),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_581),
.B(n_303),
.C(n_300),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_533),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_584),
.A2(n_443),
.B(n_434),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_573),
.A2(n_426),
.B(n_423),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_541),
.B(n_309),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_586),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_503),
.A2(n_385),
.B1(n_381),
.B2(n_426),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_569),
.A2(n_511),
.B(n_502),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_586),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_539),
.A2(n_381),
.B1(n_385),
.B2(n_359),
.Y(n_644)
);

NAND2x1p5_ASAP7_75t_L g645 ( 
.A(n_546),
.B(n_496),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_545),
.A2(n_477),
.B(n_482),
.Y(n_646)
);

AO21x1_ASAP7_75t_L g647 ( 
.A1(n_560),
.A2(n_453),
.B(n_455),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_577),
.B(n_585),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_556),
.A2(n_385),
.B1(n_309),
.B2(n_453),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_531),
.A2(n_560),
.B(n_579),
.C(n_507),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_551),
.A2(n_483),
.B(n_485),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_504),
.A2(n_309),
.B1(n_455),
.B2(n_456),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_513),
.A2(n_490),
.B(n_486),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_563),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_544),
.B(n_20),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_21),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_504),
.A2(n_463),
.B1(n_468),
.B2(n_470),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_510),
.B(n_558),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_583),
.A2(n_470),
.B1(n_346),
.B2(n_348),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_570),
.A2(n_494),
.B(n_490),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_513),
.A2(n_488),
.B(n_489),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_576),
.B(n_22),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_574),
.A2(n_494),
.B(n_488),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_578),
.A2(n_375),
.B(n_348),
.C(n_349),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_552),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_549),
.B(n_22),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_552),
.B(n_530),
.Y(n_668)
);

BUFx8_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_623),
.B(n_524),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_SL g671 ( 
.A1(n_628),
.A2(n_582),
.B(n_568),
.C(n_547),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_614),
.B(n_23),
.Y(n_672)
);

OA22x2_ASAP7_75t_L g673 ( 
.A1(n_607),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_629),
.B(n_25),
.Y(n_674)
);

AO32x2_ASAP7_75t_L g675 ( 
.A1(n_652),
.A2(n_376),
.A3(n_348),
.B1(n_349),
.B2(n_353),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_632),
.B(n_26),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_593),
.B(n_616),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_647),
.A2(n_376),
.A3(n_348),
.B(n_349),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_609),
.B(n_26),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_622),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_613),
.B(n_28),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_617),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_666),
.B(n_29),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_605),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_610),
.B(n_29),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_650),
.A2(n_375),
.B(n_348),
.C(n_349),
.Y(n_686)
);

INVxp67_ASAP7_75t_SL g687 ( 
.A(n_590),
.Y(n_687)
);

AOI21xp33_ASAP7_75t_L g688 ( 
.A1(n_612),
.A2(n_30),
.B(n_31),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_648),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_632),
.B(n_500),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_635),
.B(n_30),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_636),
.A2(n_375),
.A3(n_349),
.B(n_353),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_591),
.A2(n_592),
.B(n_599),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_594),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_615),
.B(n_31),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_663),
.B(n_32),
.Y(n_696)
);

AO31x2_ASAP7_75t_L g697 ( 
.A1(n_597),
.A2(n_372),
.A3(n_401),
.B(n_390),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_658),
.B(n_496),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_658),
.B(n_496),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_657),
.B(n_496),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_602),
.A2(n_500),
.B(n_497),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_654),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_669),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_601),
.A2(n_476),
.B(n_346),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_607),
.B(n_497),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_624),
.A2(n_375),
.B1(n_353),
.B2(n_354),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_667),
.B(n_497),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_621),
.B(n_497),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_619),
.B(n_500),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_596),
.B(n_34),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_642),
.B(n_500),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_659),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_656),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_668),
.B(n_36),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_669),
.Y(n_715)
);

AOI211x1_ASAP7_75t_L g716 ( 
.A1(n_595),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_643),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_604),
.Y(n_718)
);

BUFx12f_ASAP7_75t_L g719 ( 
.A(n_645),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_655),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_653),
.A2(n_372),
.B(n_367),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_603),
.B(n_589),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_641),
.A2(n_500),
.B(n_372),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_662),
.A2(n_372),
.B(n_367),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_630),
.B(n_354),
.Y(n_725)
);

NAND3x1_ASAP7_75t_L g726 ( 
.A(n_600),
.B(n_44),
.C(n_47),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_606),
.B(n_49),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_622),
.Y(n_728)
);

BUFx12f_ASAP7_75t_L g729 ( 
.A(n_622),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_639),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_608),
.A2(n_50),
.B(n_51),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_639),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_644),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_611),
.A2(n_55),
.B(n_56),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_633),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_639),
.B(n_63),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_620),
.A2(n_66),
.B1(n_70),
.B2(n_78),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_640),
.B(n_83),
.Y(n_738)
);

NOR2x1_ASAP7_75t_SL g739 ( 
.A(n_634),
.B(n_85),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_661),
.A2(n_87),
.B(n_89),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_627),
.A2(n_96),
.B(n_97),
.Y(n_741)
);

BUFx4f_ASAP7_75t_L g742 ( 
.A(n_631),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_649),
.B(n_111),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_618),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_665),
.A2(n_118),
.A3(n_119),
.B(n_120),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_664),
.A2(n_121),
.B(n_123),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_637),
.A2(n_124),
.B(n_126),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_651),
.A2(n_129),
.B(n_132),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_660),
.B(n_133),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_644),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_638),
.B(n_141),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_646),
.A2(n_145),
.B(n_147),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_591),
.A2(n_156),
.B(n_157),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_614),
.B(n_158),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_163),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_614),
.B(n_166),
.Y(n_756)
);

AOI221xp5_ASAP7_75t_SL g757 ( 
.A1(n_650),
.A2(n_169),
.B1(n_172),
.B2(n_176),
.C(n_177),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_614),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_758)
);

AO21x1_ASAP7_75t_L g759 ( 
.A1(n_592),
.A2(n_181),
.B(n_187),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_625),
.A2(n_197),
.B(n_598),
.Y(n_760)
);

NOR2x1_ASAP7_75t_SL g761 ( 
.A(n_614),
.B(n_616),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_629),
.B(n_427),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_623),
.B(n_525),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_591),
.A2(n_592),
.B(n_599),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_591),
.A2(n_592),
.B(n_599),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_722),
.A2(n_689),
.B1(n_695),
.B2(n_674),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_730),
.B(n_677),
.Y(n_767)
);

BUFx12f_ASAP7_75t_L g768 ( 
.A(n_719),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_729),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_687),
.A2(n_683),
.B1(n_677),
.B2(n_713),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_762),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_761),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_680),
.Y(n_773)
);

AO21x2_ASAP7_75t_L g774 ( 
.A1(n_701),
.A2(n_704),
.B(n_760),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_730),
.B(n_683),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_680),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_688),
.A2(n_685),
.B(n_696),
.C(n_671),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_672),
.Y(n_778)
);

OAI21x1_ASAP7_75t_SL g779 ( 
.A1(n_739),
.A2(n_753),
.B(n_731),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_757),
.A2(n_724),
.B(n_721),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_673),
.A2(n_715),
.B1(n_703),
.B2(n_676),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_717),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_684),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_717),
.Y(n_784)
);

OA21x2_ASAP7_75t_L g785 ( 
.A1(n_740),
.A2(n_746),
.B(n_723),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_702),
.Y(n_786)
);

OAI21x1_ASAP7_75t_SL g787 ( 
.A1(n_747),
.A2(n_759),
.B(n_758),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

NOR2x1_ASAP7_75t_L g789 ( 
.A(n_738),
.B(n_737),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_763),
.B(n_670),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_733),
.A2(n_750),
.B1(n_718),
.B2(n_679),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_725),
.A2(n_748),
.B(n_734),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_694),
.B(n_712),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_SL g794 ( 
.A1(n_744),
.A2(n_681),
.B(n_755),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_742),
.A2(n_691),
.B1(n_716),
.B2(n_749),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_720),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_705),
.B(n_732),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_710),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_710),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_709),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_711),
.B(n_692),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_752),
.A2(n_741),
.B(n_743),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_SL g803 ( 
.A1(n_742),
.A2(n_735),
.B1(n_726),
.B2(n_698),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_692),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_692),
.Y(n_805)
);

CKINVDCx6p67_ASAP7_75t_R g806 ( 
.A(n_680),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_706),
.A2(n_736),
.B(n_754),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_699),
.A2(n_756),
.B(n_727),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_SL g809 ( 
.A(n_700),
.B(n_751),
.C(n_707),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_728),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_728),
.B(n_678),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_728),
.B(n_708),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_678),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_697),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_745),
.A2(n_669),
.B1(n_722),
.B2(n_504),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_675),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_745),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_682),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_761),
.A2(n_559),
.B1(n_669),
.B2(n_555),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_762),
.B(n_677),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_719),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_677),
.B(n_761),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_677),
.B(n_629),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_719),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_729),
.B(n_730),
.Y(n_826)
);

AO31x2_ASAP7_75t_L g827 ( 
.A1(n_686),
.A2(n_693),
.A3(n_765),
.B(n_764),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_682),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_682),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_677),
.B(n_629),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_629),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_689),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_677),
.B(n_629),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_677),
.B(n_761),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_729),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_682),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_722),
.A2(n_669),
.B1(n_504),
.B2(n_535),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_729),
.B(n_730),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_722),
.A2(n_669),
.B1(n_504),
.B2(n_535),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_762),
.B(n_677),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_682),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_719),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_687),
.B(n_614),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_688),
.A2(n_650),
.B(n_615),
.C(n_543),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_762),
.B(n_677),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_677),
.B(n_629),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_687),
.A2(n_615),
.B1(n_559),
.B2(n_499),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_818),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_828),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_823),
.Y(n_851)
);

AO21x1_ASAP7_75t_SL g852 ( 
.A1(n_770),
.A2(n_844),
.B(n_811),
.Y(n_852)
);

CKINVDCx6p67_ASAP7_75t_R g853 ( 
.A(n_768),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_783),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_823),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_835),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_776),
.Y(n_857)
);

AO21x1_ASAP7_75t_SL g858 ( 
.A1(n_770),
.A2(n_844),
.B(n_798),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_829),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_791),
.B(n_782),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_784),
.B(n_837),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_801),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_822),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_776),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_825),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_842),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_793),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_796),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_821),
.B(n_841),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_846),
.B(n_771),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_824),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_843),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_831),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_810),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_843),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_832),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_771),
.B(n_833),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_834),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

NAND4xp25_ASAP7_75t_L g880 ( 
.A(n_766),
.B(n_840),
.C(n_838),
.D(n_790),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_835),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_769),
.Y(n_882)
);

NOR2x1_ASAP7_75t_R g883 ( 
.A(n_769),
.B(n_830),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_788),
.Y(n_885)
);

INVx6_ASAP7_75t_L g886 ( 
.A(n_773),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_830),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_836),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_772),
.B(n_800),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_786),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_786),
.B(n_819),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_814),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_L g893 ( 
.A1(n_848),
.A2(n_781),
.B1(n_845),
.B2(n_778),
.C(n_777),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_775),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_813),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_797),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_836),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_826),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_827),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_767),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_806),
.Y(n_901)
);

AO21x1_ASAP7_75t_L g902 ( 
.A1(n_795),
.A2(n_817),
.B(n_804),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_826),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_839),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_799),
.B(n_789),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_839),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_773),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_776),
.Y(n_908)
);

BUFx8_ASAP7_75t_L g909 ( 
.A(n_805),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_815),
.B(n_809),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_812),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_803),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_794),
.B(n_795),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_816),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_808),
.B(n_802),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_780),
.Y(n_916)
);

INVxp33_ASAP7_75t_L g917 ( 
.A(n_779),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_880),
.A2(n_787),
.B1(n_808),
.B2(n_802),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_909),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_862),
.A2(n_785),
.B1(n_792),
.B2(n_807),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_905),
.B(n_774),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_905),
.B(n_785),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_909),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_892),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_860),
.B(n_892),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_867),
.B(n_871),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_852),
.B(n_870),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_873),
.B(n_876),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_910),
.A2(n_893),
.B1(n_912),
.B2(n_891),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_849),
.B(n_850),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_890),
.B(n_914),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_859),
.B(n_866),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_896),
.B(n_861),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_886),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_861),
.B(n_895),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_868),
.B(n_899),
.Y(n_937)
);

BUFx8_ASAP7_75t_L g938 ( 
.A(n_874),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_877),
.B(n_878),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_888),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_879),
.B(n_893),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_869),
.B(n_884),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_897),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_916),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_913),
.B(n_858),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_857),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_854),
.B(n_865),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_851),
.B(n_855),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_855),
.B(n_856),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_889),
.B(n_881),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_889),
.B(n_881),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_931),
.B(n_911),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_919),
.B(n_898),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_933),
.B(n_906),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_936),
.B(n_926),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_925),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_934),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_944),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_919),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_943),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_936),
.B(n_915),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_921),
.B(n_917),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_944),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_925),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_934),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_924),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_939),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_939),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_923),
.B(n_853),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_926),
.B(n_932),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_922),
.B(n_902),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_927),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_937),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_960),
.B(n_941),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_955),
.B(n_928),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_959),
.B(n_919),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_971),
.A2(n_930),
.B(n_918),
.Y(n_977)
);

AND2x2_ASAP7_75t_SL g978 ( 
.A(n_959),
.B(n_945),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_964),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_964),
.B(n_945),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_970),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_970),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_955),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_966),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_972),
.B(n_940),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_961),
.B(n_928),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_961),
.B(n_942),
.Y(n_987)
);

NAND2x1_ASAP7_75t_L g988 ( 
.A(n_976),
.B(n_959),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_980),
.B(n_962),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_976),
.B(n_953),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_984),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_975),
.B(n_967),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_983),
.Y(n_993)
);

AO31x2_ASAP7_75t_L g994 ( 
.A1(n_974),
.A2(n_958),
.A3(n_963),
.B(n_920),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_976),
.B(n_956),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_980),
.B(n_973),
.Y(n_996)
);

NOR2x1p5_ASAP7_75t_L g997 ( 
.A(n_986),
.B(n_919),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_987),
.B(n_968),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_978),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_978),
.A2(n_923),
.B(n_969),
.C(n_898),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_974),
.B(n_938),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_1001),
.B(n_981),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_989),
.B(n_982),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_993),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_992),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_998),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_996),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_997),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_988),
.Y(n_1011)
);

AOI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_1000),
.A2(n_977),
.B1(n_985),
.B2(n_957),
.C(n_965),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_988),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_995),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1005),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_1007),
.B(n_947),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_1011),
.B(n_990),
.Y(n_1017)
);

INVxp33_ASAP7_75t_L g1018 ( 
.A(n_1013),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1007),
.A2(n_999),
.B1(n_1012),
.B2(n_990),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1008),
.B(n_1006),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1017),
.A2(n_1019),
.B(n_1018),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_1002),
.B1(n_1014),
.B2(n_1010),
.Y(n_1022)
);

AOI222xp33_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_985),
.B1(n_1005),
.B2(n_1003),
.C1(n_954),
.C2(n_1009),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1023),
.B(n_1020),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_1021),
.B(n_883),
.C(n_904),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_SL g1026 ( 
.A(n_1024),
.B(n_872),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_L g1028 ( 
.A(n_1027),
.B(n_882),
.C(n_875),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_1026),
.B(n_882),
.C(n_887),
.Y(n_1029)
);

XOR2xp5_ASAP7_75t_L g1030 ( 
.A(n_1028),
.B(n_863),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1029),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1031),
.A2(n_863),
.B1(n_953),
.B2(n_995),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1031),
.B(n_994),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1032),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1034),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_1033),
.B(n_938),
.Y(n_1037)
);

AOI321xp33_ASAP7_75t_L g1038 ( 
.A1(n_1032),
.A2(n_903),
.A3(n_938),
.B1(n_894),
.B2(n_935),
.C(n_929),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

XNOR2x1_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_938),
.Y(n_1040)
);

AO22x2_ASAP7_75t_L g1041 ( 
.A1(n_1037),
.A2(n_907),
.B1(n_900),
.B2(n_1004),
.Y(n_1041)
);

AOI22x1_ASAP7_75t_L g1042 ( 
.A1(n_1038),
.A2(n_901),
.B1(n_885),
.B2(n_953),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1037),
.A2(n_900),
.B(n_952),
.Y(n_1043)
);

XNOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_935),
.Y(n_1044)
);

OAI22x1_ASAP7_75t_L g1045 ( 
.A1(n_1039),
.A2(n_979),
.B1(n_948),
.B2(n_949),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1040),
.A2(n_935),
.B(n_979),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1046),
.A2(n_1044),
.B(n_1041),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_1045),
.A2(n_1043),
.B(n_1042),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1047),
.A2(n_950),
.B(n_951),
.Y(n_1049)
);

AOI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_1049),
.A2(n_1048),
.B1(n_908),
.B2(n_864),
.C(n_857),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_1050),
.A2(n_908),
.B(n_946),
.Y(n_1051)
);


endmodule